module Switch( // @[:@3.2]
  input  [3:0]  io_inAddr_0, // @[:@6.4]
  input  [3:0]  io_inAddr_1, // @[:@6.4]
  input  [3:0]  io_inAddr_2, // @[:@6.4]
  input  [3:0]  io_inAddr_3, // @[:@6.4]
  input  [3:0]  io_inAddr_4, // @[:@6.4]
  input  [3:0]  io_inAddr_5, // @[:@6.4]
  input  [3:0]  io_inAddr_6, // @[:@6.4]
  input  [3:0]  io_inAddr_7, // @[:@6.4]
  input  [3:0]  io_inAddr_8, // @[:@6.4]
  input  [3:0]  io_inAddr_9, // @[:@6.4]
  input  [3:0]  io_inAddr_10, // @[:@6.4]
  input  [3:0]  io_inAddr_11, // @[:@6.4]
  input  [3:0]  io_inAddr_12, // @[:@6.4]
  input  [3:0]  io_inAddr_13, // @[:@6.4]
  input  [3:0]  io_inAddr_14, // @[:@6.4]
  input  [3:0]  io_inAddr_15, // @[:@6.4]
  input  [47:0] io_inData_0, // @[:@6.4]
  input  [47:0] io_inData_1, // @[:@6.4]
  input  [47:0] io_inData_2, // @[:@6.4]
  input  [47:0] io_inData_3, // @[:@6.4]
  input  [47:0] io_inData_4, // @[:@6.4]
  input  [47:0] io_inData_5, // @[:@6.4]
  input  [47:0] io_inData_6, // @[:@6.4]
  input  [47:0] io_inData_7, // @[:@6.4]
  input  [47:0] io_inData_8, // @[:@6.4]
  input  [47:0] io_inData_9, // @[:@6.4]
  input  [47:0] io_inData_10, // @[:@6.4]
  input  [47:0] io_inData_11, // @[:@6.4]
  input  [47:0] io_inData_12, // @[:@6.4]
  input  [47:0] io_inData_13, // @[:@6.4]
  input  [47:0] io_inData_14, // @[:@6.4]
  input  [47:0] io_inData_15, // @[:@6.4]
  input         io_inValid_0, // @[:@6.4]
  input         io_inValid_1, // @[:@6.4]
  input         io_inValid_2, // @[:@6.4]
  input         io_inValid_3, // @[:@6.4]
  input         io_inValid_4, // @[:@6.4]
  input         io_inValid_5, // @[:@6.4]
  input         io_inValid_6, // @[:@6.4]
  input         io_inValid_7, // @[:@6.4]
  input         io_inValid_8, // @[:@6.4]
  input         io_inValid_9, // @[:@6.4]
  input         io_inValid_10, // @[:@6.4]
  input         io_inValid_11, // @[:@6.4]
  input         io_inValid_12, // @[:@6.4]
  input         io_inValid_13, // @[:@6.4]
  input         io_inValid_14, // @[:@6.4]
  input         io_inValid_15, // @[:@6.4]
  output        io_outAck_0, // @[:@6.4]
  output        io_outAck_1, // @[:@6.4]
  output        io_outAck_2, // @[:@6.4]
  output        io_outAck_3, // @[:@6.4]
  output        io_outAck_4, // @[:@6.4]
  output        io_outAck_5, // @[:@6.4]
  output        io_outAck_6, // @[:@6.4]
  output        io_outAck_7, // @[:@6.4]
  output        io_outAck_8, // @[:@6.4]
  output        io_outAck_9, // @[:@6.4]
  output        io_outAck_10, // @[:@6.4]
  output        io_outAck_11, // @[:@6.4]
  output        io_outAck_12, // @[:@6.4]
  output        io_outAck_13, // @[:@6.4]
  output        io_outAck_14, // @[:@6.4]
  output        io_outAck_15, // @[:@6.4]
  output [47:0] io_outData_0, // @[:@6.4]
  output [47:0] io_outData_1, // @[:@6.4]
  output [47:0] io_outData_2, // @[:@6.4]
  output [47:0] io_outData_3, // @[:@6.4]
  output [47:0] io_outData_4, // @[:@6.4]
  output [47:0] io_outData_5, // @[:@6.4]
  output [47:0] io_outData_6, // @[:@6.4]
  output [47:0] io_outData_7, // @[:@6.4]
  output [47:0] io_outData_8, // @[:@6.4]
  output [47:0] io_outData_9, // @[:@6.4]
  output [47:0] io_outData_10, // @[:@6.4]
  output [47:0] io_outData_11, // @[:@6.4]
  output [47:0] io_outData_12, // @[:@6.4]
  output [47:0] io_outData_13, // @[:@6.4]
  output [47:0] io_outData_14, // @[:@6.4]
  output [47:0] io_outData_15, // @[:@6.4]
  output        io_outValid_0, // @[:@6.4]
  output        io_outValid_1, // @[:@6.4]
  output        io_outValid_2, // @[:@6.4]
  output        io_outValid_3, // @[:@6.4]
  output        io_outValid_4, // @[:@6.4]
  output        io_outValid_5, // @[:@6.4]
  output        io_outValid_6, // @[:@6.4]
  output        io_outValid_7, // @[:@6.4]
  output        io_outValid_8, // @[:@6.4]
  output        io_outValid_9, // @[:@6.4]
  output        io_outValid_10, // @[:@6.4]
  output        io_outValid_11, // @[:@6.4]
  output        io_outValid_12, // @[:@6.4]
  output        io_outValid_13, // @[:@6.4]
  output        io_outValid_14, // @[:@6.4]
  output        io_outValid_15 // @[:@6.4]
);
  wire  _T_1382; // @[Switch.scala 30:53:@10.4]
  wire  valid_0_0; // @[Switch.scala 30:36:@11.4]
  wire  _T_1385; // @[Switch.scala 30:53:@13.4]
  wire  valid_0_1; // @[Switch.scala 30:36:@14.4]
  wire  _T_1388; // @[Switch.scala 30:53:@16.4]
  wire  valid_0_2; // @[Switch.scala 30:36:@17.4]
  wire  _T_1391; // @[Switch.scala 30:53:@19.4]
  wire  valid_0_3; // @[Switch.scala 30:36:@20.4]
  wire  _T_1394; // @[Switch.scala 30:53:@22.4]
  wire  valid_0_4; // @[Switch.scala 30:36:@23.4]
  wire  _T_1397; // @[Switch.scala 30:53:@25.4]
  wire  valid_0_5; // @[Switch.scala 30:36:@26.4]
  wire  _T_1400; // @[Switch.scala 30:53:@28.4]
  wire  valid_0_6; // @[Switch.scala 30:36:@29.4]
  wire  _T_1403; // @[Switch.scala 30:53:@31.4]
  wire  valid_0_7; // @[Switch.scala 30:36:@32.4]
  wire  _T_1406; // @[Switch.scala 30:53:@34.4]
  wire  valid_0_8; // @[Switch.scala 30:36:@35.4]
  wire  _T_1409; // @[Switch.scala 30:53:@37.4]
  wire  valid_0_9; // @[Switch.scala 30:36:@38.4]
  wire  _T_1412; // @[Switch.scala 30:53:@40.4]
  wire  valid_0_10; // @[Switch.scala 30:36:@41.4]
  wire  _T_1415; // @[Switch.scala 30:53:@43.4]
  wire  valid_0_11; // @[Switch.scala 30:36:@44.4]
  wire  _T_1418; // @[Switch.scala 30:53:@46.4]
  wire  valid_0_12; // @[Switch.scala 30:36:@47.4]
  wire  _T_1421; // @[Switch.scala 30:53:@49.4]
  wire  valid_0_13; // @[Switch.scala 30:36:@50.4]
  wire  _T_1424; // @[Switch.scala 30:53:@52.4]
  wire  valid_0_14; // @[Switch.scala 30:36:@53.4]
  wire  _T_1427; // @[Switch.scala 30:53:@55.4]
  wire  valid_0_15; // @[Switch.scala 30:36:@56.4]
  wire [3:0] _T_1445; // @[Mux.scala 31:69:@58.4]
  wire [3:0] _T_1446; // @[Mux.scala 31:69:@59.4]
  wire [3:0] _T_1447; // @[Mux.scala 31:69:@60.4]
  wire [3:0] _T_1448; // @[Mux.scala 31:69:@61.4]
  wire [3:0] _T_1449; // @[Mux.scala 31:69:@62.4]
  wire [3:0] _T_1450; // @[Mux.scala 31:69:@63.4]
  wire [3:0] _T_1451; // @[Mux.scala 31:69:@64.4]
  wire [3:0] _T_1452; // @[Mux.scala 31:69:@65.4]
  wire [3:0] _T_1453; // @[Mux.scala 31:69:@66.4]
  wire [3:0] _T_1454; // @[Mux.scala 31:69:@67.4]
  wire [3:0] _T_1455; // @[Mux.scala 31:69:@68.4]
  wire [3:0] _T_1456; // @[Mux.scala 31:69:@69.4]
  wire [3:0] _T_1457; // @[Mux.scala 31:69:@70.4]
  wire [3:0] _T_1458; // @[Mux.scala 31:69:@71.4]
  wire [3:0] select_0; // @[Mux.scala 31:69:@72.4]
  wire [47:0] _GEN_1; // @[Switch.scala 33:19:@74.4]
  wire [47:0] _GEN_2; // @[Switch.scala 33:19:@74.4]
  wire [47:0] _GEN_3; // @[Switch.scala 33:19:@74.4]
  wire [47:0] _GEN_4; // @[Switch.scala 33:19:@74.4]
  wire [47:0] _GEN_5; // @[Switch.scala 33:19:@74.4]
  wire [47:0] _GEN_6; // @[Switch.scala 33:19:@74.4]
  wire [47:0] _GEN_7; // @[Switch.scala 33:19:@74.4]
  wire [47:0] _GEN_8; // @[Switch.scala 33:19:@74.4]
  wire [47:0] _GEN_9; // @[Switch.scala 33:19:@74.4]
  wire [47:0] _GEN_10; // @[Switch.scala 33:19:@74.4]
  wire [47:0] _GEN_11; // @[Switch.scala 33:19:@74.4]
  wire [47:0] _GEN_12; // @[Switch.scala 33:19:@74.4]
  wire [47:0] _GEN_13; // @[Switch.scala 33:19:@74.4]
  wire [47:0] _GEN_14; // @[Switch.scala 33:19:@74.4]
  wire [7:0] _T_1467; // @[Switch.scala 34:32:@81.4]
  wire [15:0] _T_1475; // @[Switch.scala 34:32:@89.4]
  wire  _T_1479; // @[Switch.scala 30:53:@92.4]
  wire  valid_1_0; // @[Switch.scala 30:36:@93.4]
  wire  _T_1482; // @[Switch.scala 30:53:@95.4]
  wire  valid_1_1; // @[Switch.scala 30:36:@96.4]
  wire  _T_1485; // @[Switch.scala 30:53:@98.4]
  wire  valid_1_2; // @[Switch.scala 30:36:@99.4]
  wire  _T_1488; // @[Switch.scala 30:53:@101.4]
  wire  valid_1_3; // @[Switch.scala 30:36:@102.4]
  wire  _T_1491; // @[Switch.scala 30:53:@104.4]
  wire  valid_1_4; // @[Switch.scala 30:36:@105.4]
  wire  _T_1494; // @[Switch.scala 30:53:@107.4]
  wire  valid_1_5; // @[Switch.scala 30:36:@108.4]
  wire  _T_1497; // @[Switch.scala 30:53:@110.4]
  wire  valid_1_6; // @[Switch.scala 30:36:@111.4]
  wire  _T_1500; // @[Switch.scala 30:53:@113.4]
  wire  valid_1_7; // @[Switch.scala 30:36:@114.4]
  wire  _T_1503; // @[Switch.scala 30:53:@116.4]
  wire  valid_1_8; // @[Switch.scala 30:36:@117.4]
  wire  _T_1506; // @[Switch.scala 30:53:@119.4]
  wire  valid_1_9; // @[Switch.scala 30:36:@120.4]
  wire  _T_1509; // @[Switch.scala 30:53:@122.4]
  wire  valid_1_10; // @[Switch.scala 30:36:@123.4]
  wire  _T_1512; // @[Switch.scala 30:53:@125.4]
  wire  valid_1_11; // @[Switch.scala 30:36:@126.4]
  wire  _T_1515; // @[Switch.scala 30:53:@128.4]
  wire  valid_1_12; // @[Switch.scala 30:36:@129.4]
  wire  _T_1518; // @[Switch.scala 30:53:@131.4]
  wire  valid_1_13; // @[Switch.scala 30:36:@132.4]
  wire  _T_1521; // @[Switch.scala 30:53:@134.4]
  wire  valid_1_14; // @[Switch.scala 30:36:@135.4]
  wire  _T_1524; // @[Switch.scala 30:53:@137.4]
  wire  valid_1_15; // @[Switch.scala 30:36:@138.4]
  wire [3:0] _T_1542; // @[Mux.scala 31:69:@140.4]
  wire [3:0] _T_1543; // @[Mux.scala 31:69:@141.4]
  wire [3:0] _T_1544; // @[Mux.scala 31:69:@142.4]
  wire [3:0] _T_1545; // @[Mux.scala 31:69:@143.4]
  wire [3:0] _T_1546; // @[Mux.scala 31:69:@144.4]
  wire [3:0] _T_1547; // @[Mux.scala 31:69:@145.4]
  wire [3:0] _T_1548; // @[Mux.scala 31:69:@146.4]
  wire [3:0] _T_1549; // @[Mux.scala 31:69:@147.4]
  wire [3:0] _T_1550; // @[Mux.scala 31:69:@148.4]
  wire [3:0] _T_1551; // @[Mux.scala 31:69:@149.4]
  wire [3:0] _T_1552; // @[Mux.scala 31:69:@150.4]
  wire [3:0] _T_1553; // @[Mux.scala 31:69:@151.4]
  wire [3:0] _T_1554; // @[Mux.scala 31:69:@152.4]
  wire [3:0] _T_1555; // @[Mux.scala 31:69:@153.4]
  wire [3:0] select_1; // @[Mux.scala 31:69:@154.4]
  wire [47:0] _GEN_17; // @[Switch.scala 33:19:@156.4]
  wire [47:0] _GEN_18; // @[Switch.scala 33:19:@156.4]
  wire [47:0] _GEN_19; // @[Switch.scala 33:19:@156.4]
  wire [47:0] _GEN_20; // @[Switch.scala 33:19:@156.4]
  wire [47:0] _GEN_21; // @[Switch.scala 33:19:@156.4]
  wire [47:0] _GEN_22; // @[Switch.scala 33:19:@156.4]
  wire [47:0] _GEN_23; // @[Switch.scala 33:19:@156.4]
  wire [47:0] _GEN_24; // @[Switch.scala 33:19:@156.4]
  wire [47:0] _GEN_25; // @[Switch.scala 33:19:@156.4]
  wire [47:0] _GEN_26; // @[Switch.scala 33:19:@156.4]
  wire [47:0] _GEN_27; // @[Switch.scala 33:19:@156.4]
  wire [47:0] _GEN_28; // @[Switch.scala 33:19:@156.4]
  wire [47:0] _GEN_29; // @[Switch.scala 33:19:@156.4]
  wire [47:0] _GEN_30; // @[Switch.scala 33:19:@156.4]
  wire [7:0] _T_1564; // @[Switch.scala 34:32:@163.4]
  wire [15:0] _T_1572; // @[Switch.scala 34:32:@171.4]
  wire  _T_1576; // @[Switch.scala 30:53:@174.4]
  wire  valid_2_0; // @[Switch.scala 30:36:@175.4]
  wire  _T_1579; // @[Switch.scala 30:53:@177.4]
  wire  valid_2_1; // @[Switch.scala 30:36:@178.4]
  wire  _T_1582; // @[Switch.scala 30:53:@180.4]
  wire  valid_2_2; // @[Switch.scala 30:36:@181.4]
  wire  _T_1585; // @[Switch.scala 30:53:@183.4]
  wire  valid_2_3; // @[Switch.scala 30:36:@184.4]
  wire  _T_1588; // @[Switch.scala 30:53:@186.4]
  wire  valid_2_4; // @[Switch.scala 30:36:@187.4]
  wire  _T_1591; // @[Switch.scala 30:53:@189.4]
  wire  valid_2_5; // @[Switch.scala 30:36:@190.4]
  wire  _T_1594; // @[Switch.scala 30:53:@192.4]
  wire  valid_2_6; // @[Switch.scala 30:36:@193.4]
  wire  _T_1597; // @[Switch.scala 30:53:@195.4]
  wire  valid_2_7; // @[Switch.scala 30:36:@196.4]
  wire  _T_1600; // @[Switch.scala 30:53:@198.4]
  wire  valid_2_8; // @[Switch.scala 30:36:@199.4]
  wire  _T_1603; // @[Switch.scala 30:53:@201.4]
  wire  valid_2_9; // @[Switch.scala 30:36:@202.4]
  wire  _T_1606; // @[Switch.scala 30:53:@204.4]
  wire  valid_2_10; // @[Switch.scala 30:36:@205.4]
  wire  _T_1609; // @[Switch.scala 30:53:@207.4]
  wire  valid_2_11; // @[Switch.scala 30:36:@208.4]
  wire  _T_1612; // @[Switch.scala 30:53:@210.4]
  wire  valid_2_12; // @[Switch.scala 30:36:@211.4]
  wire  _T_1615; // @[Switch.scala 30:53:@213.4]
  wire  valid_2_13; // @[Switch.scala 30:36:@214.4]
  wire  _T_1618; // @[Switch.scala 30:53:@216.4]
  wire  valid_2_14; // @[Switch.scala 30:36:@217.4]
  wire  _T_1621; // @[Switch.scala 30:53:@219.4]
  wire  valid_2_15; // @[Switch.scala 30:36:@220.4]
  wire [3:0] _T_1639; // @[Mux.scala 31:69:@222.4]
  wire [3:0] _T_1640; // @[Mux.scala 31:69:@223.4]
  wire [3:0] _T_1641; // @[Mux.scala 31:69:@224.4]
  wire [3:0] _T_1642; // @[Mux.scala 31:69:@225.4]
  wire [3:0] _T_1643; // @[Mux.scala 31:69:@226.4]
  wire [3:0] _T_1644; // @[Mux.scala 31:69:@227.4]
  wire [3:0] _T_1645; // @[Mux.scala 31:69:@228.4]
  wire [3:0] _T_1646; // @[Mux.scala 31:69:@229.4]
  wire [3:0] _T_1647; // @[Mux.scala 31:69:@230.4]
  wire [3:0] _T_1648; // @[Mux.scala 31:69:@231.4]
  wire [3:0] _T_1649; // @[Mux.scala 31:69:@232.4]
  wire [3:0] _T_1650; // @[Mux.scala 31:69:@233.4]
  wire [3:0] _T_1651; // @[Mux.scala 31:69:@234.4]
  wire [3:0] _T_1652; // @[Mux.scala 31:69:@235.4]
  wire [3:0] select_2; // @[Mux.scala 31:69:@236.4]
  wire [47:0] _GEN_33; // @[Switch.scala 33:19:@238.4]
  wire [47:0] _GEN_34; // @[Switch.scala 33:19:@238.4]
  wire [47:0] _GEN_35; // @[Switch.scala 33:19:@238.4]
  wire [47:0] _GEN_36; // @[Switch.scala 33:19:@238.4]
  wire [47:0] _GEN_37; // @[Switch.scala 33:19:@238.4]
  wire [47:0] _GEN_38; // @[Switch.scala 33:19:@238.4]
  wire [47:0] _GEN_39; // @[Switch.scala 33:19:@238.4]
  wire [47:0] _GEN_40; // @[Switch.scala 33:19:@238.4]
  wire [47:0] _GEN_41; // @[Switch.scala 33:19:@238.4]
  wire [47:0] _GEN_42; // @[Switch.scala 33:19:@238.4]
  wire [47:0] _GEN_43; // @[Switch.scala 33:19:@238.4]
  wire [47:0] _GEN_44; // @[Switch.scala 33:19:@238.4]
  wire [47:0] _GEN_45; // @[Switch.scala 33:19:@238.4]
  wire [47:0] _GEN_46; // @[Switch.scala 33:19:@238.4]
  wire [7:0] _T_1661; // @[Switch.scala 34:32:@245.4]
  wire [15:0] _T_1669; // @[Switch.scala 34:32:@253.4]
  wire  _T_1673; // @[Switch.scala 30:53:@256.4]
  wire  valid_3_0; // @[Switch.scala 30:36:@257.4]
  wire  _T_1676; // @[Switch.scala 30:53:@259.4]
  wire  valid_3_1; // @[Switch.scala 30:36:@260.4]
  wire  _T_1679; // @[Switch.scala 30:53:@262.4]
  wire  valid_3_2; // @[Switch.scala 30:36:@263.4]
  wire  _T_1682; // @[Switch.scala 30:53:@265.4]
  wire  valid_3_3; // @[Switch.scala 30:36:@266.4]
  wire  _T_1685; // @[Switch.scala 30:53:@268.4]
  wire  valid_3_4; // @[Switch.scala 30:36:@269.4]
  wire  _T_1688; // @[Switch.scala 30:53:@271.4]
  wire  valid_3_5; // @[Switch.scala 30:36:@272.4]
  wire  _T_1691; // @[Switch.scala 30:53:@274.4]
  wire  valid_3_6; // @[Switch.scala 30:36:@275.4]
  wire  _T_1694; // @[Switch.scala 30:53:@277.4]
  wire  valid_3_7; // @[Switch.scala 30:36:@278.4]
  wire  _T_1697; // @[Switch.scala 30:53:@280.4]
  wire  valid_3_8; // @[Switch.scala 30:36:@281.4]
  wire  _T_1700; // @[Switch.scala 30:53:@283.4]
  wire  valid_3_9; // @[Switch.scala 30:36:@284.4]
  wire  _T_1703; // @[Switch.scala 30:53:@286.4]
  wire  valid_3_10; // @[Switch.scala 30:36:@287.4]
  wire  _T_1706; // @[Switch.scala 30:53:@289.4]
  wire  valid_3_11; // @[Switch.scala 30:36:@290.4]
  wire  _T_1709; // @[Switch.scala 30:53:@292.4]
  wire  valid_3_12; // @[Switch.scala 30:36:@293.4]
  wire  _T_1712; // @[Switch.scala 30:53:@295.4]
  wire  valid_3_13; // @[Switch.scala 30:36:@296.4]
  wire  _T_1715; // @[Switch.scala 30:53:@298.4]
  wire  valid_3_14; // @[Switch.scala 30:36:@299.4]
  wire  _T_1718; // @[Switch.scala 30:53:@301.4]
  wire  valid_3_15; // @[Switch.scala 30:36:@302.4]
  wire [3:0] _T_1736; // @[Mux.scala 31:69:@304.4]
  wire [3:0] _T_1737; // @[Mux.scala 31:69:@305.4]
  wire [3:0] _T_1738; // @[Mux.scala 31:69:@306.4]
  wire [3:0] _T_1739; // @[Mux.scala 31:69:@307.4]
  wire [3:0] _T_1740; // @[Mux.scala 31:69:@308.4]
  wire [3:0] _T_1741; // @[Mux.scala 31:69:@309.4]
  wire [3:0] _T_1742; // @[Mux.scala 31:69:@310.4]
  wire [3:0] _T_1743; // @[Mux.scala 31:69:@311.4]
  wire [3:0] _T_1744; // @[Mux.scala 31:69:@312.4]
  wire [3:0] _T_1745; // @[Mux.scala 31:69:@313.4]
  wire [3:0] _T_1746; // @[Mux.scala 31:69:@314.4]
  wire [3:0] _T_1747; // @[Mux.scala 31:69:@315.4]
  wire [3:0] _T_1748; // @[Mux.scala 31:69:@316.4]
  wire [3:0] _T_1749; // @[Mux.scala 31:69:@317.4]
  wire [3:0] select_3; // @[Mux.scala 31:69:@318.4]
  wire [47:0] _GEN_49; // @[Switch.scala 33:19:@320.4]
  wire [47:0] _GEN_50; // @[Switch.scala 33:19:@320.4]
  wire [47:0] _GEN_51; // @[Switch.scala 33:19:@320.4]
  wire [47:0] _GEN_52; // @[Switch.scala 33:19:@320.4]
  wire [47:0] _GEN_53; // @[Switch.scala 33:19:@320.4]
  wire [47:0] _GEN_54; // @[Switch.scala 33:19:@320.4]
  wire [47:0] _GEN_55; // @[Switch.scala 33:19:@320.4]
  wire [47:0] _GEN_56; // @[Switch.scala 33:19:@320.4]
  wire [47:0] _GEN_57; // @[Switch.scala 33:19:@320.4]
  wire [47:0] _GEN_58; // @[Switch.scala 33:19:@320.4]
  wire [47:0] _GEN_59; // @[Switch.scala 33:19:@320.4]
  wire [47:0] _GEN_60; // @[Switch.scala 33:19:@320.4]
  wire [47:0] _GEN_61; // @[Switch.scala 33:19:@320.4]
  wire [47:0] _GEN_62; // @[Switch.scala 33:19:@320.4]
  wire [7:0] _T_1758; // @[Switch.scala 34:32:@327.4]
  wire [15:0] _T_1766; // @[Switch.scala 34:32:@335.4]
  wire  _T_1770; // @[Switch.scala 30:53:@338.4]
  wire  valid_4_0; // @[Switch.scala 30:36:@339.4]
  wire  _T_1773; // @[Switch.scala 30:53:@341.4]
  wire  valid_4_1; // @[Switch.scala 30:36:@342.4]
  wire  _T_1776; // @[Switch.scala 30:53:@344.4]
  wire  valid_4_2; // @[Switch.scala 30:36:@345.4]
  wire  _T_1779; // @[Switch.scala 30:53:@347.4]
  wire  valid_4_3; // @[Switch.scala 30:36:@348.4]
  wire  _T_1782; // @[Switch.scala 30:53:@350.4]
  wire  valid_4_4; // @[Switch.scala 30:36:@351.4]
  wire  _T_1785; // @[Switch.scala 30:53:@353.4]
  wire  valid_4_5; // @[Switch.scala 30:36:@354.4]
  wire  _T_1788; // @[Switch.scala 30:53:@356.4]
  wire  valid_4_6; // @[Switch.scala 30:36:@357.4]
  wire  _T_1791; // @[Switch.scala 30:53:@359.4]
  wire  valid_4_7; // @[Switch.scala 30:36:@360.4]
  wire  _T_1794; // @[Switch.scala 30:53:@362.4]
  wire  valid_4_8; // @[Switch.scala 30:36:@363.4]
  wire  _T_1797; // @[Switch.scala 30:53:@365.4]
  wire  valid_4_9; // @[Switch.scala 30:36:@366.4]
  wire  _T_1800; // @[Switch.scala 30:53:@368.4]
  wire  valid_4_10; // @[Switch.scala 30:36:@369.4]
  wire  _T_1803; // @[Switch.scala 30:53:@371.4]
  wire  valid_4_11; // @[Switch.scala 30:36:@372.4]
  wire  _T_1806; // @[Switch.scala 30:53:@374.4]
  wire  valid_4_12; // @[Switch.scala 30:36:@375.4]
  wire  _T_1809; // @[Switch.scala 30:53:@377.4]
  wire  valid_4_13; // @[Switch.scala 30:36:@378.4]
  wire  _T_1812; // @[Switch.scala 30:53:@380.4]
  wire  valid_4_14; // @[Switch.scala 30:36:@381.4]
  wire  _T_1815; // @[Switch.scala 30:53:@383.4]
  wire  valid_4_15; // @[Switch.scala 30:36:@384.4]
  wire [3:0] _T_1833; // @[Mux.scala 31:69:@386.4]
  wire [3:0] _T_1834; // @[Mux.scala 31:69:@387.4]
  wire [3:0] _T_1835; // @[Mux.scala 31:69:@388.4]
  wire [3:0] _T_1836; // @[Mux.scala 31:69:@389.4]
  wire [3:0] _T_1837; // @[Mux.scala 31:69:@390.4]
  wire [3:0] _T_1838; // @[Mux.scala 31:69:@391.4]
  wire [3:0] _T_1839; // @[Mux.scala 31:69:@392.4]
  wire [3:0] _T_1840; // @[Mux.scala 31:69:@393.4]
  wire [3:0] _T_1841; // @[Mux.scala 31:69:@394.4]
  wire [3:0] _T_1842; // @[Mux.scala 31:69:@395.4]
  wire [3:0] _T_1843; // @[Mux.scala 31:69:@396.4]
  wire [3:0] _T_1844; // @[Mux.scala 31:69:@397.4]
  wire [3:0] _T_1845; // @[Mux.scala 31:69:@398.4]
  wire [3:0] _T_1846; // @[Mux.scala 31:69:@399.4]
  wire [3:0] select_4; // @[Mux.scala 31:69:@400.4]
  wire [47:0] _GEN_65; // @[Switch.scala 33:19:@402.4]
  wire [47:0] _GEN_66; // @[Switch.scala 33:19:@402.4]
  wire [47:0] _GEN_67; // @[Switch.scala 33:19:@402.4]
  wire [47:0] _GEN_68; // @[Switch.scala 33:19:@402.4]
  wire [47:0] _GEN_69; // @[Switch.scala 33:19:@402.4]
  wire [47:0] _GEN_70; // @[Switch.scala 33:19:@402.4]
  wire [47:0] _GEN_71; // @[Switch.scala 33:19:@402.4]
  wire [47:0] _GEN_72; // @[Switch.scala 33:19:@402.4]
  wire [47:0] _GEN_73; // @[Switch.scala 33:19:@402.4]
  wire [47:0] _GEN_74; // @[Switch.scala 33:19:@402.4]
  wire [47:0] _GEN_75; // @[Switch.scala 33:19:@402.4]
  wire [47:0] _GEN_76; // @[Switch.scala 33:19:@402.4]
  wire [47:0] _GEN_77; // @[Switch.scala 33:19:@402.4]
  wire [47:0] _GEN_78; // @[Switch.scala 33:19:@402.4]
  wire [7:0] _T_1855; // @[Switch.scala 34:32:@409.4]
  wire [15:0] _T_1863; // @[Switch.scala 34:32:@417.4]
  wire  _T_1867; // @[Switch.scala 30:53:@420.4]
  wire  valid_5_0; // @[Switch.scala 30:36:@421.4]
  wire  _T_1870; // @[Switch.scala 30:53:@423.4]
  wire  valid_5_1; // @[Switch.scala 30:36:@424.4]
  wire  _T_1873; // @[Switch.scala 30:53:@426.4]
  wire  valid_5_2; // @[Switch.scala 30:36:@427.4]
  wire  _T_1876; // @[Switch.scala 30:53:@429.4]
  wire  valid_5_3; // @[Switch.scala 30:36:@430.4]
  wire  _T_1879; // @[Switch.scala 30:53:@432.4]
  wire  valid_5_4; // @[Switch.scala 30:36:@433.4]
  wire  _T_1882; // @[Switch.scala 30:53:@435.4]
  wire  valid_5_5; // @[Switch.scala 30:36:@436.4]
  wire  _T_1885; // @[Switch.scala 30:53:@438.4]
  wire  valid_5_6; // @[Switch.scala 30:36:@439.4]
  wire  _T_1888; // @[Switch.scala 30:53:@441.4]
  wire  valid_5_7; // @[Switch.scala 30:36:@442.4]
  wire  _T_1891; // @[Switch.scala 30:53:@444.4]
  wire  valid_5_8; // @[Switch.scala 30:36:@445.4]
  wire  _T_1894; // @[Switch.scala 30:53:@447.4]
  wire  valid_5_9; // @[Switch.scala 30:36:@448.4]
  wire  _T_1897; // @[Switch.scala 30:53:@450.4]
  wire  valid_5_10; // @[Switch.scala 30:36:@451.4]
  wire  _T_1900; // @[Switch.scala 30:53:@453.4]
  wire  valid_5_11; // @[Switch.scala 30:36:@454.4]
  wire  _T_1903; // @[Switch.scala 30:53:@456.4]
  wire  valid_5_12; // @[Switch.scala 30:36:@457.4]
  wire  _T_1906; // @[Switch.scala 30:53:@459.4]
  wire  valid_5_13; // @[Switch.scala 30:36:@460.4]
  wire  _T_1909; // @[Switch.scala 30:53:@462.4]
  wire  valid_5_14; // @[Switch.scala 30:36:@463.4]
  wire  _T_1912; // @[Switch.scala 30:53:@465.4]
  wire  valid_5_15; // @[Switch.scala 30:36:@466.4]
  wire [3:0] _T_1930; // @[Mux.scala 31:69:@468.4]
  wire [3:0] _T_1931; // @[Mux.scala 31:69:@469.4]
  wire [3:0] _T_1932; // @[Mux.scala 31:69:@470.4]
  wire [3:0] _T_1933; // @[Mux.scala 31:69:@471.4]
  wire [3:0] _T_1934; // @[Mux.scala 31:69:@472.4]
  wire [3:0] _T_1935; // @[Mux.scala 31:69:@473.4]
  wire [3:0] _T_1936; // @[Mux.scala 31:69:@474.4]
  wire [3:0] _T_1937; // @[Mux.scala 31:69:@475.4]
  wire [3:0] _T_1938; // @[Mux.scala 31:69:@476.4]
  wire [3:0] _T_1939; // @[Mux.scala 31:69:@477.4]
  wire [3:0] _T_1940; // @[Mux.scala 31:69:@478.4]
  wire [3:0] _T_1941; // @[Mux.scala 31:69:@479.4]
  wire [3:0] _T_1942; // @[Mux.scala 31:69:@480.4]
  wire [3:0] _T_1943; // @[Mux.scala 31:69:@481.4]
  wire [3:0] select_5; // @[Mux.scala 31:69:@482.4]
  wire [47:0] _GEN_81; // @[Switch.scala 33:19:@484.4]
  wire [47:0] _GEN_82; // @[Switch.scala 33:19:@484.4]
  wire [47:0] _GEN_83; // @[Switch.scala 33:19:@484.4]
  wire [47:0] _GEN_84; // @[Switch.scala 33:19:@484.4]
  wire [47:0] _GEN_85; // @[Switch.scala 33:19:@484.4]
  wire [47:0] _GEN_86; // @[Switch.scala 33:19:@484.4]
  wire [47:0] _GEN_87; // @[Switch.scala 33:19:@484.4]
  wire [47:0] _GEN_88; // @[Switch.scala 33:19:@484.4]
  wire [47:0] _GEN_89; // @[Switch.scala 33:19:@484.4]
  wire [47:0] _GEN_90; // @[Switch.scala 33:19:@484.4]
  wire [47:0] _GEN_91; // @[Switch.scala 33:19:@484.4]
  wire [47:0] _GEN_92; // @[Switch.scala 33:19:@484.4]
  wire [47:0] _GEN_93; // @[Switch.scala 33:19:@484.4]
  wire [47:0] _GEN_94; // @[Switch.scala 33:19:@484.4]
  wire [7:0] _T_1952; // @[Switch.scala 34:32:@491.4]
  wire [15:0] _T_1960; // @[Switch.scala 34:32:@499.4]
  wire  _T_1964; // @[Switch.scala 30:53:@502.4]
  wire  valid_6_0; // @[Switch.scala 30:36:@503.4]
  wire  _T_1967; // @[Switch.scala 30:53:@505.4]
  wire  valid_6_1; // @[Switch.scala 30:36:@506.4]
  wire  _T_1970; // @[Switch.scala 30:53:@508.4]
  wire  valid_6_2; // @[Switch.scala 30:36:@509.4]
  wire  _T_1973; // @[Switch.scala 30:53:@511.4]
  wire  valid_6_3; // @[Switch.scala 30:36:@512.4]
  wire  _T_1976; // @[Switch.scala 30:53:@514.4]
  wire  valid_6_4; // @[Switch.scala 30:36:@515.4]
  wire  _T_1979; // @[Switch.scala 30:53:@517.4]
  wire  valid_6_5; // @[Switch.scala 30:36:@518.4]
  wire  _T_1982; // @[Switch.scala 30:53:@520.4]
  wire  valid_6_6; // @[Switch.scala 30:36:@521.4]
  wire  _T_1985; // @[Switch.scala 30:53:@523.4]
  wire  valid_6_7; // @[Switch.scala 30:36:@524.4]
  wire  _T_1988; // @[Switch.scala 30:53:@526.4]
  wire  valid_6_8; // @[Switch.scala 30:36:@527.4]
  wire  _T_1991; // @[Switch.scala 30:53:@529.4]
  wire  valid_6_9; // @[Switch.scala 30:36:@530.4]
  wire  _T_1994; // @[Switch.scala 30:53:@532.4]
  wire  valid_6_10; // @[Switch.scala 30:36:@533.4]
  wire  _T_1997; // @[Switch.scala 30:53:@535.4]
  wire  valid_6_11; // @[Switch.scala 30:36:@536.4]
  wire  _T_2000; // @[Switch.scala 30:53:@538.4]
  wire  valid_6_12; // @[Switch.scala 30:36:@539.4]
  wire  _T_2003; // @[Switch.scala 30:53:@541.4]
  wire  valid_6_13; // @[Switch.scala 30:36:@542.4]
  wire  _T_2006; // @[Switch.scala 30:53:@544.4]
  wire  valid_6_14; // @[Switch.scala 30:36:@545.4]
  wire  _T_2009; // @[Switch.scala 30:53:@547.4]
  wire  valid_6_15; // @[Switch.scala 30:36:@548.4]
  wire [3:0] _T_2027; // @[Mux.scala 31:69:@550.4]
  wire [3:0] _T_2028; // @[Mux.scala 31:69:@551.4]
  wire [3:0] _T_2029; // @[Mux.scala 31:69:@552.4]
  wire [3:0] _T_2030; // @[Mux.scala 31:69:@553.4]
  wire [3:0] _T_2031; // @[Mux.scala 31:69:@554.4]
  wire [3:0] _T_2032; // @[Mux.scala 31:69:@555.4]
  wire [3:0] _T_2033; // @[Mux.scala 31:69:@556.4]
  wire [3:0] _T_2034; // @[Mux.scala 31:69:@557.4]
  wire [3:0] _T_2035; // @[Mux.scala 31:69:@558.4]
  wire [3:0] _T_2036; // @[Mux.scala 31:69:@559.4]
  wire [3:0] _T_2037; // @[Mux.scala 31:69:@560.4]
  wire [3:0] _T_2038; // @[Mux.scala 31:69:@561.4]
  wire [3:0] _T_2039; // @[Mux.scala 31:69:@562.4]
  wire [3:0] _T_2040; // @[Mux.scala 31:69:@563.4]
  wire [3:0] select_6; // @[Mux.scala 31:69:@564.4]
  wire [47:0] _GEN_97; // @[Switch.scala 33:19:@566.4]
  wire [47:0] _GEN_98; // @[Switch.scala 33:19:@566.4]
  wire [47:0] _GEN_99; // @[Switch.scala 33:19:@566.4]
  wire [47:0] _GEN_100; // @[Switch.scala 33:19:@566.4]
  wire [47:0] _GEN_101; // @[Switch.scala 33:19:@566.4]
  wire [47:0] _GEN_102; // @[Switch.scala 33:19:@566.4]
  wire [47:0] _GEN_103; // @[Switch.scala 33:19:@566.4]
  wire [47:0] _GEN_104; // @[Switch.scala 33:19:@566.4]
  wire [47:0] _GEN_105; // @[Switch.scala 33:19:@566.4]
  wire [47:0] _GEN_106; // @[Switch.scala 33:19:@566.4]
  wire [47:0] _GEN_107; // @[Switch.scala 33:19:@566.4]
  wire [47:0] _GEN_108; // @[Switch.scala 33:19:@566.4]
  wire [47:0] _GEN_109; // @[Switch.scala 33:19:@566.4]
  wire [47:0] _GEN_110; // @[Switch.scala 33:19:@566.4]
  wire [7:0] _T_2049; // @[Switch.scala 34:32:@573.4]
  wire [15:0] _T_2057; // @[Switch.scala 34:32:@581.4]
  wire  _T_2061; // @[Switch.scala 30:53:@584.4]
  wire  valid_7_0; // @[Switch.scala 30:36:@585.4]
  wire  _T_2064; // @[Switch.scala 30:53:@587.4]
  wire  valid_7_1; // @[Switch.scala 30:36:@588.4]
  wire  _T_2067; // @[Switch.scala 30:53:@590.4]
  wire  valid_7_2; // @[Switch.scala 30:36:@591.4]
  wire  _T_2070; // @[Switch.scala 30:53:@593.4]
  wire  valid_7_3; // @[Switch.scala 30:36:@594.4]
  wire  _T_2073; // @[Switch.scala 30:53:@596.4]
  wire  valid_7_4; // @[Switch.scala 30:36:@597.4]
  wire  _T_2076; // @[Switch.scala 30:53:@599.4]
  wire  valid_7_5; // @[Switch.scala 30:36:@600.4]
  wire  _T_2079; // @[Switch.scala 30:53:@602.4]
  wire  valid_7_6; // @[Switch.scala 30:36:@603.4]
  wire  _T_2082; // @[Switch.scala 30:53:@605.4]
  wire  valid_7_7; // @[Switch.scala 30:36:@606.4]
  wire  _T_2085; // @[Switch.scala 30:53:@608.4]
  wire  valid_7_8; // @[Switch.scala 30:36:@609.4]
  wire  _T_2088; // @[Switch.scala 30:53:@611.4]
  wire  valid_7_9; // @[Switch.scala 30:36:@612.4]
  wire  _T_2091; // @[Switch.scala 30:53:@614.4]
  wire  valid_7_10; // @[Switch.scala 30:36:@615.4]
  wire  _T_2094; // @[Switch.scala 30:53:@617.4]
  wire  valid_7_11; // @[Switch.scala 30:36:@618.4]
  wire  _T_2097; // @[Switch.scala 30:53:@620.4]
  wire  valid_7_12; // @[Switch.scala 30:36:@621.4]
  wire  _T_2100; // @[Switch.scala 30:53:@623.4]
  wire  valid_7_13; // @[Switch.scala 30:36:@624.4]
  wire  _T_2103; // @[Switch.scala 30:53:@626.4]
  wire  valid_7_14; // @[Switch.scala 30:36:@627.4]
  wire  _T_2106; // @[Switch.scala 30:53:@629.4]
  wire  valid_7_15; // @[Switch.scala 30:36:@630.4]
  wire [3:0] _T_2124; // @[Mux.scala 31:69:@632.4]
  wire [3:0] _T_2125; // @[Mux.scala 31:69:@633.4]
  wire [3:0] _T_2126; // @[Mux.scala 31:69:@634.4]
  wire [3:0] _T_2127; // @[Mux.scala 31:69:@635.4]
  wire [3:0] _T_2128; // @[Mux.scala 31:69:@636.4]
  wire [3:0] _T_2129; // @[Mux.scala 31:69:@637.4]
  wire [3:0] _T_2130; // @[Mux.scala 31:69:@638.4]
  wire [3:0] _T_2131; // @[Mux.scala 31:69:@639.4]
  wire [3:0] _T_2132; // @[Mux.scala 31:69:@640.4]
  wire [3:0] _T_2133; // @[Mux.scala 31:69:@641.4]
  wire [3:0] _T_2134; // @[Mux.scala 31:69:@642.4]
  wire [3:0] _T_2135; // @[Mux.scala 31:69:@643.4]
  wire [3:0] _T_2136; // @[Mux.scala 31:69:@644.4]
  wire [3:0] _T_2137; // @[Mux.scala 31:69:@645.4]
  wire [3:0] select_7; // @[Mux.scala 31:69:@646.4]
  wire [47:0] _GEN_113; // @[Switch.scala 33:19:@648.4]
  wire [47:0] _GEN_114; // @[Switch.scala 33:19:@648.4]
  wire [47:0] _GEN_115; // @[Switch.scala 33:19:@648.4]
  wire [47:0] _GEN_116; // @[Switch.scala 33:19:@648.4]
  wire [47:0] _GEN_117; // @[Switch.scala 33:19:@648.4]
  wire [47:0] _GEN_118; // @[Switch.scala 33:19:@648.4]
  wire [47:0] _GEN_119; // @[Switch.scala 33:19:@648.4]
  wire [47:0] _GEN_120; // @[Switch.scala 33:19:@648.4]
  wire [47:0] _GEN_121; // @[Switch.scala 33:19:@648.4]
  wire [47:0] _GEN_122; // @[Switch.scala 33:19:@648.4]
  wire [47:0] _GEN_123; // @[Switch.scala 33:19:@648.4]
  wire [47:0] _GEN_124; // @[Switch.scala 33:19:@648.4]
  wire [47:0] _GEN_125; // @[Switch.scala 33:19:@648.4]
  wire [47:0] _GEN_126; // @[Switch.scala 33:19:@648.4]
  wire [7:0] _T_2146; // @[Switch.scala 34:32:@655.4]
  wire [15:0] _T_2154; // @[Switch.scala 34:32:@663.4]
  wire  _T_2158; // @[Switch.scala 30:53:@666.4]
  wire  valid_8_0; // @[Switch.scala 30:36:@667.4]
  wire  _T_2161; // @[Switch.scala 30:53:@669.4]
  wire  valid_8_1; // @[Switch.scala 30:36:@670.4]
  wire  _T_2164; // @[Switch.scala 30:53:@672.4]
  wire  valid_8_2; // @[Switch.scala 30:36:@673.4]
  wire  _T_2167; // @[Switch.scala 30:53:@675.4]
  wire  valid_8_3; // @[Switch.scala 30:36:@676.4]
  wire  _T_2170; // @[Switch.scala 30:53:@678.4]
  wire  valid_8_4; // @[Switch.scala 30:36:@679.4]
  wire  _T_2173; // @[Switch.scala 30:53:@681.4]
  wire  valid_8_5; // @[Switch.scala 30:36:@682.4]
  wire  _T_2176; // @[Switch.scala 30:53:@684.4]
  wire  valid_8_6; // @[Switch.scala 30:36:@685.4]
  wire  _T_2179; // @[Switch.scala 30:53:@687.4]
  wire  valid_8_7; // @[Switch.scala 30:36:@688.4]
  wire  _T_2182; // @[Switch.scala 30:53:@690.4]
  wire  valid_8_8; // @[Switch.scala 30:36:@691.4]
  wire  _T_2185; // @[Switch.scala 30:53:@693.4]
  wire  valid_8_9; // @[Switch.scala 30:36:@694.4]
  wire  _T_2188; // @[Switch.scala 30:53:@696.4]
  wire  valid_8_10; // @[Switch.scala 30:36:@697.4]
  wire  _T_2191; // @[Switch.scala 30:53:@699.4]
  wire  valid_8_11; // @[Switch.scala 30:36:@700.4]
  wire  _T_2194; // @[Switch.scala 30:53:@702.4]
  wire  valid_8_12; // @[Switch.scala 30:36:@703.4]
  wire  _T_2197; // @[Switch.scala 30:53:@705.4]
  wire  valid_8_13; // @[Switch.scala 30:36:@706.4]
  wire  _T_2200; // @[Switch.scala 30:53:@708.4]
  wire  valid_8_14; // @[Switch.scala 30:36:@709.4]
  wire  _T_2203; // @[Switch.scala 30:53:@711.4]
  wire  valid_8_15; // @[Switch.scala 30:36:@712.4]
  wire [3:0] _T_2221; // @[Mux.scala 31:69:@714.4]
  wire [3:0] _T_2222; // @[Mux.scala 31:69:@715.4]
  wire [3:0] _T_2223; // @[Mux.scala 31:69:@716.4]
  wire [3:0] _T_2224; // @[Mux.scala 31:69:@717.4]
  wire [3:0] _T_2225; // @[Mux.scala 31:69:@718.4]
  wire [3:0] _T_2226; // @[Mux.scala 31:69:@719.4]
  wire [3:0] _T_2227; // @[Mux.scala 31:69:@720.4]
  wire [3:0] _T_2228; // @[Mux.scala 31:69:@721.4]
  wire [3:0] _T_2229; // @[Mux.scala 31:69:@722.4]
  wire [3:0] _T_2230; // @[Mux.scala 31:69:@723.4]
  wire [3:0] _T_2231; // @[Mux.scala 31:69:@724.4]
  wire [3:0] _T_2232; // @[Mux.scala 31:69:@725.4]
  wire [3:0] _T_2233; // @[Mux.scala 31:69:@726.4]
  wire [3:0] _T_2234; // @[Mux.scala 31:69:@727.4]
  wire [3:0] select_8; // @[Mux.scala 31:69:@728.4]
  wire [47:0] _GEN_129; // @[Switch.scala 33:19:@730.4]
  wire [47:0] _GEN_130; // @[Switch.scala 33:19:@730.4]
  wire [47:0] _GEN_131; // @[Switch.scala 33:19:@730.4]
  wire [47:0] _GEN_132; // @[Switch.scala 33:19:@730.4]
  wire [47:0] _GEN_133; // @[Switch.scala 33:19:@730.4]
  wire [47:0] _GEN_134; // @[Switch.scala 33:19:@730.4]
  wire [47:0] _GEN_135; // @[Switch.scala 33:19:@730.4]
  wire [47:0] _GEN_136; // @[Switch.scala 33:19:@730.4]
  wire [47:0] _GEN_137; // @[Switch.scala 33:19:@730.4]
  wire [47:0] _GEN_138; // @[Switch.scala 33:19:@730.4]
  wire [47:0] _GEN_139; // @[Switch.scala 33:19:@730.4]
  wire [47:0] _GEN_140; // @[Switch.scala 33:19:@730.4]
  wire [47:0] _GEN_141; // @[Switch.scala 33:19:@730.4]
  wire [47:0] _GEN_142; // @[Switch.scala 33:19:@730.4]
  wire [7:0] _T_2243; // @[Switch.scala 34:32:@737.4]
  wire [15:0] _T_2251; // @[Switch.scala 34:32:@745.4]
  wire  _T_2255; // @[Switch.scala 30:53:@748.4]
  wire  valid_9_0; // @[Switch.scala 30:36:@749.4]
  wire  _T_2258; // @[Switch.scala 30:53:@751.4]
  wire  valid_9_1; // @[Switch.scala 30:36:@752.4]
  wire  _T_2261; // @[Switch.scala 30:53:@754.4]
  wire  valid_9_2; // @[Switch.scala 30:36:@755.4]
  wire  _T_2264; // @[Switch.scala 30:53:@757.4]
  wire  valid_9_3; // @[Switch.scala 30:36:@758.4]
  wire  _T_2267; // @[Switch.scala 30:53:@760.4]
  wire  valid_9_4; // @[Switch.scala 30:36:@761.4]
  wire  _T_2270; // @[Switch.scala 30:53:@763.4]
  wire  valid_9_5; // @[Switch.scala 30:36:@764.4]
  wire  _T_2273; // @[Switch.scala 30:53:@766.4]
  wire  valid_9_6; // @[Switch.scala 30:36:@767.4]
  wire  _T_2276; // @[Switch.scala 30:53:@769.4]
  wire  valid_9_7; // @[Switch.scala 30:36:@770.4]
  wire  _T_2279; // @[Switch.scala 30:53:@772.4]
  wire  valid_9_8; // @[Switch.scala 30:36:@773.4]
  wire  _T_2282; // @[Switch.scala 30:53:@775.4]
  wire  valid_9_9; // @[Switch.scala 30:36:@776.4]
  wire  _T_2285; // @[Switch.scala 30:53:@778.4]
  wire  valid_9_10; // @[Switch.scala 30:36:@779.4]
  wire  _T_2288; // @[Switch.scala 30:53:@781.4]
  wire  valid_9_11; // @[Switch.scala 30:36:@782.4]
  wire  _T_2291; // @[Switch.scala 30:53:@784.4]
  wire  valid_9_12; // @[Switch.scala 30:36:@785.4]
  wire  _T_2294; // @[Switch.scala 30:53:@787.4]
  wire  valid_9_13; // @[Switch.scala 30:36:@788.4]
  wire  _T_2297; // @[Switch.scala 30:53:@790.4]
  wire  valid_9_14; // @[Switch.scala 30:36:@791.4]
  wire  _T_2300; // @[Switch.scala 30:53:@793.4]
  wire  valid_9_15; // @[Switch.scala 30:36:@794.4]
  wire [3:0] _T_2318; // @[Mux.scala 31:69:@796.4]
  wire [3:0] _T_2319; // @[Mux.scala 31:69:@797.4]
  wire [3:0] _T_2320; // @[Mux.scala 31:69:@798.4]
  wire [3:0] _T_2321; // @[Mux.scala 31:69:@799.4]
  wire [3:0] _T_2322; // @[Mux.scala 31:69:@800.4]
  wire [3:0] _T_2323; // @[Mux.scala 31:69:@801.4]
  wire [3:0] _T_2324; // @[Mux.scala 31:69:@802.4]
  wire [3:0] _T_2325; // @[Mux.scala 31:69:@803.4]
  wire [3:0] _T_2326; // @[Mux.scala 31:69:@804.4]
  wire [3:0] _T_2327; // @[Mux.scala 31:69:@805.4]
  wire [3:0] _T_2328; // @[Mux.scala 31:69:@806.4]
  wire [3:0] _T_2329; // @[Mux.scala 31:69:@807.4]
  wire [3:0] _T_2330; // @[Mux.scala 31:69:@808.4]
  wire [3:0] _T_2331; // @[Mux.scala 31:69:@809.4]
  wire [3:0] select_9; // @[Mux.scala 31:69:@810.4]
  wire [47:0] _GEN_145; // @[Switch.scala 33:19:@812.4]
  wire [47:0] _GEN_146; // @[Switch.scala 33:19:@812.4]
  wire [47:0] _GEN_147; // @[Switch.scala 33:19:@812.4]
  wire [47:0] _GEN_148; // @[Switch.scala 33:19:@812.4]
  wire [47:0] _GEN_149; // @[Switch.scala 33:19:@812.4]
  wire [47:0] _GEN_150; // @[Switch.scala 33:19:@812.4]
  wire [47:0] _GEN_151; // @[Switch.scala 33:19:@812.4]
  wire [47:0] _GEN_152; // @[Switch.scala 33:19:@812.4]
  wire [47:0] _GEN_153; // @[Switch.scala 33:19:@812.4]
  wire [47:0] _GEN_154; // @[Switch.scala 33:19:@812.4]
  wire [47:0] _GEN_155; // @[Switch.scala 33:19:@812.4]
  wire [47:0] _GEN_156; // @[Switch.scala 33:19:@812.4]
  wire [47:0] _GEN_157; // @[Switch.scala 33:19:@812.4]
  wire [47:0] _GEN_158; // @[Switch.scala 33:19:@812.4]
  wire [7:0] _T_2340; // @[Switch.scala 34:32:@819.4]
  wire [15:0] _T_2348; // @[Switch.scala 34:32:@827.4]
  wire  _T_2352; // @[Switch.scala 30:53:@830.4]
  wire  valid_10_0; // @[Switch.scala 30:36:@831.4]
  wire  _T_2355; // @[Switch.scala 30:53:@833.4]
  wire  valid_10_1; // @[Switch.scala 30:36:@834.4]
  wire  _T_2358; // @[Switch.scala 30:53:@836.4]
  wire  valid_10_2; // @[Switch.scala 30:36:@837.4]
  wire  _T_2361; // @[Switch.scala 30:53:@839.4]
  wire  valid_10_3; // @[Switch.scala 30:36:@840.4]
  wire  _T_2364; // @[Switch.scala 30:53:@842.4]
  wire  valid_10_4; // @[Switch.scala 30:36:@843.4]
  wire  _T_2367; // @[Switch.scala 30:53:@845.4]
  wire  valid_10_5; // @[Switch.scala 30:36:@846.4]
  wire  _T_2370; // @[Switch.scala 30:53:@848.4]
  wire  valid_10_6; // @[Switch.scala 30:36:@849.4]
  wire  _T_2373; // @[Switch.scala 30:53:@851.4]
  wire  valid_10_7; // @[Switch.scala 30:36:@852.4]
  wire  _T_2376; // @[Switch.scala 30:53:@854.4]
  wire  valid_10_8; // @[Switch.scala 30:36:@855.4]
  wire  _T_2379; // @[Switch.scala 30:53:@857.4]
  wire  valid_10_9; // @[Switch.scala 30:36:@858.4]
  wire  _T_2382; // @[Switch.scala 30:53:@860.4]
  wire  valid_10_10; // @[Switch.scala 30:36:@861.4]
  wire  _T_2385; // @[Switch.scala 30:53:@863.4]
  wire  valid_10_11; // @[Switch.scala 30:36:@864.4]
  wire  _T_2388; // @[Switch.scala 30:53:@866.4]
  wire  valid_10_12; // @[Switch.scala 30:36:@867.4]
  wire  _T_2391; // @[Switch.scala 30:53:@869.4]
  wire  valid_10_13; // @[Switch.scala 30:36:@870.4]
  wire  _T_2394; // @[Switch.scala 30:53:@872.4]
  wire  valid_10_14; // @[Switch.scala 30:36:@873.4]
  wire  _T_2397; // @[Switch.scala 30:53:@875.4]
  wire  valid_10_15; // @[Switch.scala 30:36:@876.4]
  wire [3:0] _T_2415; // @[Mux.scala 31:69:@878.4]
  wire [3:0] _T_2416; // @[Mux.scala 31:69:@879.4]
  wire [3:0] _T_2417; // @[Mux.scala 31:69:@880.4]
  wire [3:0] _T_2418; // @[Mux.scala 31:69:@881.4]
  wire [3:0] _T_2419; // @[Mux.scala 31:69:@882.4]
  wire [3:0] _T_2420; // @[Mux.scala 31:69:@883.4]
  wire [3:0] _T_2421; // @[Mux.scala 31:69:@884.4]
  wire [3:0] _T_2422; // @[Mux.scala 31:69:@885.4]
  wire [3:0] _T_2423; // @[Mux.scala 31:69:@886.4]
  wire [3:0] _T_2424; // @[Mux.scala 31:69:@887.4]
  wire [3:0] _T_2425; // @[Mux.scala 31:69:@888.4]
  wire [3:0] _T_2426; // @[Mux.scala 31:69:@889.4]
  wire [3:0] _T_2427; // @[Mux.scala 31:69:@890.4]
  wire [3:0] _T_2428; // @[Mux.scala 31:69:@891.4]
  wire [3:0] select_10; // @[Mux.scala 31:69:@892.4]
  wire [47:0] _GEN_161; // @[Switch.scala 33:19:@894.4]
  wire [47:0] _GEN_162; // @[Switch.scala 33:19:@894.4]
  wire [47:0] _GEN_163; // @[Switch.scala 33:19:@894.4]
  wire [47:0] _GEN_164; // @[Switch.scala 33:19:@894.4]
  wire [47:0] _GEN_165; // @[Switch.scala 33:19:@894.4]
  wire [47:0] _GEN_166; // @[Switch.scala 33:19:@894.4]
  wire [47:0] _GEN_167; // @[Switch.scala 33:19:@894.4]
  wire [47:0] _GEN_168; // @[Switch.scala 33:19:@894.4]
  wire [47:0] _GEN_169; // @[Switch.scala 33:19:@894.4]
  wire [47:0] _GEN_170; // @[Switch.scala 33:19:@894.4]
  wire [47:0] _GEN_171; // @[Switch.scala 33:19:@894.4]
  wire [47:0] _GEN_172; // @[Switch.scala 33:19:@894.4]
  wire [47:0] _GEN_173; // @[Switch.scala 33:19:@894.4]
  wire [47:0] _GEN_174; // @[Switch.scala 33:19:@894.4]
  wire [7:0] _T_2437; // @[Switch.scala 34:32:@901.4]
  wire [15:0] _T_2445; // @[Switch.scala 34:32:@909.4]
  wire  _T_2449; // @[Switch.scala 30:53:@912.4]
  wire  valid_11_0; // @[Switch.scala 30:36:@913.4]
  wire  _T_2452; // @[Switch.scala 30:53:@915.4]
  wire  valid_11_1; // @[Switch.scala 30:36:@916.4]
  wire  _T_2455; // @[Switch.scala 30:53:@918.4]
  wire  valid_11_2; // @[Switch.scala 30:36:@919.4]
  wire  _T_2458; // @[Switch.scala 30:53:@921.4]
  wire  valid_11_3; // @[Switch.scala 30:36:@922.4]
  wire  _T_2461; // @[Switch.scala 30:53:@924.4]
  wire  valid_11_4; // @[Switch.scala 30:36:@925.4]
  wire  _T_2464; // @[Switch.scala 30:53:@927.4]
  wire  valid_11_5; // @[Switch.scala 30:36:@928.4]
  wire  _T_2467; // @[Switch.scala 30:53:@930.4]
  wire  valid_11_6; // @[Switch.scala 30:36:@931.4]
  wire  _T_2470; // @[Switch.scala 30:53:@933.4]
  wire  valid_11_7; // @[Switch.scala 30:36:@934.4]
  wire  _T_2473; // @[Switch.scala 30:53:@936.4]
  wire  valid_11_8; // @[Switch.scala 30:36:@937.4]
  wire  _T_2476; // @[Switch.scala 30:53:@939.4]
  wire  valid_11_9; // @[Switch.scala 30:36:@940.4]
  wire  _T_2479; // @[Switch.scala 30:53:@942.4]
  wire  valid_11_10; // @[Switch.scala 30:36:@943.4]
  wire  _T_2482; // @[Switch.scala 30:53:@945.4]
  wire  valid_11_11; // @[Switch.scala 30:36:@946.4]
  wire  _T_2485; // @[Switch.scala 30:53:@948.4]
  wire  valid_11_12; // @[Switch.scala 30:36:@949.4]
  wire  _T_2488; // @[Switch.scala 30:53:@951.4]
  wire  valid_11_13; // @[Switch.scala 30:36:@952.4]
  wire  _T_2491; // @[Switch.scala 30:53:@954.4]
  wire  valid_11_14; // @[Switch.scala 30:36:@955.4]
  wire  _T_2494; // @[Switch.scala 30:53:@957.4]
  wire  valid_11_15; // @[Switch.scala 30:36:@958.4]
  wire [3:0] _T_2512; // @[Mux.scala 31:69:@960.4]
  wire [3:0] _T_2513; // @[Mux.scala 31:69:@961.4]
  wire [3:0] _T_2514; // @[Mux.scala 31:69:@962.4]
  wire [3:0] _T_2515; // @[Mux.scala 31:69:@963.4]
  wire [3:0] _T_2516; // @[Mux.scala 31:69:@964.4]
  wire [3:0] _T_2517; // @[Mux.scala 31:69:@965.4]
  wire [3:0] _T_2518; // @[Mux.scala 31:69:@966.4]
  wire [3:0] _T_2519; // @[Mux.scala 31:69:@967.4]
  wire [3:0] _T_2520; // @[Mux.scala 31:69:@968.4]
  wire [3:0] _T_2521; // @[Mux.scala 31:69:@969.4]
  wire [3:0] _T_2522; // @[Mux.scala 31:69:@970.4]
  wire [3:0] _T_2523; // @[Mux.scala 31:69:@971.4]
  wire [3:0] _T_2524; // @[Mux.scala 31:69:@972.4]
  wire [3:0] _T_2525; // @[Mux.scala 31:69:@973.4]
  wire [3:0] select_11; // @[Mux.scala 31:69:@974.4]
  wire [47:0] _GEN_177; // @[Switch.scala 33:19:@976.4]
  wire [47:0] _GEN_178; // @[Switch.scala 33:19:@976.4]
  wire [47:0] _GEN_179; // @[Switch.scala 33:19:@976.4]
  wire [47:0] _GEN_180; // @[Switch.scala 33:19:@976.4]
  wire [47:0] _GEN_181; // @[Switch.scala 33:19:@976.4]
  wire [47:0] _GEN_182; // @[Switch.scala 33:19:@976.4]
  wire [47:0] _GEN_183; // @[Switch.scala 33:19:@976.4]
  wire [47:0] _GEN_184; // @[Switch.scala 33:19:@976.4]
  wire [47:0] _GEN_185; // @[Switch.scala 33:19:@976.4]
  wire [47:0] _GEN_186; // @[Switch.scala 33:19:@976.4]
  wire [47:0] _GEN_187; // @[Switch.scala 33:19:@976.4]
  wire [47:0] _GEN_188; // @[Switch.scala 33:19:@976.4]
  wire [47:0] _GEN_189; // @[Switch.scala 33:19:@976.4]
  wire [47:0] _GEN_190; // @[Switch.scala 33:19:@976.4]
  wire [7:0] _T_2534; // @[Switch.scala 34:32:@983.4]
  wire [15:0] _T_2542; // @[Switch.scala 34:32:@991.4]
  wire  _T_2546; // @[Switch.scala 30:53:@994.4]
  wire  valid_12_0; // @[Switch.scala 30:36:@995.4]
  wire  _T_2549; // @[Switch.scala 30:53:@997.4]
  wire  valid_12_1; // @[Switch.scala 30:36:@998.4]
  wire  _T_2552; // @[Switch.scala 30:53:@1000.4]
  wire  valid_12_2; // @[Switch.scala 30:36:@1001.4]
  wire  _T_2555; // @[Switch.scala 30:53:@1003.4]
  wire  valid_12_3; // @[Switch.scala 30:36:@1004.4]
  wire  _T_2558; // @[Switch.scala 30:53:@1006.4]
  wire  valid_12_4; // @[Switch.scala 30:36:@1007.4]
  wire  _T_2561; // @[Switch.scala 30:53:@1009.4]
  wire  valid_12_5; // @[Switch.scala 30:36:@1010.4]
  wire  _T_2564; // @[Switch.scala 30:53:@1012.4]
  wire  valid_12_6; // @[Switch.scala 30:36:@1013.4]
  wire  _T_2567; // @[Switch.scala 30:53:@1015.4]
  wire  valid_12_7; // @[Switch.scala 30:36:@1016.4]
  wire  _T_2570; // @[Switch.scala 30:53:@1018.4]
  wire  valid_12_8; // @[Switch.scala 30:36:@1019.4]
  wire  _T_2573; // @[Switch.scala 30:53:@1021.4]
  wire  valid_12_9; // @[Switch.scala 30:36:@1022.4]
  wire  _T_2576; // @[Switch.scala 30:53:@1024.4]
  wire  valid_12_10; // @[Switch.scala 30:36:@1025.4]
  wire  _T_2579; // @[Switch.scala 30:53:@1027.4]
  wire  valid_12_11; // @[Switch.scala 30:36:@1028.4]
  wire  _T_2582; // @[Switch.scala 30:53:@1030.4]
  wire  valid_12_12; // @[Switch.scala 30:36:@1031.4]
  wire  _T_2585; // @[Switch.scala 30:53:@1033.4]
  wire  valid_12_13; // @[Switch.scala 30:36:@1034.4]
  wire  _T_2588; // @[Switch.scala 30:53:@1036.4]
  wire  valid_12_14; // @[Switch.scala 30:36:@1037.4]
  wire  _T_2591; // @[Switch.scala 30:53:@1039.4]
  wire  valid_12_15; // @[Switch.scala 30:36:@1040.4]
  wire [3:0] _T_2609; // @[Mux.scala 31:69:@1042.4]
  wire [3:0] _T_2610; // @[Mux.scala 31:69:@1043.4]
  wire [3:0] _T_2611; // @[Mux.scala 31:69:@1044.4]
  wire [3:0] _T_2612; // @[Mux.scala 31:69:@1045.4]
  wire [3:0] _T_2613; // @[Mux.scala 31:69:@1046.4]
  wire [3:0] _T_2614; // @[Mux.scala 31:69:@1047.4]
  wire [3:0] _T_2615; // @[Mux.scala 31:69:@1048.4]
  wire [3:0] _T_2616; // @[Mux.scala 31:69:@1049.4]
  wire [3:0] _T_2617; // @[Mux.scala 31:69:@1050.4]
  wire [3:0] _T_2618; // @[Mux.scala 31:69:@1051.4]
  wire [3:0] _T_2619; // @[Mux.scala 31:69:@1052.4]
  wire [3:0] _T_2620; // @[Mux.scala 31:69:@1053.4]
  wire [3:0] _T_2621; // @[Mux.scala 31:69:@1054.4]
  wire [3:0] _T_2622; // @[Mux.scala 31:69:@1055.4]
  wire [3:0] select_12; // @[Mux.scala 31:69:@1056.4]
  wire [47:0] _GEN_193; // @[Switch.scala 33:19:@1058.4]
  wire [47:0] _GEN_194; // @[Switch.scala 33:19:@1058.4]
  wire [47:0] _GEN_195; // @[Switch.scala 33:19:@1058.4]
  wire [47:0] _GEN_196; // @[Switch.scala 33:19:@1058.4]
  wire [47:0] _GEN_197; // @[Switch.scala 33:19:@1058.4]
  wire [47:0] _GEN_198; // @[Switch.scala 33:19:@1058.4]
  wire [47:0] _GEN_199; // @[Switch.scala 33:19:@1058.4]
  wire [47:0] _GEN_200; // @[Switch.scala 33:19:@1058.4]
  wire [47:0] _GEN_201; // @[Switch.scala 33:19:@1058.4]
  wire [47:0] _GEN_202; // @[Switch.scala 33:19:@1058.4]
  wire [47:0] _GEN_203; // @[Switch.scala 33:19:@1058.4]
  wire [47:0] _GEN_204; // @[Switch.scala 33:19:@1058.4]
  wire [47:0] _GEN_205; // @[Switch.scala 33:19:@1058.4]
  wire [47:0] _GEN_206; // @[Switch.scala 33:19:@1058.4]
  wire [7:0] _T_2631; // @[Switch.scala 34:32:@1065.4]
  wire [15:0] _T_2639; // @[Switch.scala 34:32:@1073.4]
  wire  _T_2643; // @[Switch.scala 30:53:@1076.4]
  wire  valid_13_0; // @[Switch.scala 30:36:@1077.4]
  wire  _T_2646; // @[Switch.scala 30:53:@1079.4]
  wire  valid_13_1; // @[Switch.scala 30:36:@1080.4]
  wire  _T_2649; // @[Switch.scala 30:53:@1082.4]
  wire  valid_13_2; // @[Switch.scala 30:36:@1083.4]
  wire  _T_2652; // @[Switch.scala 30:53:@1085.4]
  wire  valid_13_3; // @[Switch.scala 30:36:@1086.4]
  wire  _T_2655; // @[Switch.scala 30:53:@1088.4]
  wire  valid_13_4; // @[Switch.scala 30:36:@1089.4]
  wire  _T_2658; // @[Switch.scala 30:53:@1091.4]
  wire  valid_13_5; // @[Switch.scala 30:36:@1092.4]
  wire  _T_2661; // @[Switch.scala 30:53:@1094.4]
  wire  valid_13_6; // @[Switch.scala 30:36:@1095.4]
  wire  _T_2664; // @[Switch.scala 30:53:@1097.4]
  wire  valid_13_7; // @[Switch.scala 30:36:@1098.4]
  wire  _T_2667; // @[Switch.scala 30:53:@1100.4]
  wire  valid_13_8; // @[Switch.scala 30:36:@1101.4]
  wire  _T_2670; // @[Switch.scala 30:53:@1103.4]
  wire  valid_13_9; // @[Switch.scala 30:36:@1104.4]
  wire  _T_2673; // @[Switch.scala 30:53:@1106.4]
  wire  valid_13_10; // @[Switch.scala 30:36:@1107.4]
  wire  _T_2676; // @[Switch.scala 30:53:@1109.4]
  wire  valid_13_11; // @[Switch.scala 30:36:@1110.4]
  wire  _T_2679; // @[Switch.scala 30:53:@1112.4]
  wire  valid_13_12; // @[Switch.scala 30:36:@1113.4]
  wire  _T_2682; // @[Switch.scala 30:53:@1115.4]
  wire  valid_13_13; // @[Switch.scala 30:36:@1116.4]
  wire  _T_2685; // @[Switch.scala 30:53:@1118.4]
  wire  valid_13_14; // @[Switch.scala 30:36:@1119.4]
  wire  _T_2688; // @[Switch.scala 30:53:@1121.4]
  wire  valid_13_15; // @[Switch.scala 30:36:@1122.4]
  wire [3:0] _T_2706; // @[Mux.scala 31:69:@1124.4]
  wire [3:0] _T_2707; // @[Mux.scala 31:69:@1125.4]
  wire [3:0] _T_2708; // @[Mux.scala 31:69:@1126.4]
  wire [3:0] _T_2709; // @[Mux.scala 31:69:@1127.4]
  wire [3:0] _T_2710; // @[Mux.scala 31:69:@1128.4]
  wire [3:0] _T_2711; // @[Mux.scala 31:69:@1129.4]
  wire [3:0] _T_2712; // @[Mux.scala 31:69:@1130.4]
  wire [3:0] _T_2713; // @[Mux.scala 31:69:@1131.4]
  wire [3:0] _T_2714; // @[Mux.scala 31:69:@1132.4]
  wire [3:0] _T_2715; // @[Mux.scala 31:69:@1133.4]
  wire [3:0] _T_2716; // @[Mux.scala 31:69:@1134.4]
  wire [3:0] _T_2717; // @[Mux.scala 31:69:@1135.4]
  wire [3:0] _T_2718; // @[Mux.scala 31:69:@1136.4]
  wire [3:0] _T_2719; // @[Mux.scala 31:69:@1137.4]
  wire [3:0] select_13; // @[Mux.scala 31:69:@1138.4]
  wire [47:0] _GEN_209; // @[Switch.scala 33:19:@1140.4]
  wire [47:0] _GEN_210; // @[Switch.scala 33:19:@1140.4]
  wire [47:0] _GEN_211; // @[Switch.scala 33:19:@1140.4]
  wire [47:0] _GEN_212; // @[Switch.scala 33:19:@1140.4]
  wire [47:0] _GEN_213; // @[Switch.scala 33:19:@1140.4]
  wire [47:0] _GEN_214; // @[Switch.scala 33:19:@1140.4]
  wire [47:0] _GEN_215; // @[Switch.scala 33:19:@1140.4]
  wire [47:0] _GEN_216; // @[Switch.scala 33:19:@1140.4]
  wire [47:0] _GEN_217; // @[Switch.scala 33:19:@1140.4]
  wire [47:0] _GEN_218; // @[Switch.scala 33:19:@1140.4]
  wire [47:0] _GEN_219; // @[Switch.scala 33:19:@1140.4]
  wire [47:0] _GEN_220; // @[Switch.scala 33:19:@1140.4]
  wire [47:0] _GEN_221; // @[Switch.scala 33:19:@1140.4]
  wire [47:0] _GEN_222; // @[Switch.scala 33:19:@1140.4]
  wire [7:0] _T_2728; // @[Switch.scala 34:32:@1147.4]
  wire [15:0] _T_2736; // @[Switch.scala 34:32:@1155.4]
  wire  _T_2740; // @[Switch.scala 30:53:@1158.4]
  wire  valid_14_0; // @[Switch.scala 30:36:@1159.4]
  wire  _T_2743; // @[Switch.scala 30:53:@1161.4]
  wire  valid_14_1; // @[Switch.scala 30:36:@1162.4]
  wire  _T_2746; // @[Switch.scala 30:53:@1164.4]
  wire  valid_14_2; // @[Switch.scala 30:36:@1165.4]
  wire  _T_2749; // @[Switch.scala 30:53:@1167.4]
  wire  valid_14_3; // @[Switch.scala 30:36:@1168.4]
  wire  _T_2752; // @[Switch.scala 30:53:@1170.4]
  wire  valid_14_4; // @[Switch.scala 30:36:@1171.4]
  wire  _T_2755; // @[Switch.scala 30:53:@1173.4]
  wire  valid_14_5; // @[Switch.scala 30:36:@1174.4]
  wire  _T_2758; // @[Switch.scala 30:53:@1176.4]
  wire  valid_14_6; // @[Switch.scala 30:36:@1177.4]
  wire  _T_2761; // @[Switch.scala 30:53:@1179.4]
  wire  valid_14_7; // @[Switch.scala 30:36:@1180.4]
  wire  _T_2764; // @[Switch.scala 30:53:@1182.4]
  wire  valid_14_8; // @[Switch.scala 30:36:@1183.4]
  wire  _T_2767; // @[Switch.scala 30:53:@1185.4]
  wire  valid_14_9; // @[Switch.scala 30:36:@1186.4]
  wire  _T_2770; // @[Switch.scala 30:53:@1188.4]
  wire  valid_14_10; // @[Switch.scala 30:36:@1189.4]
  wire  _T_2773; // @[Switch.scala 30:53:@1191.4]
  wire  valid_14_11; // @[Switch.scala 30:36:@1192.4]
  wire  _T_2776; // @[Switch.scala 30:53:@1194.4]
  wire  valid_14_12; // @[Switch.scala 30:36:@1195.4]
  wire  _T_2779; // @[Switch.scala 30:53:@1197.4]
  wire  valid_14_13; // @[Switch.scala 30:36:@1198.4]
  wire  _T_2782; // @[Switch.scala 30:53:@1200.4]
  wire  valid_14_14; // @[Switch.scala 30:36:@1201.4]
  wire  _T_2785; // @[Switch.scala 30:53:@1203.4]
  wire  valid_14_15; // @[Switch.scala 30:36:@1204.4]
  wire [3:0] _T_2803; // @[Mux.scala 31:69:@1206.4]
  wire [3:0] _T_2804; // @[Mux.scala 31:69:@1207.4]
  wire [3:0] _T_2805; // @[Mux.scala 31:69:@1208.4]
  wire [3:0] _T_2806; // @[Mux.scala 31:69:@1209.4]
  wire [3:0] _T_2807; // @[Mux.scala 31:69:@1210.4]
  wire [3:0] _T_2808; // @[Mux.scala 31:69:@1211.4]
  wire [3:0] _T_2809; // @[Mux.scala 31:69:@1212.4]
  wire [3:0] _T_2810; // @[Mux.scala 31:69:@1213.4]
  wire [3:0] _T_2811; // @[Mux.scala 31:69:@1214.4]
  wire [3:0] _T_2812; // @[Mux.scala 31:69:@1215.4]
  wire [3:0] _T_2813; // @[Mux.scala 31:69:@1216.4]
  wire [3:0] _T_2814; // @[Mux.scala 31:69:@1217.4]
  wire [3:0] _T_2815; // @[Mux.scala 31:69:@1218.4]
  wire [3:0] _T_2816; // @[Mux.scala 31:69:@1219.4]
  wire [3:0] select_14; // @[Mux.scala 31:69:@1220.4]
  wire [47:0] _GEN_225; // @[Switch.scala 33:19:@1222.4]
  wire [47:0] _GEN_226; // @[Switch.scala 33:19:@1222.4]
  wire [47:0] _GEN_227; // @[Switch.scala 33:19:@1222.4]
  wire [47:0] _GEN_228; // @[Switch.scala 33:19:@1222.4]
  wire [47:0] _GEN_229; // @[Switch.scala 33:19:@1222.4]
  wire [47:0] _GEN_230; // @[Switch.scala 33:19:@1222.4]
  wire [47:0] _GEN_231; // @[Switch.scala 33:19:@1222.4]
  wire [47:0] _GEN_232; // @[Switch.scala 33:19:@1222.4]
  wire [47:0] _GEN_233; // @[Switch.scala 33:19:@1222.4]
  wire [47:0] _GEN_234; // @[Switch.scala 33:19:@1222.4]
  wire [47:0] _GEN_235; // @[Switch.scala 33:19:@1222.4]
  wire [47:0] _GEN_236; // @[Switch.scala 33:19:@1222.4]
  wire [47:0] _GEN_237; // @[Switch.scala 33:19:@1222.4]
  wire [47:0] _GEN_238; // @[Switch.scala 33:19:@1222.4]
  wire [7:0] _T_2825; // @[Switch.scala 34:32:@1229.4]
  wire [15:0] _T_2833; // @[Switch.scala 34:32:@1237.4]
  wire  _T_2837; // @[Switch.scala 30:53:@1240.4]
  wire  valid_15_0; // @[Switch.scala 30:36:@1241.4]
  wire  _T_2840; // @[Switch.scala 30:53:@1243.4]
  wire  valid_15_1; // @[Switch.scala 30:36:@1244.4]
  wire  _T_2843; // @[Switch.scala 30:53:@1246.4]
  wire  valid_15_2; // @[Switch.scala 30:36:@1247.4]
  wire  _T_2846; // @[Switch.scala 30:53:@1249.4]
  wire  valid_15_3; // @[Switch.scala 30:36:@1250.4]
  wire  _T_2849; // @[Switch.scala 30:53:@1252.4]
  wire  valid_15_4; // @[Switch.scala 30:36:@1253.4]
  wire  _T_2852; // @[Switch.scala 30:53:@1255.4]
  wire  valid_15_5; // @[Switch.scala 30:36:@1256.4]
  wire  _T_2855; // @[Switch.scala 30:53:@1258.4]
  wire  valid_15_6; // @[Switch.scala 30:36:@1259.4]
  wire  _T_2858; // @[Switch.scala 30:53:@1261.4]
  wire  valid_15_7; // @[Switch.scala 30:36:@1262.4]
  wire  _T_2861; // @[Switch.scala 30:53:@1264.4]
  wire  valid_15_8; // @[Switch.scala 30:36:@1265.4]
  wire  _T_2864; // @[Switch.scala 30:53:@1267.4]
  wire  valid_15_9; // @[Switch.scala 30:36:@1268.4]
  wire  _T_2867; // @[Switch.scala 30:53:@1270.4]
  wire  valid_15_10; // @[Switch.scala 30:36:@1271.4]
  wire  _T_2870; // @[Switch.scala 30:53:@1273.4]
  wire  valid_15_11; // @[Switch.scala 30:36:@1274.4]
  wire  _T_2873; // @[Switch.scala 30:53:@1276.4]
  wire  valid_15_12; // @[Switch.scala 30:36:@1277.4]
  wire  _T_2876; // @[Switch.scala 30:53:@1279.4]
  wire  valid_15_13; // @[Switch.scala 30:36:@1280.4]
  wire  _T_2879; // @[Switch.scala 30:53:@1282.4]
  wire  valid_15_14; // @[Switch.scala 30:36:@1283.4]
  wire  _T_2882; // @[Switch.scala 30:53:@1285.4]
  wire  valid_15_15; // @[Switch.scala 30:36:@1286.4]
  wire [3:0] _T_2900; // @[Mux.scala 31:69:@1288.4]
  wire [3:0] _T_2901; // @[Mux.scala 31:69:@1289.4]
  wire [3:0] _T_2902; // @[Mux.scala 31:69:@1290.4]
  wire [3:0] _T_2903; // @[Mux.scala 31:69:@1291.4]
  wire [3:0] _T_2904; // @[Mux.scala 31:69:@1292.4]
  wire [3:0] _T_2905; // @[Mux.scala 31:69:@1293.4]
  wire [3:0] _T_2906; // @[Mux.scala 31:69:@1294.4]
  wire [3:0] _T_2907; // @[Mux.scala 31:69:@1295.4]
  wire [3:0] _T_2908; // @[Mux.scala 31:69:@1296.4]
  wire [3:0] _T_2909; // @[Mux.scala 31:69:@1297.4]
  wire [3:0] _T_2910; // @[Mux.scala 31:69:@1298.4]
  wire [3:0] _T_2911; // @[Mux.scala 31:69:@1299.4]
  wire [3:0] _T_2912; // @[Mux.scala 31:69:@1300.4]
  wire [3:0] _T_2913; // @[Mux.scala 31:69:@1301.4]
  wire [3:0] select_15; // @[Mux.scala 31:69:@1302.4]
  wire [47:0] _GEN_241; // @[Switch.scala 33:19:@1304.4]
  wire [47:0] _GEN_242; // @[Switch.scala 33:19:@1304.4]
  wire [47:0] _GEN_243; // @[Switch.scala 33:19:@1304.4]
  wire [47:0] _GEN_244; // @[Switch.scala 33:19:@1304.4]
  wire [47:0] _GEN_245; // @[Switch.scala 33:19:@1304.4]
  wire [47:0] _GEN_246; // @[Switch.scala 33:19:@1304.4]
  wire [47:0] _GEN_247; // @[Switch.scala 33:19:@1304.4]
  wire [47:0] _GEN_248; // @[Switch.scala 33:19:@1304.4]
  wire [47:0] _GEN_249; // @[Switch.scala 33:19:@1304.4]
  wire [47:0] _GEN_250; // @[Switch.scala 33:19:@1304.4]
  wire [47:0] _GEN_251; // @[Switch.scala 33:19:@1304.4]
  wire [47:0] _GEN_252; // @[Switch.scala 33:19:@1304.4]
  wire [47:0] _GEN_253; // @[Switch.scala 33:19:@1304.4]
  wire [47:0] _GEN_254; // @[Switch.scala 33:19:@1304.4]
  wire [7:0] _T_2922; // @[Switch.scala 34:32:@1311.4]
  wire [15:0] _T_2930; // @[Switch.scala 34:32:@1319.4]
  wire  _T_4164; // @[Switch.scala 41:52:@1323.4]
  wire  output_0_0; // @[Switch.scala 41:38:@1324.4]
  wire  _T_4167; // @[Switch.scala 41:52:@1326.4]
  wire  output_0_1; // @[Switch.scala 41:38:@1327.4]
  wire  _T_4170; // @[Switch.scala 41:52:@1329.4]
  wire  output_0_2; // @[Switch.scala 41:38:@1330.4]
  wire  _T_4173; // @[Switch.scala 41:52:@1332.4]
  wire  output_0_3; // @[Switch.scala 41:38:@1333.4]
  wire  _T_4176; // @[Switch.scala 41:52:@1335.4]
  wire  output_0_4; // @[Switch.scala 41:38:@1336.4]
  wire  _T_4179; // @[Switch.scala 41:52:@1338.4]
  wire  output_0_5; // @[Switch.scala 41:38:@1339.4]
  wire  _T_4182; // @[Switch.scala 41:52:@1341.4]
  wire  output_0_6; // @[Switch.scala 41:38:@1342.4]
  wire  _T_4185; // @[Switch.scala 41:52:@1344.4]
  wire  output_0_7; // @[Switch.scala 41:38:@1345.4]
  wire  _T_4188; // @[Switch.scala 41:52:@1347.4]
  wire  output_0_8; // @[Switch.scala 41:38:@1348.4]
  wire  _T_4191; // @[Switch.scala 41:52:@1350.4]
  wire  output_0_9; // @[Switch.scala 41:38:@1351.4]
  wire  _T_4194; // @[Switch.scala 41:52:@1353.4]
  wire  output_0_10; // @[Switch.scala 41:38:@1354.4]
  wire  _T_4197; // @[Switch.scala 41:52:@1356.4]
  wire  output_0_11; // @[Switch.scala 41:38:@1357.4]
  wire  _T_4200; // @[Switch.scala 41:52:@1359.4]
  wire  output_0_12; // @[Switch.scala 41:38:@1360.4]
  wire  _T_4203; // @[Switch.scala 41:52:@1362.4]
  wire  output_0_13; // @[Switch.scala 41:38:@1363.4]
  wire  _T_4206; // @[Switch.scala 41:52:@1365.4]
  wire  output_0_14; // @[Switch.scala 41:38:@1366.4]
  wire  _T_4209; // @[Switch.scala 41:52:@1368.4]
  wire  output_0_15; // @[Switch.scala 41:38:@1369.4]
  wire [7:0] _T_4217; // @[Switch.scala 43:31:@1377.4]
  wire [15:0] _T_4225; // @[Switch.scala 43:31:@1385.4]
  wire  _T_4229; // @[Switch.scala 41:52:@1388.4]
  wire  output_1_0; // @[Switch.scala 41:38:@1389.4]
  wire  _T_4232; // @[Switch.scala 41:52:@1391.4]
  wire  output_1_1; // @[Switch.scala 41:38:@1392.4]
  wire  _T_4235; // @[Switch.scala 41:52:@1394.4]
  wire  output_1_2; // @[Switch.scala 41:38:@1395.4]
  wire  _T_4238; // @[Switch.scala 41:52:@1397.4]
  wire  output_1_3; // @[Switch.scala 41:38:@1398.4]
  wire  _T_4241; // @[Switch.scala 41:52:@1400.4]
  wire  output_1_4; // @[Switch.scala 41:38:@1401.4]
  wire  _T_4244; // @[Switch.scala 41:52:@1403.4]
  wire  output_1_5; // @[Switch.scala 41:38:@1404.4]
  wire  _T_4247; // @[Switch.scala 41:52:@1406.4]
  wire  output_1_6; // @[Switch.scala 41:38:@1407.4]
  wire  _T_4250; // @[Switch.scala 41:52:@1409.4]
  wire  output_1_7; // @[Switch.scala 41:38:@1410.4]
  wire  _T_4253; // @[Switch.scala 41:52:@1412.4]
  wire  output_1_8; // @[Switch.scala 41:38:@1413.4]
  wire  _T_4256; // @[Switch.scala 41:52:@1415.4]
  wire  output_1_9; // @[Switch.scala 41:38:@1416.4]
  wire  _T_4259; // @[Switch.scala 41:52:@1418.4]
  wire  output_1_10; // @[Switch.scala 41:38:@1419.4]
  wire  _T_4262; // @[Switch.scala 41:52:@1421.4]
  wire  output_1_11; // @[Switch.scala 41:38:@1422.4]
  wire  _T_4265; // @[Switch.scala 41:52:@1424.4]
  wire  output_1_12; // @[Switch.scala 41:38:@1425.4]
  wire  _T_4268; // @[Switch.scala 41:52:@1427.4]
  wire  output_1_13; // @[Switch.scala 41:38:@1428.4]
  wire  _T_4271; // @[Switch.scala 41:52:@1430.4]
  wire  output_1_14; // @[Switch.scala 41:38:@1431.4]
  wire  _T_4274; // @[Switch.scala 41:52:@1433.4]
  wire  output_1_15; // @[Switch.scala 41:38:@1434.4]
  wire [7:0] _T_4282; // @[Switch.scala 43:31:@1442.4]
  wire [15:0] _T_4290; // @[Switch.scala 43:31:@1450.4]
  wire  _T_4294; // @[Switch.scala 41:52:@1453.4]
  wire  output_2_0; // @[Switch.scala 41:38:@1454.4]
  wire  _T_4297; // @[Switch.scala 41:52:@1456.4]
  wire  output_2_1; // @[Switch.scala 41:38:@1457.4]
  wire  _T_4300; // @[Switch.scala 41:52:@1459.4]
  wire  output_2_2; // @[Switch.scala 41:38:@1460.4]
  wire  _T_4303; // @[Switch.scala 41:52:@1462.4]
  wire  output_2_3; // @[Switch.scala 41:38:@1463.4]
  wire  _T_4306; // @[Switch.scala 41:52:@1465.4]
  wire  output_2_4; // @[Switch.scala 41:38:@1466.4]
  wire  _T_4309; // @[Switch.scala 41:52:@1468.4]
  wire  output_2_5; // @[Switch.scala 41:38:@1469.4]
  wire  _T_4312; // @[Switch.scala 41:52:@1471.4]
  wire  output_2_6; // @[Switch.scala 41:38:@1472.4]
  wire  _T_4315; // @[Switch.scala 41:52:@1474.4]
  wire  output_2_7; // @[Switch.scala 41:38:@1475.4]
  wire  _T_4318; // @[Switch.scala 41:52:@1477.4]
  wire  output_2_8; // @[Switch.scala 41:38:@1478.4]
  wire  _T_4321; // @[Switch.scala 41:52:@1480.4]
  wire  output_2_9; // @[Switch.scala 41:38:@1481.4]
  wire  _T_4324; // @[Switch.scala 41:52:@1483.4]
  wire  output_2_10; // @[Switch.scala 41:38:@1484.4]
  wire  _T_4327; // @[Switch.scala 41:52:@1486.4]
  wire  output_2_11; // @[Switch.scala 41:38:@1487.4]
  wire  _T_4330; // @[Switch.scala 41:52:@1489.4]
  wire  output_2_12; // @[Switch.scala 41:38:@1490.4]
  wire  _T_4333; // @[Switch.scala 41:52:@1492.4]
  wire  output_2_13; // @[Switch.scala 41:38:@1493.4]
  wire  _T_4336; // @[Switch.scala 41:52:@1495.4]
  wire  output_2_14; // @[Switch.scala 41:38:@1496.4]
  wire  _T_4339; // @[Switch.scala 41:52:@1498.4]
  wire  output_2_15; // @[Switch.scala 41:38:@1499.4]
  wire [7:0] _T_4347; // @[Switch.scala 43:31:@1507.4]
  wire [15:0] _T_4355; // @[Switch.scala 43:31:@1515.4]
  wire  _T_4359; // @[Switch.scala 41:52:@1518.4]
  wire  output_3_0; // @[Switch.scala 41:38:@1519.4]
  wire  _T_4362; // @[Switch.scala 41:52:@1521.4]
  wire  output_3_1; // @[Switch.scala 41:38:@1522.4]
  wire  _T_4365; // @[Switch.scala 41:52:@1524.4]
  wire  output_3_2; // @[Switch.scala 41:38:@1525.4]
  wire  _T_4368; // @[Switch.scala 41:52:@1527.4]
  wire  output_3_3; // @[Switch.scala 41:38:@1528.4]
  wire  _T_4371; // @[Switch.scala 41:52:@1530.4]
  wire  output_3_4; // @[Switch.scala 41:38:@1531.4]
  wire  _T_4374; // @[Switch.scala 41:52:@1533.4]
  wire  output_3_5; // @[Switch.scala 41:38:@1534.4]
  wire  _T_4377; // @[Switch.scala 41:52:@1536.4]
  wire  output_3_6; // @[Switch.scala 41:38:@1537.4]
  wire  _T_4380; // @[Switch.scala 41:52:@1539.4]
  wire  output_3_7; // @[Switch.scala 41:38:@1540.4]
  wire  _T_4383; // @[Switch.scala 41:52:@1542.4]
  wire  output_3_8; // @[Switch.scala 41:38:@1543.4]
  wire  _T_4386; // @[Switch.scala 41:52:@1545.4]
  wire  output_3_9; // @[Switch.scala 41:38:@1546.4]
  wire  _T_4389; // @[Switch.scala 41:52:@1548.4]
  wire  output_3_10; // @[Switch.scala 41:38:@1549.4]
  wire  _T_4392; // @[Switch.scala 41:52:@1551.4]
  wire  output_3_11; // @[Switch.scala 41:38:@1552.4]
  wire  _T_4395; // @[Switch.scala 41:52:@1554.4]
  wire  output_3_12; // @[Switch.scala 41:38:@1555.4]
  wire  _T_4398; // @[Switch.scala 41:52:@1557.4]
  wire  output_3_13; // @[Switch.scala 41:38:@1558.4]
  wire  _T_4401; // @[Switch.scala 41:52:@1560.4]
  wire  output_3_14; // @[Switch.scala 41:38:@1561.4]
  wire  _T_4404; // @[Switch.scala 41:52:@1563.4]
  wire  output_3_15; // @[Switch.scala 41:38:@1564.4]
  wire [7:0] _T_4412; // @[Switch.scala 43:31:@1572.4]
  wire [15:0] _T_4420; // @[Switch.scala 43:31:@1580.4]
  wire  _T_4424; // @[Switch.scala 41:52:@1583.4]
  wire  output_4_0; // @[Switch.scala 41:38:@1584.4]
  wire  _T_4427; // @[Switch.scala 41:52:@1586.4]
  wire  output_4_1; // @[Switch.scala 41:38:@1587.4]
  wire  _T_4430; // @[Switch.scala 41:52:@1589.4]
  wire  output_4_2; // @[Switch.scala 41:38:@1590.4]
  wire  _T_4433; // @[Switch.scala 41:52:@1592.4]
  wire  output_4_3; // @[Switch.scala 41:38:@1593.4]
  wire  _T_4436; // @[Switch.scala 41:52:@1595.4]
  wire  output_4_4; // @[Switch.scala 41:38:@1596.4]
  wire  _T_4439; // @[Switch.scala 41:52:@1598.4]
  wire  output_4_5; // @[Switch.scala 41:38:@1599.4]
  wire  _T_4442; // @[Switch.scala 41:52:@1601.4]
  wire  output_4_6; // @[Switch.scala 41:38:@1602.4]
  wire  _T_4445; // @[Switch.scala 41:52:@1604.4]
  wire  output_4_7; // @[Switch.scala 41:38:@1605.4]
  wire  _T_4448; // @[Switch.scala 41:52:@1607.4]
  wire  output_4_8; // @[Switch.scala 41:38:@1608.4]
  wire  _T_4451; // @[Switch.scala 41:52:@1610.4]
  wire  output_4_9; // @[Switch.scala 41:38:@1611.4]
  wire  _T_4454; // @[Switch.scala 41:52:@1613.4]
  wire  output_4_10; // @[Switch.scala 41:38:@1614.4]
  wire  _T_4457; // @[Switch.scala 41:52:@1616.4]
  wire  output_4_11; // @[Switch.scala 41:38:@1617.4]
  wire  _T_4460; // @[Switch.scala 41:52:@1619.4]
  wire  output_4_12; // @[Switch.scala 41:38:@1620.4]
  wire  _T_4463; // @[Switch.scala 41:52:@1622.4]
  wire  output_4_13; // @[Switch.scala 41:38:@1623.4]
  wire  _T_4466; // @[Switch.scala 41:52:@1625.4]
  wire  output_4_14; // @[Switch.scala 41:38:@1626.4]
  wire  _T_4469; // @[Switch.scala 41:52:@1628.4]
  wire  output_4_15; // @[Switch.scala 41:38:@1629.4]
  wire [7:0] _T_4477; // @[Switch.scala 43:31:@1637.4]
  wire [15:0] _T_4485; // @[Switch.scala 43:31:@1645.4]
  wire  _T_4489; // @[Switch.scala 41:52:@1648.4]
  wire  output_5_0; // @[Switch.scala 41:38:@1649.4]
  wire  _T_4492; // @[Switch.scala 41:52:@1651.4]
  wire  output_5_1; // @[Switch.scala 41:38:@1652.4]
  wire  _T_4495; // @[Switch.scala 41:52:@1654.4]
  wire  output_5_2; // @[Switch.scala 41:38:@1655.4]
  wire  _T_4498; // @[Switch.scala 41:52:@1657.4]
  wire  output_5_3; // @[Switch.scala 41:38:@1658.4]
  wire  _T_4501; // @[Switch.scala 41:52:@1660.4]
  wire  output_5_4; // @[Switch.scala 41:38:@1661.4]
  wire  _T_4504; // @[Switch.scala 41:52:@1663.4]
  wire  output_5_5; // @[Switch.scala 41:38:@1664.4]
  wire  _T_4507; // @[Switch.scala 41:52:@1666.4]
  wire  output_5_6; // @[Switch.scala 41:38:@1667.4]
  wire  _T_4510; // @[Switch.scala 41:52:@1669.4]
  wire  output_5_7; // @[Switch.scala 41:38:@1670.4]
  wire  _T_4513; // @[Switch.scala 41:52:@1672.4]
  wire  output_5_8; // @[Switch.scala 41:38:@1673.4]
  wire  _T_4516; // @[Switch.scala 41:52:@1675.4]
  wire  output_5_9; // @[Switch.scala 41:38:@1676.4]
  wire  _T_4519; // @[Switch.scala 41:52:@1678.4]
  wire  output_5_10; // @[Switch.scala 41:38:@1679.4]
  wire  _T_4522; // @[Switch.scala 41:52:@1681.4]
  wire  output_5_11; // @[Switch.scala 41:38:@1682.4]
  wire  _T_4525; // @[Switch.scala 41:52:@1684.4]
  wire  output_5_12; // @[Switch.scala 41:38:@1685.4]
  wire  _T_4528; // @[Switch.scala 41:52:@1687.4]
  wire  output_5_13; // @[Switch.scala 41:38:@1688.4]
  wire  _T_4531; // @[Switch.scala 41:52:@1690.4]
  wire  output_5_14; // @[Switch.scala 41:38:@1691.4]
  wire  _T_4534; // @[Switch.scala 41:52:@1693.4]
  wire  output_5_15; // @[Switch.scala 41:38:@1694.4]
  wire [7:0] _T_4542; // @[Switch.scala 43:31:@1702.4]
  wire [15:0] _T_4550; // @[Switch.scala 43:31:@1710.4]
  wire  _T_4554; // @[Switch.scala 41:52:@1713.4]
  wire  output_6_0; // @[Switch.scala 41:38:@1714.4]
  wire  _T_4557; // @[Switch.scala 41:52:@1716.4]
  wire  output_6_1; // @[Switch.scala 41:38:@1717.4]
  wire  _T_4560; // @[Switch.scala 41:52:@1719.4]
  wire  output_6_2; // @[Switch.scala 41:38:@1720.4]
  wire  _T_4563; // @[Switch.scala 41:52:@1722.4]
  wire  output_6_3; // @[Switch.scala 41:38:@1723.4]
  wire  _T_4566; // @[Switch.scala 41:52:@1725.4]
  wire  output_6_4; // @[Switch.scala 41:38:@1726.4]
  wire  _T_4569; // @[Switch.scala 41:52:@1728.4]
  wire  output_6_5; // @[Switch.scala 41:38:@1729.4]
  wire  _T_4572; // @[Switch.scala 41:52:@1731.4]
  wire  output_6_6; // @[Switch.scala 41:38:@1732.4]
  wire  _T_4575; // @[Switch.scala 41:52:@1734.4]
  wire  output_6_7; // @[Switch.scala 41:38:@1735.4]
  wire  _T_4578; // @[Switch.scala 41:52:@1737.4]
  wire  output_6_8; // @[Switch.scala 41:38:@1738.4]
  wire  _T_4581; // @[Switch.scala 41:52:@1740.4]
  wire  output_6_9; // @[Switch.scala 41:38:@1741.4]
  wire  _T_4584; // @[Switch.scala 41:52:@1743.4]
  wire  output_6_10; // @[Switch.scala 41:38:@1744.4]
  wire  _T_4587; // @[Switch.scala 41:52:@1746.4]
  wire  output_6_11; // @[Switch.scala 41:38:@1747.4]
  wire  _T_4590; // @[Switch.scala 41:52:@1749.4]
  wire  output_6_12; // @[Switch.scala 41:38:@1750.4]
  wire  _T_4593; // @[Switch.scala 41:52:@1752.4]
  wire  output_6_13; // @[Switch.scala 41:38:@1753.4]
  wire  _T_4596; // @[Switch.scala 41:52:@1755.4]
  wire  output_6_14; // @[Switch.scala 41:38:@1756.4]
  wire  _T_4599; // @[Switch.scala 41:52:@1758.4]
  wire  output_6_15; // @[Switch.scala 41:38:@1759.4]
  wire [7:0] _T_4607; // @[Switch.scala 43:31:@1767.4]
  wire [15:0] _T_4615; // @[Switch.scala 43:31:@1775.4]
  wire  _T_4619; // @[Switch.scala 41:52:@1778.4]
  wire  output_7_0; // @[Switch.scala 41:38:@1779.4]
  wire  _T_4622; // @[Switch.scala 41:52:@1781.4]
  wire  output_7_1; // @[Switch.scala 41:38:@1782.4]
  wire  _T_4625; // @[Switch.scala 41:52:@1784.4]
  wire  output_7_2; // @[Switch.scala 41:38:@1785.4]
  wire  _T_4628; // @[Switch.scala 41:52:@1787.4]
  wire  output_7_3; // @[Switch.scala 41:38:@1788.4]
  wire  _T_4631; // @[Switch.scala 41:52:@1790.4]
  wire  output_7_4; // @[Switch.scala 41:38:@1791.4]
  wire  _T_4634; // @[Switch.scala 41:52:@1793.4]
  wire  output_7_5; // @[Switch.scala 41:38:@1794.4]
  wire  _T_4637; // @[Switch.scala 41:52:@1796.4]
  wire  output_7_6; // @[Switch.scala 41:38:@1797.4]
  wire  _T_4640; // @[Switch.scala 41:52:@1799.4]
  wire  output_7_7; // @[Switch.scala 41:38:@1800.4]
  wire  _T_4643; // @[Switch.scala 41:52:@1802.4]
  wire  output_7_8; // @[Switch.scala 41:38:@1803.4]
  wire  _T_4646; // @[Switch.scala 41:52:@1805.4]
  wire  output_7_9; // @[Switch.scala 41:38:@1806.4]
  wire  _T_4649; // @[Switch.scala 41:52:@1808.4]
  wire  output_7_10; // @[Switch.scala 41:38:@1809.4]
  wire  _T_4652; // @[Switch.scala 41:52:@1811.4]
  wire  output_7_11; // @[Switch.scala 41:38:@1812.4]
  wire  _T_4655; // @[Switch.scala 41:52:@1814.4]
  wire  output_7_12; // @[Switch.scala 41:38:@1815.4]
  wire  _T_4658; // @[Switch.scala 41:52:@1817.4]
  wire  output_7_13; // @[Switch.scala 41:38:@1818.4]
  wire  _T_4661; // @[Switch.scala 41:52:@1820.4]
  wire  output_7_14; // @[Switch.scala 41:38:@1821.4]
  wire  _T_4664; // @[Switch.scala 41:52:@1823.4]
  wire  output_7_15; // @[Switch.scala 41:38:@1824.4]
  wire [7:0] _T_4672; // @[Switch.scala 43:31:@1832.4]
  wire [15:0] _T_4680; // @[Switch.scala 43:31:@1840.4]
  wire  _T_4684; // @[Switch.scala 41:52:@1843.4]
  wire  output_8_0; // @[Switch.scala 41:38:@1844.4]
  wire  _T_4687; // @[Switch.scala 41:52:@1846.4]
  wire  output_8_1; // @[Switch.scala 41:38:@1847.4]
  wire  _T_4690; // @[Switch.scala 41:52:@1849.4]
  wire  output_8_2; // @[Switch.scala 41:38:@1850.4]
  wire  _T_4693; // @[Switch.scala 41:52:@1852.4]
  wire  output_8_3; // @[Switch.scala 41:38:@1853.4]
  wire  _T_4696; // @[Switch.scala 41:52:@1855.4]
  wire  output_8_4; // @[Switch.scala 41:38:@1856.4]
  wire  _T_4699; // @[Switch.scala 41:52:@1858.4]
  wire  output_8_5; // @[Switch.scala 41:38:@1859.4]
  wire  _T_4702; // @[Switch.scala 41:52:@1861.4]
  wire  output_8_6; // @[Switch.scala 41:38:@1862.4]
  wire  _T_4705; // @[Switch.scala 41:52:@1864.4]
  wire  output_8_7; // @[Switch.scala 41:38:@1865.4]
  wire  _T_4708; // @[Switch.scala 41:52:@1867.4]
  wire  output_8_8; // @[Switch.scala 41:38:@1868.4]
  wire  _T_4711; // @[Switch.scala 41:52:@1870.4]
  wire  output_8_9; // @[Switch.scala 41:38:@1871.4]
  wire  _T_4714; // @[Switch.scala 41:52:@1873.4]
  wire  output_8_10; // @[Switch.scala 41:38:@1874.4]
  wire  _T_4717; // @[Switch.scala 41:52:@1876.4]
  wire  output_8_11; // @[Switch.scala 41:38:@1877.4]
  wire  _T_4720; // @[Switch.scala 41:52:@1879.4]
  wire  output_8_12; // @[Switch.scala 41:38:@1880.4]
  wire  _T_4723; // @[Switch.scala 41:52:@1882.4]
  wire  output_8_13; // @[Switch.scala 41:38:@1883.4]
  wire  _T_4726; // @[Switch.scala 41:52:@1885.4]
  wire  output_8_14; // @[Switch.scala 41:38:@1886.4]
  wire  _T_4729; // @[Switch.scala 41:52:@1888.4]
  wire  output_8_15; // @[Switch.scala 41:38:@1889.4]
  wire [7:0] _T_4737; // @[Switch.scala 43:31:@1897.4]
  wire [15:0] _T_4745; // @[Switch.scala 43:31:@1905.4]
  wire  _T_4749; // @[Switch.scala 41:52:@1908.4]
  wire  output_9_0; // @[Switch.scala 41:38:@1909.4]
  wire  _T_4752; // @[Switch.scala 41:52:@1911.4]
  wire  output_9_1; // @[Switch.scala 41:38:@1912.4]
  wire  _T_4755; // @[Switch.scala 41:52:@1914.4]
  wire  output_9_2; // @[Switch.scala 41:38:@1915.4]
  wire  _T_4758; // @[Switch.scala 41:52:@1917.4]
  wire  output_9_3; // @[Switch.scala 41:38:@1918.4]
  wire  _T_4761; // @[Switch.scala 41:52:@1920.4]
  wire  output_9_4; // @[Switch.scala 41:38:@1921.4]
  wire  _T_4764; // @[Switch.scala 41:52:@1923.4]
  wire  output_9_5; // @[Switch.scala 41:38:@1924.4]
  wire  _T_4767; // @[Switch.scala 41:52:@1926.4]
  wire  output_9_6; // @[Switch.scala 41:38:@1927.4]
  wire  _T_4770; // @[Switch.scala 41:52:@1929.4]
  wire  output_9_7; // @[Switch.scala 41:38:@1930.4]
  wire  _T_4773; // @[Switch.scala 41:52:@1932.4]
  wire  output_9_8; // @[Switch.scala 41:38:@1933.4]
  wire  _T_4776; // @[Switch.scala 41:52:@1935.4]
  wire  output_9_9; // @[Switch.scala 41:38:@1936.4]
  wire  _T_4779; // @[Switch.scala 41:52:@1938.4]
  wire  output_9_10; // @[Switch.scala 41:38:@1939.4]
  wire  _T_4782; // @[Switch.scala 41:52:@1941.4]
  wire  output_9_11; // @[Switch.scala 41:38:@1942.4]
  wire  _T_4785; // @[Switch.scala 41:52:@1944.4]
  wire  output_9_12; // @[Switch.scala 41:38:@1945.4]
  wire  _T_4788; // @[Switch.scala 41:52:@1947.4]
  wire  output_9_13; // @[Switch.scala 41:38:@1948.4]
  wire  _T_4791; // @[Switch.scala 41:52:@1950.4]
  wire  output_9_14; // @[Switch.scala 41:38:@1951.4]
  wire  _T_4794; // @[Switch.scala 41:52:@1953.4]
  wire  output_9_15; // @[Switch.scala 41:38:@1954.4]
  wire [7:0] _T_4802; // @[Switch.scala 43:31:@1962.4]
  wire [15:0] _T_4810; // @[Switch.scala 43:31:@1970.4]
  wire  _T_4814; // @[Switch.scala 41:52:@1973.4]
  wire  output_10_0; // @[Switch.scala 41:38:@1974.4]
  wire  _T_4817; // @[Switch.scala 41:52:@1976.4]
  wire  output_10_1; // @[Switch.scala 41:38:@1977.4]
  wire  _T_4820; // @[Switch.scala 41:52:@1979.4]
  wire  output_10_2; // @[Switch.scala 41:38:@1980.4]
  wire  _T_4823; // @[Switch.scala 41:52:@1982.4]
  wire  output_10_3; // @[Switch.scala 41:38:@1983.4]
  wire  _T_4826; // @[Switch.scala 41:52:@1985.4]
  wire  output_10_4; // @[Switch.scala 41:38:@1986.4]
  wire  _T_4829; // @[Switch.scala 41:52:@1988.4]
  wire  output_10_5; // @[Switch.scala 41:38:@1989.4]
  wire  _T_4832; // @[Switch.scala 41:52:@1991.4]
  wire  output_10_6; // @[Switch.scala 41:38:@1992.4]
  wire  _T_4835; // @[Switch.scala 41:52:@1994.4]
  wire  output_10_7; // @[Switch.scala 41:38:@1995.4]
  wire  _T_4838; // @[Switch.scala 41:52:@1997.4]
  wire  output_10_8; // @[Switch.scala 41:38:@1998.4]
  wire  _T_4841; // @[Switch.scala 41:52:@2000.4]
  wire  output_10_9; // @[Switch.scala 41:38:@2001.4]
  wire  _T_4844; // @[Switch.scala 41:52:@2003.4]
  wire  output_10_10; // @[Switch.scala 41:38:@2004.4]
  wire  _T_4847; // @[Switch.scala 41:52:@2006.4]
  wire  output_10_11; // @[Switch.scala 41:38:@2007.4]
  wire  _T_4850; // @[Switch.scala 41:52:@2009.4]
  wire  output_10_12; // @[Switch.scala 41:38:@2010.4]
  wire  _T_4853; // @[Switch.scala 41:52:@2012.4]
  wire  output_10_13; // @[Switch.scala 41:38:@2013.4]
  wire  _T_4856; // @[Switch.scala 41:52:@2015.4]
  wire  output_10_14; // @[Switch.scala 41:38:@2016.4]
  wire  _T_4859; // @[Switch.scala 41:52:@2018.4]
  wire  output_10_15; // @[Switch.scala 41:38:@2019.4]
  wire [7:0] _T_4867; // @[Switch.scala 43:31:@2027.4]
  wire [15:0] _T_4875; // @[Switch.scala 43:31:@2035.4]
  wire  _T_4879; // @[Switch.scala 41:52:@2038.4]
  wire  output_11_0; // @[Switch.scala 41:38:@2039.4]
  wire  _T_4882; // @[Switch.scala 41:52:@2041.4]
  wire  output_11_1; // @[Switch.scala 41:38:@2042.4]
  wire  _T_4885; // @[Switch.scala 41:52:@2044.4]
  wire  output_11_2; // @[Switch.scala 41:38:@2045.4]
  wire  _T_4888; // @[Switch.scala 41:52:@2047.4]
  wire  output_11_3; // @[Switch.scala 41:38:@2048.4]
  wire  _T_4891; // @[Switch.scala 41:52:@2050.4]
  wire  output_11_4; // @[Switch.scala 41:38:@2051.4]
  wire  _T_4894; // @[Switch.scala 41:52:@2053.4]
  wire  output_11_5; // @[Switch.scala 41:38:@2054.4]
  wire  _T_4897; // @[Switch.scala 41:52:@2056.4]
  wire  output_11_6; // @[Switch.scala 41:38:@2057.4]
  wire  _T_4900; // @[Switch.scala 41:52:@2059.4]
  wire  output_11_7; // @[Switch.scala 41:38:@2060.4]
  wire  _T_4903; // @[Switch.scala 41:52:@2062.4]
  wire  output_11_8; // @[Switch.scala 41:38:@2063.4]
  wire  _T_4906; // @[Switch.scala 41:52:@2065.4]
  wire  output_11_9; // @[Switch.scala 41:38:@2066.4]
  wire  _T_4909; // @[Switch.scala 41:52:@2068.4]
  wire  output_11_10; // @[Switch.scala 41:38:@2069.4]
  wire  _T_4912; // @[Switch.scala 41:52:@2071.4]
  wire  output_11_11; // @[Switch.scala 41:38:@2072.4]
  wire  _T_4915; // @[Switch.scala 41:52:@2074.4]
  wire  output_11_12; // @[Switch.scala 41:38:@2075.4]
  wire  _T_4918; // @[Switch.scala 41:52:@2077.4]
  wire  output_11_13; // @[Switch.scala 41:38:@2078.4]
  wire  _T_4921; // @[Switch.scala 41:52:@2080.4]
  wire  output_11_14; // @[Switch.scala 41:38:@2081.4]
  wire  _T_4924; // @[Switch.scala 41:52:@2083.4]
  wire  output_11_15; // @[Switch.scala 41:38:@2084.4]
  wire [7:0] _T_4932; // @[Switch.scala 43:31:@2092.4]
  wire [15:0] _T_4940; // @[Switch.scala 43:31:@2100.4]
  wire  _T_4944; // @[Switch.scala 41:52:@2103.4]
  wire  output_12_0; // @[Switch.scala 41:38:@2104.4]
  wire  _T_4947; // @[Switch.scala 41:52:@2106.4]
  wire  output_12_1; // @[Switch.scala 41:38:@2107.4]
  wire  _T_4950; // @[Switch.scala 41:52:@2109.4]
  wire  output_12_2; // @[Switch.scala 41:38:@2110.4]
  wire  _T_4953; // @[Switch.scala 41:52:@2112.4]
  wire  output_12_3; // @[Switch.scala 41:38:@2113.4]
  wire  _T_4956; // @[Switch.scala 41:52:@2115.4]
  wire  output_12_4; // @[Switch.scala 41:38:@2116.4]
  wire  _T_4959; // @[Switch.scala 41:52:@2118.4]
  wire  output_12_5; // @[Switch.scala 41:38:@2119.4]
  wire  _T_4962; // @[Switch.scala 41:52:@2121.4]
  wire  output_12_6; // @[Switch.scala 41:38:@2122.4]
  wire  _T_4965; // @[Switch.scala 41:52:@2124.4]
  wire  output_12_7; // @[Switch.scala 41:38:@2125.4]
  wire  _T_4968; // @[Switch.scala 41:52:@2127.4]
  wire  output_12_8; // @[Switch.scala 41:38:@2128.4]
  wire  _T_4971; // @[Switch.scala 41:52:@2130.4]
  wire  output_12_9; // @[Switch.scala 41:38:@2131.4]
  wire  _T_4974; // @[Switch.scala 41:52:@2133.4]
  wire  output_12_10; // @[Switch.scala 41:38:@2134.4]
  wire  _T_4977; // @[Switch.scala 41:52:@2136.4]
  wire  output_12_11; // @[Switch.scala 41:38:@2137.4]
  wire  _T_4980; // @[Switch.scala 41:52:@2139.4]
  wire  output_12_12; // @[Switch.scala 41:38:@2140.4]
  wire  _T_4983; // @[Switch.scala 41:52:@2142.4]
  wire  output_12_13; // @[Switch.scala 41:38:@2143.4]
  wire  _T_4986; // @[Switch.scala 41:52:@2145.4]
  wire  output_12_14; // @[Switch.scala 41:38:@2146.4]
  wire  _T_4989; // @[Switch.scala 41:52:@2148.4]
  wire  output_12_15; // @[Switch.scala 41:38:@2149.4]
  wire [7:0] _T_4997; // @[Switch.scala 43:31:@2157.4]
  wire [15:0] _T_5005; // @[Switch.scala 43:31:@2165.4]
  wire  _T_5009; // @[Switch.scala 41:52:@2168.4]
  wire  output_13_0; // @[Switch.scala 41:38:@2169.4]
  wire  _T_5012; // @[Switch.scala 41:52:@2171.4]
  wire  output_13_1; // @[Switch.scala 41:38:@2172.4]
  wire  _T_5015; // @[Switch.scala 41:52:@2174.4]
  wire  output_13_2; // @[Switch.scala 41:38:@2175.4]
  wire  _T_5018; // @[Switch.scala 41:52:@2177.4]
  wire  output_13_3; // @[Switch.scala 41:38:@2178.4]
  wire  _T_5021; // @[Switch.scala 41:52:@2180.4]
  wire  output_13_4; // @[Switch.scala 41:38:@2181.4]
  wire  _T_5024; // @[Switch.scala 41:52:@2183.4]
  wire  output_13_5; // @[Switch.scala 41:38:@2184.4]
  wire  _T_5027; // @[Switch.scala 41:52:@2186.4]
  wire  output_13_6; // @[Switch.scala 41:38:@2187.4]
  wire  _T_5030; // @[Switch.scala 41:52:@2189.4]
  wire  output_13_7; // @[Switch.scala 41:38:@2190.4]
  wire  _T_5033; // @[Switch.scala 41:52:@2192.4]
  wire  output_13_8; // @[Switch.scala 41:38:@2193.4]
  wire  _T_5036; // @[Switch.scala 41:52:@2195.4]
  wire  output_13_9; // @[Switch.scala 41:38:@2196.4]
  wire  _T_5039; // @[Switch.scala 41:52:@2198.4]
  wire  output_13_10; // @[Switch.scala 41:38:@2199.4]
  wire  _T_5042; // @[Switch.scala 41:52:@2201.4]
  wire  output_13_11; // @[Switch.scala 41:38:@2202.4]
  wire  _T_5045; // @[Switch.scala 41:52:@2204.4]
  wire  output_13_12; // @[Switch.scala 41:38:@2205.4]
  wire  _T_5048; // @[Switch.scala 41:52:@2207.4]
  wire  output_13_13; // @[Switch.scala 41:38:@2208.4]
  wire  _T_5051; // @[Switch.scala 41:52:@2210.4]
  wire  output_13_14; // @[Switch.scala 41:38:@2211.4]
  wire  _T_5054; // @[Switch.scala 41:52:@2213.4]
  wire  output_13_15; // @[Switch.scala 41:38:@2214.4]
  wire [7:0] _T_5062; // @[Switch.scala 43:31:@2222.4]
  wire [15:0] _T_5070; // @[Switch.scala 43:31:@2230.4]
  wire  _T_5074; // @[Switch.scala 41:52:@2233.4]
  wire  output_14_0; // @[Switch.scala 41:38:@2234.4]
  wire  _T_5077; // @[Switch.scala 41:52:@2236.4]
  wire  output_14_1; // @[Switch.scala 41:38:@2237.4]
  wire  _T_5080; // @[Switch.scala 41:52:@2239.4]
  wire  output_14_2; // @[Switch.scala 41:38:@2240.4]
  wire  _T_5083; // @[Switch.scala 41:52:@2242.4]
  wire  output_14_3; // @[Switch.scala 41:38:@2243.4]
  wire  _T_5086; // @[Switch.scala 41:52:@2245.4]
  wire  output_14_4; // @[Switch.scala 41:38:@2246.4]
  wire  _T_5089; // @[Switch.scala 41:52:@2248.4]
  wire  output_14_5; // @[Switch.scala 41:38:@2249.4]
  wire  _T_5092; // @[Switch.scala 41:52:@2251.4]
  wire  output_14_6; // @[Switch.scala 41:38:@2252.4]
  wire  _T_5095; // @[Switch.scala 41:52:@2254.4]
  wire  output_14_7; // @[Switch.scala 41:38:@2255.4]
  wire  _T_5098; // @[Switch.scala 41:52:@2257.4]
  wire  output_14_8; // @[Switch.scala 41:38:@2258.4]
  wire  _T_5101; // @[Switch.scala 41:52:@2260.4]
  wire  output_14_9; // @[Switch.scala 41:38:@2261.4]
  wire  _T_5104; // @[Switch.scala 41:52:@2263.4]
  wire  output_14_10; // @[Switch.scala 41:38:@2264.4]
  wire  _T_5107; // @[Switch.scala 41:52:@2266.4]
  wire  output_14_11; // @[Switch.scala 41:38:@2267.4]
  wire  _T_5110; // @[Switch.scala 41:52:@2269.4]
  wire  output_14_12; // @[Switch.scala 41:38:@2270.4]
  wire  _T_5113; // @[Switch.scala 41:52:@2272.4]
  wire  output_14_13; // @[Switch.scala 41:38:@2273.4]
  wire  _T_5116; // @[Switch.scala 41:52:@2275.4]
  wire  output_14_14; // @[Switch.scala 41:38:@2276.4]
  wire  _T_5119; // @[Switch.scala 41:52:@2278.4]
  wire  output_14_15; // @[Switch.scala 41:38:@2279.4]
  wire [7:0] _T_5127; // @[Switch.scala 43:31:@2287.4]
  wire [15:0] _T_5135; // @[Switch.scala 43:31:@2295.4]
  wire  _T_5139; // @[Switch.scala 41:52:@2298.4]
  wire  output_15_0; // @[Switch.scala 41:38:@2299.4]
  wire  _T_5142; // @[Switch.scala 41:52:@2301.4]
  wire  output_15_1; // @[Switch.scala 41:38:@2302.4]
  wire  _T_5145; // @[Switch.scala 41:52:@2304.4]
  wire  output_15_2; // @[Switch.scala 41:38:@2305.4]
  wire  _T_5148; // @[Switch.scala 41:52:@2307.4]
  wire  output_15_3; // @[Switch.scala 41:38:@2308.4]
  wire  _T_5151; // @[Switch.scala 41:52:@2310.4]
  wire  output_15_4; // @[Switch.scala 41:38:@2311.4]
  wire  _T_5154; // @[Switch.scala 41:52:@2313.4]
  wire  output_15_5; // @[Switch.scala 41:38:@2314.4]
  wire  _T_5157; // @[Switch.scala 41:52:@2316.4]
  wire  output_15_6; // @[Switch.scala 41:38:@2317.4]
  wire  _T_5160; // @[Switch.scala 41:52:@2319.4]
  wire  output_15_7; // @[Switch.scala 41:38:@2320.4]
  wire  _T_5163; // @[Switch.scala 41:52:@2322.4]
  wire  output_15_8; // @[Switch.scala 41:38:@2323.4]
  wire  _T_5166; // @[Switch.scala 41:52:@2325.4]
  wire  output_15_9; // @[Switch.scala 41:38:@2326.4]
  wire  _T_5169; // @[Switch.scala 41:52:@2328.4]
  wire  output_15_10; // @[Switch.scala 41:38:@2329.4]
  wire  _T_5172; // @[Switch.scala 41:52:@2331.4]
  wire  output_15_11; // @[Switch.scala 41:38:@2332.4]
  wire  _T_5175; // @[Switch.scala 41:52:@2334.4]
  wire  output_15_12; // @[Switch.scala 41:38:@2335.4]
  wire  _T_5178; // @[Switch.scala 41:52:@2337.4]
  wire  output_15_13; // @[Switch.scala 41:38:@2338.4]
  wire  _T_5181; // @[Switch.scala 41:52:@2340.4]
  wire  output_15_14; // @[Switch.scala 41:38:@2341.4]
  wire  _T_5184; // @[Switch.scala 41:52:@2343.4]
  wire  output_15_15; // @[Switch.scala 41:38:@2344.4]
  wire [7:0] _T_5192; // @[Switch.scala 43:31:@2352.4]
  wire [15:0] _T_5200; // @[Switch.scala 43:31:@2360.4]
  assign _T_1382 = io_inAddr_0 == 4'h0; // @[Switch.scala 30:53:@10.4]
  assign valid_0_0 = io_inValid_0 & _T_1382; // @[Switch.scala 30:36:@11.4]
  assign _T_1385 = io_inAddr_1 == 4'h0; // @[Switch.scala 30:53:@13.4]
  assign valid_0_1 = io_inValid_1 & _T_1385; // @[Switch.scala 30:36:@14.4]
  assign _T_1388 = io_inAddr_2 == 4'h0; // @[Switch.scala 30:53:@16.4]
  assign valid_0_2 = io_inValid_2 & _T_1388; // @[Switch.scala 30:36:@17.4]
  assign _T_1391 = io_inAddr_3 == 4'h0; // @[Switch.scala 30:53:@19.4]
  assign valid_0_3 = io_inValid_3 & _T_1391; // @[Switch.scala 30:36:@20.4]
  assign _T_1394 = io_inAddr_4 == 4'h0; // @[Switch.scala 30:53:@22.4]
  assign valid_0_4 = io_inValid_4 & _T_1394; // @[Switch.scala 30:36:@23.4]
  assign _T_1397 = io_inAddr_5 == 4'h0; // @[Switch.scala 30:53:@25.4]
  assign valid_0_5 = io_inValid_5 & _T_1397; // @[Switch.scala 30:36:@26.4]
  assign _T_1400 = io_inAddr_6 == 4'h0; // @[Switch.scala 30:53:@28.4]
  assign valid_0_6 = io_inValid_6 & _T_1400; // @[Switch.scala 30:36:@29.4]
  assign _T_1403 = io_inAddr_7 == 4'h0; // @[Switch.scala 30:53:@31.4]
  assign valid_0_7 = io_inValid_7 & _T_1403; // @[Switch.scala 30:36:@32.4]
  assign _T_1406 = io_inAddr_8 == 4'h0; // @[Switch.scala 30:53:@34.4]
  assign valid_0_8 = io_inValid_8 & _T_1406; // @[Switch.scala 30:36:@35.4]
  assign _T_1409 = io_inAddr_9 == 4'h0; // @[Switch.scala 30:53:@37.4]
  assign valid_0_9 = io_inValid_9 & _T_1409; // @[Switch.scala 30:36:@38.4]
  assign _T_1412 = io_inAddr_10 == 4'h0; // @[Switch.scala 30:53:@40.4]
  assign valid_0_10 = io_inValid_10 & _T_1412; // @[Switch.scala 30:36:@41.4]
  assign _T_1415 = io_inAddr_11 == 4'h0; // @[Switch.scala 30:53:@43.4]
  assign valid_0_11 = io_inValid_11 & _T_1415; // @[Switch.scala 30:36:@44.4]
  assign _T_1418 = io_inAddr_12 == 4'h0; // @[Switch.scala 30:53:@46.4]
  assign valid_0_12 = io_inValid_12 & _T_1418; // @[Switch.scala 30:36:@47.4]
  assign _T_1421 = io_inAddr_13 == 4'h0; // @[Switch.scala 30:53:@49.4]
  assign valid_0_13 = io_inValid_13 & _T_1421; // @[Switch.scala 30:36:@50.4]
  assign _T_1424 = io_inAddr_14 == 4'h0; // @[Switch.scala 30:53:@52.4]
  assign valid_0_14 = io_inValid_14 & _T_1424; // @[Switch.scala 30:36:@53.4]
  assign _T_1427 = io_inAddr_15 == 4'h0; // @[Switch.scala 30:53:@55.4]
  assign valid_0_15 = io_inValid_15 & _T_1427; // @[Switch.scala 30:36:@56.4]
  assign _T_1445 = valid_0_14 ? 4'he : 4'hf; // @[Mux.scala 31:69:@58.4]
  assign _T_1446 = valid_0_13 ? 4'hd : _T_1445; // @[Mux.scala 31:69:@59.4]
  assign _T_1447 = valid_0_12 ? 4'hc : _T_1446; // @[Mux.scala 31:69:@60.4]
  assign _T_1448 = valid_0_11 ? 4'hb : _T_1447; // @[Mux.scala 31:69:@61.4]
  assign _T_1449 = valid_0_10 ? 4'ha : _T_1448; // @[Mux.scala 31:69:@62.4]
  assign _T_1450 = valid_0_9 ? 4'h9 : _T_1449; // @[Mux.scala 31:69:@63.4]
  assign _T_1451 = valid_0_8 ? 4'h8 : _T_1450; // @[Mux.scala 31:69:@64.4]
  assign _T_1452 = valid_0_7 ? 4'h7 : _T_1451; // @[Mux.scala 31:69:@65.4]
  assign _T_1453 = valid_0_6 ? 4'h6 : _T_1452; // @[Mux.scala 31:69:@66.4]
  assign _T_1454 = valid_0_5 ? 4'h5 : _T_1453; // @[Mux.scala 31:69:@67.4]
  assign _T_1455 = valid_0_4 ? 4'h4 : _T_1454; // @[Mux.scala 31:69:@68.4]
  assign _T_1456 = valid_0_3 ? 4'h3 : _T_1455; // @[Mux.scala 31:69:@69.4]
  assign _T_1457 = valid_0_2 ? 4'h2 : _T_1456; // @[Mux.scala 31:69:@70.4]
  assign _T_1458 = valid_0_1 ? 4'h1 : _T_1457; // @[Mux.scala 31:69:@71.4]
  assign select_0 = valid_0_0 ? 4'h0 : _T_1458; // @[Mux.scala 31:69:@72.4]
  assign _GEN_1 = 4'h1 == select_0 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@74.4]
  assign _GEN_2 = 4'h2 == select_0 ? io_inData_2 : _GEN_1; // @[Switch.scala 33:19:@74.4]
  assign _GEN_3 = 4'h3 == select_0 ? io_inData_3 : _GEN_2; // @[Switch.scala 33:19:@74.4]
  assign _GEN_4 = 4'h4 == select_0 ? io_inData_4 : _GEN_3; // @[Switch.scala 33:19:@74.4]
  assign _GEN_5 = 4'h5 == select_0 ? io_inData_5 : _GEN_4; // @[Switch.scala 33:19:@74.4]
  assign _GEN_6 = 4'h6 == select_0 ? io_inData_6 : _GEN_5; // @[Switch.scala 33:19:@74.4]
  assign _GEN_7 = 4'h7 == select_0 ? io_inData_7 : _GEN_6; // @[Switch.scala 33:19:@74.4]
  assign _GEN_8 = 4'h8 == select_0 ? io_inData_8 : _GEN_7; // @[Switch.scala 33:19:@74.4]
  assign _GEN_9 = 4'h9 == select_0 ? io_inData_9 : _GEN_8; // @[Switch.scala 33:19:@74.4]
  assign _GEN_10 = 4'ha == select_0 ? io_inData_10 : _GEN_9; // @[Switch.scala 33:19:@74.4]
  assign _GEN_11 = 4'hb == select_0 ? io_inData_11 : _GEN_10; // @[Switch.scala 33:19:@74.4]
  assign _GEN_12 = 4'hc == select_0 ? io_inData_12 : _GEN_11; // @[Switch.scala 33:19:@74.4]
  assign _GEN_13 = 4'hd == select_0 ? io_inData_13 : _GEN_12; // @[Switch.scala 33:19:@74.4]
  assign _GEN_14 = 4'he == select_0 ? io_inData_14 : _GEN_13; // @[Switch.scala 33:19:@74.4]
  assign _T_1467 = {valid_0_7,valid_0_6,valid_0_5,valid_0_4,valid_0_3,valid_0_2,valid_0_1,valid_0_0}; // @[Switch.scala 34:32:@81.4]
  assign _T_1475 = {valid_0_15,valid_0_14,valid_0_13,valid_0_12,valid_0_11,valid_0_10,valid_0_9,valid_0_8,_T_1467}; // @[Switch.scala 34:32:@89.4]
  assign _T_1479 = io_inAddr_0 == 4'h1; // @[Switch.scala 30:53:@92.4]
  assign valid_1_0 = io_inValid_0 & _T_1479; // @[Switch.scala 30:36:@93.4]
  assign _T_1482 = io_inAddr_1 == 4'h1; // @[Switch.scala 30:53:@95.4]
  assign valid_1_1 = io_inValid_1 & _T_1482; // @[Switch.scala 30:36:@96.4]
  assign _T_1485 = io_inAddr_2 == 4'h1; // @[Switch.scala 30:53:@98.4]
  assign valid_1_2 = io_inValid_2 & _T_1485; // @[Switch.scala 30:36:@99.4]
  assign _T_1488 = io_inAddr_3 == 4'h1; // @[Switch.scala 30:53:@101.4]
  assign valid_1_3 = io_inValid_3 & _T_1488; // @[Switch.scala 30:36:@102.4]
  assign _T_1491 = io_inAddr_4 == 4'h1; // @[Switch.scala 30:53:@104.4]
  assign valid_1_4 = io_inValid_4 & _T_1491; // @[Switch.scala 30:36:@105.4]
  assign _T_1494 = io_inAddr_5 == 4'h1; // @[Switch.scala 30:53:@107.4]
  assign valid_1_5 = io_inValid_5 & _T_1494; // @[Switch.scala 30:36:@108.4]
  assign _T_1497 = io_inAddr_6 == 4'h1; // @[Switch.scala 30:53:@110.4]
  assign valid_1_6 = io_inValid_6 & _T_1497; // @[Switch.scala 30:36:@111.4]
  assign _T_1500 = io_inAddr_7 == 4'h1; // @[Switch.scala 30:53:@113.4]
  assign valid_1_7 = io_inValid_7 & _T_1500; // @[Switch.scala 30:36:@114.4]
  assign _T_1503 = io_inAddr_8 == 4'h1; // @[Switch.scala 30:53:@116.4]
  assign valid_1_8 = io_inValid_8 & _T_1503; // @[Switch.scala 30:36:@117.4]
  assign _T_1506 = io_inAddr_9 == 4'h1; // @[Switch.scala 30:53:@119.4]
  assign valid_1_9 = io_inValid_9 & _T_1506; // @[Switch.scala 30:36:@120.4]
  assign _T_1509 = io_inAddr_10 == 4'h1; // @[Switch.scala 30:53:@122.4]
  assign valid_1_10 = io_inValid_10 & _T_1509; // @[Switch.scala 30:36:@123.4]
  assign _T_1512 = io_inAddr_11 == 4'h1; // @[Switch.scala 30:53:@125.4]
  assign valid_1_11 = io_inValid_11 & _T_1512; // @[Switch.scala 30:36:@126.4]
  assign _T_1515 = io_inAddr_12 == 4'h1; // @[Switch.scala 30:53:@128.4]
  assign valid_1_12 = io_inValid_12 & _T_1515; // @[Switch.scala 30:36:@129.4]
  assign _T_1518 = io_inAddr_13 == 4'h1; // @[Switch.scala 30:53:@131.4]
  assign valid_1_13 = io_inValid_13 & _T_1518; // @[Switch.scala 30:36:@132.4]
  assign _T_1521 = io_inAddr_14 == 4'h1; // @[Switch.scala 30:53:@134.4]
  assign valid_1_14 = io_inValid_14 & _T_1521; // @[Switch.scala 30:36:@135.4]
  assign _T_1524 = io_inAddr_15 == 4'h1; // @[Switch.scala 30:53:@137.4]
  assign valid_1_15 = io_inValid_15 & _T_1524; // @[Switch.scala 30:36:@138.4]
  assign _T_1542 = valid_1_14 ? 4'he : 4'hf; // @[Mux.scala 31:69:@140.4]
  assign _T_1543 = valid_1_13 ? 4'hd : _T_1542; // @[Mux.scala 31:69:@141.4]
  assign _T_1544 = valid_1_12 ? 4'hc : _T_1543; // @[Mux.scala 31:69:@142.4]
  assign _T_1545 = valid_1_11 ? 4'hb : _T_1544; // @[Mux.scala 31:69:@143.4]
  assign _T_1546 = valid_1_10 ? 4'ha : _T_1545; // @[Mux.scala 31:69:@144.4]
  assign _T_1547 = valid_1_9 ? 4'h9 : _T_1546; // @[Mux.scala 31:69:@145.4]
  assign _T_1548 = valid_1_8 ? 4'h8 : _T_1547; // @[Mux.scala 31:69:@146.4]
  assign _T_1549 = valid_1_7 ? 4'h7 : _T_1548; // @[Mux.scala 31:69:@147.4]
  assign _T_1550 = valid_1_6 ? 4'h6 : _T_1549; // @[Mux.scala 31:69:@148.4]
  assign _T_1551 = valid_1_5 ? 4'h5 : _T_1550; // @[Mux.scala 31:69:@149.4]
  assign _T_1552 = valid_1_4 ? 4'h4 : _T_1551; // @[Mux.scala 31:69:@150.4]
  assign _T_1553 = valid_1_3 ? 4'h3 : _T_1552; // @[Mux.scala 31:69:@151.4]
  assign _T_1554 = valid_1_2 ? 4'h2 : _T_1553; // @[Mux.scala 31:69:@152.4]
  assign _T_1555 = valid_1_1 ? 4'h1 : _T_1554; // @[Mux.scala 31:69:@153.4]
  assign select_1 = valid_1_0 ? 4'h0 : _T_1555; // @[Mux.scala 31:69:@154.4]
  assign _GEN_17 = 4'h1 == select_1 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@156.4]
  assign _GEN_18 = 4'h2 == select_1 ? io_inData_2 : _GEN_17; // @[Switch.scala 33:19:@156.4]
  assign _GEN_19 = 4'h3 == select_1 ? io_inData_3 : _GEN_18; // @[Switch.scala 33:19:@156.4]
  assign _GEN_20 = 4'h4 == select_1 ? io_inData_4 : _GEN_19; // @[Switch.scala 33:19:@156.4]
  assign _GEN_21 = 4'h5 == select_1 ? io_inData_5 : _GEN_20; // @[Switch.scala 33:19:@156.4]
  assign _GEN_22 = 4'h6 == select_1 ? io_inData_6 : _GEN_21; // @[Switch.scala 33:19:@156.4]
  assign _GEN_23 = 4'h7 == select_1 ? io_inData_7 : _GEN_22; // @[Switch.scala 33:19:@156.4]
  assign _GEN_24 = 4'h8 == select_1 ? io_inData_8 : _GEN_23; // @[Switch.scala 33:19:@156.4]
  assign _GEN_25 = 4'h9 == select_1 ? io_inData_9 : _GEN_24; // @[Switch.scala 33:19:@156.4]
  assign _GEN_26 = 4'ha == select_1 ? io_inData_10 : _GEN_25; // @[Switch.scala 33:19:@156.4]
  assign _GEN_27 = 4'hb == select_1 ? io_inData_11 : _GEN_26; // @[Switch.scala 33:19:@156.4]
  assign _GEN_28 = 4'hc == select_1 ? io_inData_12 : _GEN_27; // @[Switch.scala 33:19:@156.4]
  assign _GEN_29 = 4'hd == select_1 ? io_inData_13 : _GEN_28; // @[Switch.scala 33:19:@156.4]
  assign _GEN_30 = 4'he == select_1 ? io_inData_14 : _GEN_29; // @[Switch.scala 33:19:@156.4]
  assign _T_1564 = {valid_1_7,valid_1_6,valid_1_5,valid_1_4,valid_1_3,valid_1_2,valid_1_1,valid_1_0}; // @[Switch.scala 34:32:@163.4]
  assign _T_1572 = {valid_1_15,valid_1_14,valid_1_13,valid_1_12,valid_1_11,valid_1_10,valid_1_9,valid_1_8,_T_1564}; // @[Switch.scala 34:32:@171.4]
  assign _T_1576 = io_inAddr_0 == 4'h2; // @[Switch.scala 30:53:@174.4]
  assign valid_2_0 = io_inValid_0 & _T_1576; // @[Switch.scala 30:36:@175.4]
  assign _T_1579 = io_inAddr_1 == 4'h2; // @[Switch.scala 30:53:@177.4]
  assign valid_2_1 = io_inValid_1 & _T_1579; // @[Switch.scala 30:36:@178.4]
  assign _T_1582 = io_inAddr_2 == 4'h2; // @[Switch.scala 30:53:@180.4]
  assign valid_2_2 = io_inValid_2 & _T_1582; // @[Switch.scala 30:36:@181.4]
  assign _T_1585 = io_inAddr_3 == 4'h2; // @[Switch.scala 30:53:@183.4]
  assign valid_2_3 = io_inValid_3 & _T_1585; // @[Switch.scala 30:36:@184.4]
  assign _T_1588 = io_inAddr_4 == 4'h2; // @[Switch.scala 30:53:@186.4]
  assign valid_2_4 = io_inValid_4 & _T_1588; // @[Switch.scala 30:36:@187.4]
  assign _T_1591 = io_inAddr_5 == 4'h2; // @[Switch.scala 30:53:@189.4]
  assign valid_2_5 = io_inValid_5 & _T_1591; // @[Switch.scala 30:36:@190.4]
  assign _T_1594 = io_inAddr_6 == 4'h2; // @[Switch.scala 30:53:@192.4]
  assign valid_2_6 = io_inValid_6 & _T_1594; // @[Switch.scala 30:36:@193.4]
  assign _T_1597 = io_inAddr_7 == 4'h2; // @[Switch.scala 30:53:@195.4]
  assign valid_2_7 = io_inValid_7 & _T_1597; // @[Switch.scala 30:36:@196.4]
  assign _T_1600 = io_inAddr_8 == 4'h2; // @[Switch.scala 30:53:@198.4]
  assign valid_2_8 = io_inValid_8 & _T_1600; // @[Switch.scala 30:36:@199.4]
  assign _T_1603 = io_inAddr_9 == 4'h2; // @[Switch.scala 30:53:@201.4]
  assign valid_2_9 = io_inValid_9 & _T_1603; // @[Switch.scala 30:36:@202.4]
  assign _T_1606 = io_inAddr_10 == 4'h2; // @[Switch.scala 30:53:@204.4]
  assign valid_2_10 = io_inValid_10 & _T_1606; // @[Switch.scala 30:36:@205.4]
  assign _T_1609 = io_inAddr_11 == 4'h2; // @[Switch.scala 30:53:@207.4]
  assign valid_2_11 = io_inValid_11 & _T_1609; // @[Switch.scala 30:36:@208.4]
  assign _T_1612 = io_inAddr_12 == 4'h2; // @[Switch.scala 30:53:@210.4]
  assign valid_2_12 = io_inValid_12 & _T_1612; // @[Switch.scala 30:36:@211.4]
  assign _T_1615 = io_inAddr_13 == 4'h2; // @[Switch.scala 30:53:@213.4]
  assign valid_2_13 = io_inValid_13 & _T_1615; // @[Switch.scala 30:36:@214.4]
  assign _T_1618 = io_inAddr_14 == 4'h2; // @[Switch.scala 30:53:@216.4]
  assign valid_2_14 = io_inValid_14 & _T_1618; // @[Switch.scala 30:36:@217.4]
  assign _T_1621 = io_inAddr_15 == 4'h2; // @[Switch.scala 30:53:@219.4]
  assign valid_2_15 = io_inValid_15 & _T_1621; // @[Switch.scala 30:36:@220.4]
  assign _T_1639 = valid_2_14 ? 4'he : 4'hf; // @[Mux.scala 31:69:@222.4]
  assign _T_1640 = valid_2_13 ? 4'hd : _T_1639; // @[Mux.scala 31:69:@223.4]
  assign _T_1641 = valid_2_12 ? 4'hc : _T_1640; // @[Mux.scala 31:69:@224.4]
  assign _T_1642 = valid_2_11 ? 4'hb : _T_1641; // @[Mux.scala 31:69:@225.4]
  assign _T_1643 = valid_2_10 ? 4'ha : _T_1642; // @[Mux.scala 31:69:@226.4]
  assign _T_1644 = valid_2_9 ? 4'h9 : _T_1643; // @[Mux.scala 31:69:@227.4]
  assign _T_1645 = valid_2_8 ? 4'h8 : _T_1644; // @[Mux.scala 31:69:@228.4]
  assign _T_1646 = valid_2_7 ? 4'h7 : _T_1645; // @[Mux.scala 31:69:@229.4]
  assign _T_1647 = valid_2_6 ? 4'h6 : _T_1646; // @[Mux.scala 31:69:@230.4]
  assign _T_1648 = valid_2_5 ? 4'h5 : _T_1647; // @[Mux.scala 31:69:@231.4]
  assign _T_1649 = valid_2_4 ? 4'h4 : _T_1648; // @[Mux.scala 31:69:@232.4]
  assign _T_1650 = valid_2_3 ? 4'h3 : _T_1649; // @[Mux.scala 31:69:@233.4]
  assign _T_1651 = valid_2_2 ? 4'h2 : _T_1650; // @[Mux.scala 31:69:@234.4]
  assign _T_1652 = valid_2_1 ? 4'h1 : _T_1651; // @[Mux.scala 31:69:@235.4]
  assign select_2 = valid_2_0 ? 4'h0 : _T_1652; // @[Mux.scala 31:69:@236.4]
  assign _GEN_33 = 4'h1 == select_2 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@238.4]
  assign _GEN_34 = 4'h2 == select_2 ? io_inData_2 : _GEN_33; // @[Switch.scala 33:19:@238.4]
  assign _GEN_35 = 4'h3 == select_2 ? io_inData_3 : _GEN_34; // @[Switch.scala 33:19:@238.4]
  assign _GEN_36 = 4'h4 == select_2 ? io_inData_4 : _GEN_35; // @[Switch.scala 33:19:@238.4]
  assign _GEN_37 = 4'h5 == select_2 ? io_inData_5 : _GEN_36; // @[Switch.scala 33:19:@238.4]
  assign _GEN_38 = 4'h6 == select_2 ? io_inData_6 : _GEN_37; // @[Switch.scala 33:19:@238.4]
  assign _GEN_39 = 4'h7 == select_2 ? io_inData_7 : _GEN_38; // @[Switch.scala 33:19:@238.4]
  assign _GEN_40 = 4'h8 == select_2 ? io_inData_8 : _GEN_39; // @[Switch.scala 33:19:@238.4]
  assign _GEN_41 = 4'h9 == select_2 ? io_inData_9 : _GEN_40; // @[Switch.scala 33:19:@238.4]
  assign _GEN_42 = 4'ha == select_2 ? io_inData_10 : _GEN_41; // @[Switch.scala 33:19:@238.4]
  assign _GEN_43 = 4'hb == select_2 ? io_inData_11 : _GEN_42; // @[Switch.scala 33:19:@238.4]
  assign _GEN_44 = 4'hc == select_2 ? io_inData_12 : _GEN_43; // @[Switch.scala 33:19:@238.4]
  assign _GEN_45 = 4'hd == select_2 ? io_inData_13 : _GEN_44; // @[Switch.scala 33:19:@238.4]
  assign _GEN_46 = 4'he == select_2 ? io_inData_14 : _GEN_45; // @[Switch.scala 33:19:@238.4]
  assign _T_1661 = {valid_2_7,valid_2_6,valid_2_5,valid_2_4,valid_2_3,valid_2_2,valid_2_1,valid_2_0}; // @[Switch.scala 34:32:@245.4]
  assign _T_1669 = {valid_2_15,valid_2_14,valid_2_13,valid_2_12,valid_2_11,valid_2_10,valid_2_9,valid_2_8,_T_1661}; // @[Switch.scala 34:32:@253.4]
  assign _T_1673 = io_inAddr_0 == 4'h3; // @[Switch.scala 30:53:@256.4]
  assign valid_3_0 = io_inValid_0 & _T_1673; // @[Switch.scala 30:36:@257.4]
  assign _T_1676 = io_inAddr_1 == 4'h3; // @[Switch.scala 30:53:@259.4]
  assign valid_3_1 = io_inValid_1 & _T_1676; // @[Switch.scala 30:36:@260.4]
  assign _T_1679 = io_inAddr_2 == 4'h3; // @[Switch.scala 30:53:@262.4]
  assign valid_3_2 = io_inValid_2 & _T_1679; // @[Switch.scala 30:36:@263.4]
  assign _T_1682 = io_inAddr_3 == 4'h3; // @[Switch.scala 30:53:@265.4]
  assign valid_3_3 = io_inValid_3 & _T_1682; // @[Switch.scala 30:36:@266.4]
  assign _T_1685 = io_inAddr_4 == 4'h3; // @[Switch.scala 30:53:@268.4]
  assign valid_3_4 = io_inValid_4 & _T_1685; // @[Switch.scala 30:36:@269.4]
  assign _T_1688 = io_inAddr_5 == 4'h3; // @[Switch.scala 30:53:@271.4]
  assign valid_3_5 = io_inValid_5 & _T_1688; // @[Switch.scala 30:36:@272.4]
  assign _T_1691 = io_inAddr_6 == 4'h3; // @[Switch.scala 30:53:@274.4]
  assign valid_3_6 = io_inValid_6 & _T_1691; // @[Switch.scala 30:36:@275.4]
  assign _T_1694 = io_inAddr_7 == 4'h3; // @[Switch.scala 30:53:@277.4]
  assign valid_3_7 = io_inValid_7 & _T_1694; // @[Switch.scala 30:36:@278.4]
  assign _T_1697 = io_inAddr_8 == 4'h3; // @[Switch.scala 30:53:@280.4]
  assign valid_3_8 = io_inValid_8 & _T_1697; // @[Switch.scala 30:36:@281.4]
  assign _T_1700 = io_inAddr_9 == 4'h3; // @[Switch.scala 30:53:@283.4]
  assign valid_3_9 = io_inValid_9 & _T_1700; // @[Switch.scala 30:36:@284.4]
  assign _T_1703 = io_inAddr_10 == 4'h3; // @[Switch.scala 30:53:@286.4]
  assign valid_3_10 = io_inValid_10 & _T_1703; // @[Switch.scala 30:36:@287.4]
  assign _T_1706 = io_inAddr_11 == 4'h3; // @[Switch.scala 30:53:@289.4]
  assign valid_3_11 = io_inValid_11 & _T_1706; // @[Switch.scala 30:36:@290.4]
  assign _T_1709 = io_inAddr_12 == 4'h3; // @[Switch.scala 30:53:@292.4]
  assign valid_3_12 = io_inValid_12 & _T_1709; // @[Switch.scala 30:36:@293.4]
  assign _T_1712 = io_inAddr_13 == 4'h3; // @[Switch.scala 30:53:@295.4]
  assign valid_3_13 = io_inValid_13 & _T_1712; // @[Switch.scala 30:36:@296.4]
  assign _T_1715 = io_inAddr_14 == 4'h3; // @[Switch.scala 30:53:@298.4]
  assign valid_3_14 = io_inValid_14 & _T_1715; // @[Switch.scala 30:36:@299.4]
  assign _T_1718 = io_inAddr_15 == 4'h3; // @[Switch.scala 30:53:@301.4]
  assign valid_3_15 = io_inValid_15 & _T_1718; // @[Switch.scala 30:36:@302.4]
  assign _T_1736 = valid_3_14 ? 4'he : 4'hf; // @[Mux.scala 31:69:@304.4]
  assign _T_1737 = valid_3_13 ? 4'hd : _T_1736; // @[Mux.scala 31:69:@305.4]
  assign _T_1738 = valid_3_12 ? 4'hc : _T_1737; // @[Mux.scala 31:69:@306.4]
  assign _T_1739 = valid_3_11 ? 4'hb : _T_1738; // @[Mux.scala 31:69:@307.4]
  assign _T_1740 = valid_3_10 ? 4'ha : _T_1739; // @[Mux.scala 31:69:@308.4]
  assign _T_1741 = valid_3_9 ? 4'h9 : _T_1740; // @[Mux.scala 31:69:@309.4]
  assign _T_1742 = valid_3_8 ? 4'h8 : _T_1741; // @[Mux.scala 31:69:@310.4]
  assign _T_1743 = valid_3_7 ? 4'h7 : _T_1742; // @[Mux.scala 31:69:@311.4]
  assign _T_1744 = valid_3_6 ? 4'h6 : _T_1743; // @[Mux.scala 31:69:@312.4]
  assign _T_1745 = valid_3_5 ? 4'h5 : _T_1744; // @[Mux.scala 31:69:@313.4]
  assign _T_1746 = valid_3_4 ? 4'h4 : _T_1745; // @[Mux.scala 31:69:@314.4]
  assign _T_1747 = valid_3_3 ? 4'h3 : _T_1746; // @[Mux.scala 31:69:@315.4]
  assign _T_1748 = valid_3_2 ? 4'h2 : _T_1747; // @[Mux.scala 31:69:@316.4]
  assign _T_1749 = valid_3_1 ? 4'h1 : _T_1748; // @[Mux.scala 31:69:@317.4]
  assign select_3 = valid_3_0 ? 4'h0 : _T_1749; // @[Mux.scala 31:69:@318.4]
  assign _GEN_49 = 4'h1 == select_3 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@320.4]
  assign _GEN_50 = 4'h2 == select_3 ? io_inData_2 : _GEN_49; // @[Switch.scala 33:19:@320.4]
  assign _GEN_51 = 4'h3 == select_3 ? io_inData_3 : _GEN_50; // @[Switch.scala 33:19:@320.4]
  assign _GEN_52 = 4'h4 == select_3 ? io_inData_4 : _GEN_51; // @[Switch.scala 33:19:@320.4]
  assign _GEN_53 = 4'h5 == select_3 ? io_inData_5 : _GEN_52; // @[Switch.scala 33:19:@320.4]
  assign _GEN_54 = 4'h6 == select_3 ? io_inData_6 : _GEN_53; // @[Switch.scala 33:19:@320.4]
  assign _GEN_55 = 4'h7 == select_3 ? io_inData_7 : _GEN_54; // @[Switch.scala 33:19:@320.4]
  assign _GEN_56 = 4'h8 == select_3 ? io_inData_8 : _GEN_55; // @[Switch.scala 33:19:@320.4]
  assign _GEN_57 = 4'h9 == select_3 ? io_inData_9 : _GEN_56; // @[Switch.scala 33:19:@320.4]
  assign _GEN_58 = 4'ha == select_3 ? io_inData_10 : _GEN_57; // @[Switch.scala 33:19:@320.4]
  assign _GEN_59 = 4'hb == select_3 ? io_inData_11 : _GEN_58; // @[Switch.scala 33:19:@320.4]
  assign _GEN_60 = 4'hc == select_3 ? io_inData_12 : _GEN_59; // @[Switch.scala 33:19:@320.4]
  assign _GEN_61 = 4'hd == select_3 ? io_inData_13 : _GEN_60; // @[Switch.scala 33:19:@320.4]
  assign _GEN_62 = 4'he == select_3 ? io_inData_14 : _GEN_61; // @[Switch.scala 33:19:@320.4]
  assign _T_1758 = {valid_3_7,valid_3_6,valid_3_5,valid_3_4,valid_3_3,valid_3_2,valid_3_1,valid_3_0}; // @[Switch.scala 34:32:@327.4]
  assign _T_1766 = {valid_3_15,valid_3_14,valid_3_13,valid_3_12,valid_3_11,valid_3_10,valid_3_9,valid_3_8,_T_1758}; // @[Switch.scala 34:32:@335.4]
  assign _T_1770 = io_inAddr_0 == 4'h4; // @[Switch.scala 30:53:@338.4]
  assign valid_4_0 = io_inValid_0 & _T_1770; // @[Switch.scala 30:36:@339.4]
  assign _T_1773 = io_inAddr_1 == 4'h4; // @[Switch.scala 30:53:@341.4]
  assign valid_4_1 = io_inValid_1 & _T_1773; // @[Switch.scala 30:36:@342.4]
  assign _T_1776 = io_inAddr_2 == 4'h4; // @[Switch.scala 30:53:@344.4]
  assign valid_4_2 = io_inValid_2 & _T_1776; // @[Switch.scala 30:36:@345.4]
  assign _T_1779 = io_inAddr_3 == 4'h4; // @[Switch.scala 30:53:@347.4]
  assign valid_4_3 = io_inValid_3 & _T_1779; // @[Switch.scala 30:36:@348.4]
  assign _T_1782 = io_inAddr_4 == 4'h4; // @[Switch.scala 30:53:@350.4]
  assign valid_4_4 = io_inValid_4 & _T_1782; // @[Switch.scala 30:36:@351.4]
  assign _T_1785 = io_inAddr_5 == 4'h4; // @[Switch.scala 30:53:@353.4]
  assign valid_4_5 = io_inValid_5 & _T_1785; // @[Switch.scala 30:36:@354.4]
  assign _T_1788 = io_inAddr_6 == 4'h4; // @[Switch.scala 30:53:@356.4]
  assign valid_4_6 = io_inValid_6 & _T_1788; // @[Switch.scala 30:36:@357.4]
  assign _T_1791 = io_inAddr_7 == 4'h4; // @[Switch.scala 30:53:@359.4]
  assign valid_4_7 = io_inValid_7 & _T_1791; // @[Switch.scala 30:36:@360.4]
  assign _T_1794 = io_inAddr_8 == 4'h4; // @[Switch.scala 30:53:@362.4]
  assign valid_4_8 = io_inValid_8 & _T_1794; // @[Switch.scala 30:36:@363.4]
  assign _T_1797 = io_inAddr_9 == 4'h4; // @[Switch.scala 30:53:@365.4]
  assign valid_4_9 = io_inValid_9 & _T_1797; // @[Switch.scala 30:36:@366.4]
  assign _T_1800 = io_inAddr_10 == 4'h4; // @[Switch.scala 30:53:@368.4]
  assign valid_4_10 = io_inValid_10 & _T_1800; // @[Switch.scala 30:36:@369.4]
  assign _T_1803 = io_inAddr_11 == 4'h4; // @[Switch.scala 30:53:@371.4]
  assign valid_4_11 = io_inValid_11 & _T_1803; // @[Switch.scala 30:36:@372.4]
  assign _T_1806 = io_inAddr_12 == 4'h4; // @[Switch.scala 30:53:@374.4]
  assign valid_4_12 = io_inValid_12 & _T_1806; // @[Switch.scala 30:36:@375.4]
  assign _T_1809 = io_inAddr_13 == 4'h4; // @[Switch.scala 30:53:@377.4]
  assign valid_4_13 = io_inValid_13 & _T_1809; // @[Switch.scala 30:36:@378.4]
  assign _T_1812 = io_inAddr_14 == 4'h4; // @[Switch.scala 30:53:@380.4]
  assign valid_4_14 = io_inValid_14 & _T_1812; // @[Switch.scala 30:36:@381.4]
  assign _T_1815 = io_inAddr_15 == 4'h4; // @[Switch.scala 30:53:@383.4]
  assign valid_4_15 = io_inValid_15 & _T_1815; // @[Switch.scala 30:36:@384.4]
  assign _T_1833 = valid_4_14 ? 4'he : 4'hf; // @[Mux.scala 31:69:@386.4]
  assign _T_1834 = valid_4_13 ? 4'hd : _T_1833; // @[Mux.scala 31:69:@387.4]
  assign _T_1835 = valid_4_12 ? 4'hc : _T_1834; // @[Mux.scala 31:69:@388.4]
  assign _T_1836 = valid_4_11 ? 4'hb : _T_1835; // @[Mux.scala 31:69:@389.4]
  assign _T_1837 = valid_4_10 ? 4'ha : _T_1836; // @[Mux.scala 31:69:@390.4]
  assign _T_1838 = valid_4_9 ? 4'h9 : _T_1837; // @[Mux.scala 31:69:@391.4]
  assign _T_1839 = valid_4_8 ? 4'h8 : _T_1838; // @[Mux.scala 31:69:@392.4]
  assign _T_1840 = valid_4_7 ? 4'h7 : _T_1839; // @[Mux.scala 31:69:@393.4]
  assign _T_1841 = valid_4_6 ? 4'h6 : _T_1840; // @[Mux.scala 31:69:@394.4]
  assign _T_1842 = valid_4_5 ? 4'h5 : _T_1841; // @[Mux.scala 31:69:@395.4]
  assign _T_1843 = valid_4_4 ? 4'h4 : _T_1842; // @[Mux.scala 31:69:@396.4]
  assign _T_1844 = valid_4_3 ? 4'h3 : _T_1843; // @[Mux.scala 31:69:@397.4]
  assign _T_1845 = valid_4_2 ? 4'h2 : _T_1844; // @[Mux.scala 31:69:@398.4]
  assign _T_1846 = valid_4_1 ? 4'h1 : _T_1845; // @[Mux.scala 31:69:@399.4]
  assign select_4 = valid_4_0 ? 4'h0 : _T_1846; // @[Mux.scala 31:69:@400.4]
  assign _GEN_65 = 4'h1 == select_4 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@402.4]
  assign _GEN_66 = 4'h2 == select_4 ? io_inData_2 : _GEN_65; // @[Switch.scala 33:19:@402.4]
  assign _GEN_67 = 4'h3 == select_4 ? io_inData_3 : _GEN_66; // @[Switch.scala 33:19:@402.4]
  assign _GEN_68 = 4'h4 == select_4 ? io_inData_4 : _GEN_67; // @[Switch.scala 33:19:@402.4]
  assign _GEN_69 = 4'h5 == select_4 ? io_inData_5 : _GEN_68; // @[Switch.scala 33:19:@402.4]
  assign _GEN_70 = 4'h6 == select_4 ? io_inData_6 : _GEN_69; // @[Switch.scala 33:19:@402.4]
  assign _GEN_71 = 4'h7 == select_4 ? io_inData_7 : _GEN_70; // @[Switch.scala 33:19:@402.4]
  assign _GEN_72 = 4'h8 == select_4 ? io_inData_8 : _GEN_71; // @[Switch.scala 33:19:@402.4]
  assign _GEN_73 = 4'h9 == select_4 ? io_inData_9 : _GEN_72; // @[Switch.scala 33:19:@402.4]
  assign _GEN_74 = 4'ha == select_4 ? io_inData_10 : _GEN_73; // @[Switch.scala 33:19:@402.4]
  assign _GEN_75 = 4'hb == select_4 ? io_inData_11 : _GEN_74; // @[Switch.scala 33:19:@402.4]
  assign _GEN_76 = 4'hc == select_4 ? io_inData_12 : _GEN_75; // @[Switch.scala 33:19:@402.4]
  assign _GEN_77 = 4'hd == select_4 ? io_inData_13 : _GEN_76; // @[Switch.scala 33:19:@402.4]
  assign _GEN_78 = 4'he == select_4 ? io_inData_14 : _GEN_77; // @[Switch.scala 33:19:@402.4]
  assign _T_1855 = {valid_4_7,valid_4_6,valid_4_5,valid_4_4,valid_4_3,valid_4_2,valid_4_1,valid_4_0}; // @[Switch.scala 34:32:@409.4]
  assign _T_1863 = {valid_4_15,valid_4_14,valid_4_13,valid_4_12,valid_4_11,valid_4_10,valid_4_9,valid_4_8,_T_1855}; // @[Switch.scala 34:32:@417.4]
  assign _T_1867 = io_inAddr_0 == 4'h5; // @[Switch.scala 30:53:@420.4]
  assign valid_5_0 = io_inValid_0 & _T_1867; // @[Switch.scala 30:36:@421.4]
  assign _T_1870 = io_inAddr_1 == 4'h5; // @[Switch.scala 30:53:@423.4]
  assign valid_5_1 = io_inValid_1 & _T_1870; // @[Switch.scala 30:36:@424.4]
  assign _T_1873 = io_inAddr_2 == 4'h5; // @[Switch.scala 30:53:@426.4]
  assign valid_5_2 = io_inValid_2 & _T_1873; // @[Switch.scala 30:36:@427.4]
  assign _T_1876 = io_inAddr_3 == 4'h5; // @[Switch.scala 30:53:@429.4]
  assign valid_5_3 = io_inValid_3 & _T_1876; // @[Switch.scala 30:36:@430.4]
  assign _T_1879 = io_inAddr_4 == 4'h5; // @[Switch.scala 30:53:@432.4]
  assign valid_5_4 = io_inValid_4 & _T_1879; // @[Switch.scala 30:36:@433.4]
  assign _T_1882 = io_inAddr_5 == 4'h5; // @[Switch.scala 30:53:@435.4]
  assign valid_5_5 = io_inValid_5 & _T_1882; // @[Switch.scala 30:36:@436.4]
  assign _T_1885 = io_inAddr_6 == 4'h5; // @[Switch.scala 30:53:@438.4]
  assign valid_5_6 = io_inValid_6 & _T_1885; // @[Switch.scala 30:36:@439.4]
  assign _T_1888 = io_inAddr_7 == 4'h5; // @[Switch.scala 30:53:@441.4]
  assign valid_5_7 = io_inValid_7 & _T_1888; // @[Switch.scala 30:36:@442.4]
  assign _T_1891 = io_inAddr_8 == 4'h5; // @[Switch.scala 30:53:@444.4]
  assign valid_5_8 = io_inValid_8 & _T_1891; // @[Switch.scala 30:36:@445.4]
  assign _T_1894 = io_inAddr_9 == 4'h5; // @[Switch.scala 30:53:@447.4]
  assign valid_5_9 = io_inValid_9 & _T_1894; // @[Switch.scala 30:36:@448.4]
  assign _T_1897 = io_inAddr_10 == 4'h5; // @[Switch.scala 30:53:@450.4]
  assign valid_5_10 = io_inValid_10 & _T_1897; // @[Switch.scala 30:36:@451.4]
  assign _T_1900 = io_inAddr_11 == 4'h5; // @[Switch.scala 30:53:@453.4]
  assign valid_5_11 = io_inValid_11 & _T_1900; // @[Switch.scala 30:36:@454.4]
  assign _T_1903 = io_inAddr_12 == 4'h5; // @[Switch.scala 30:53:@456.4]
  assign valid_5_12 = io_inValid_12 & _T_1903; // @[Switch.scala 30:36:@457.4]
  assign _T_1906 = io_inAddr_13 == 4'h5; // @[Switch.scala 30:53:@459.4]
  assign valid_5_13 = io_inValid_13 & _T_1906; // @[Switch.scala 30:36:@460.4]
  assign _T_1909 = io_inAddr_14 == 4'h5; // @[Switch.scala 30:53:@462.4]
  assign valid_5_14 = io_inValid_14 & _T_1909; // @[Switch.scala 30:36:@463.4]
  assign _T_1912 = io_inAddr_15 == 4'h5; // @[Switch.scala 30:53:@465.4]
  assign valid_5_15 = io_inValid_15 & _T_1912; // @[Switch.scala 30:36:@466.4]
  assign _T_1930 = valid_5_14 ? 4'he : 4'hf; // @[Mux.scala 31:69:@468.4]
  assign _T_1931 = valid_5_13 ? 4'hd : _T_1930; // @[Mux.scala 31:69:@469.4]
  assign _T_1932 = valid_5_12 ? 4'hc : _T_1931; // @[Mux.scala 31:69:@470.4]
  assign _T_1933 = valid_5_11 ? 4'hb : _T_1932; // @[Mux.scala 31:69:@471.4]
  assign _T_1934 = valid_5_10 ? 4'ha : _T_1933; // @[Mux.scala 31:69:@472.4]
  assign _T_1935 = valid_5_9 ? 4'h9 : _T_1934; // @[Mux.scala 31:69:@473.4]
  assign _T_1936 = valid_5_8 ? 4'h8 : _T_1935; // @[Mux.scala 31:69:@474.4]
  assign _T_1937 = valid_5_7 ? 4'h7 : _T_1936; // @[Mux.scala 31:69:@475.4]
  assign _T_1938 = valid_5_6 ? 4'h6 : _T_1937; // @[Mux.scala 31:69:@476.4]
  assign _T_1939 = valid_5_5 ? 4'h5 : _T_1938; // @[Mux.scala 31:69:@477.4]
  assign _T_1940 = valid_5_4 ? 4'h4 : _T_1939; // @[Mux.scala 31:69:@478.4]
  assign _T_1941 = valid_5_3 ? 4'h3 : _T_1940; // @[Mux.scala 31:69:@479.4]
  assign _T_1942 = valid_5_2 ? 4'h2 : _T_1941; // @[Mux.scala 31:69:@480.4]
  assign _T_1943 = valid_5_1 ? 4'h1 : _T_1942; // @[Mux.scala 31:69:@481.4]
  assign select_5 = valid_5_0 ? 4'h0 : _T_1943; // @[Mux.scala 31:69:@482.4]
  assign _GEN_81 = 4'h1 == select_5 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@484.4]
  assign _GEN_82 = 4'h2 == select_5 ? io_inData_2 : _GEN_81; // @[Switch.scala 33:19:@484.4]
  assign _GEN_83 = 4'h3 == select_5 ? io_inData_3 : _GEN_82; // @[Switch.scala 33:19:@484.4]
  assign _GEN_84 = 4'h4 == select_5 ? io_inData_4 : _GEN_83; // @[Switch.scala 33:19:@484.4]
  assign _GEN_85 = 4'h5 == select_5 ? io_inData_5 : _GEN_84; // @[Switch.scala 33:19:@484.4]
  assign _GEN_86 = 4'h6 == select_5 ? io_inData_6 : _GEN_85; // @[Switch.scala 33:19:@484.4]
  assign _GEN_87 = 4'h7 == select_5 ? io_inData_7 : _GEN_86; // @[Switch.scala 33:19:@484.4]
  assign _GEN_88 = 4'h8 == select_5 ? io_inData_8 : _GEN_87; // @[Switch.scala 33:19:@484.4]
  assign _GEN_89 = 4'h9 == select_5 ? io_inData_9 : _GEN_88; // @[Switch.scala 33:19:@484.4]
  assign _GEN_90 = 4'ha == select_5 ? io_inData_10 : _GEN_89; // @[Switch.scala 33:19:@484.4]
  assign _GEN_91 = 4'hb == select_5 ? io_inData_11 : _GEN_90; // @[Switch.scala 33:19:@484.4]
  assign _GEN_92 = 4'hc == select_5 ? io_inData_12 : _GEN_91; // @[Switch.scala 33:19:@484.4]
  assign _GEN_93 = 4'hd == select_5 ? io_inData_13 : _GEN_92; // @[Switch.scala 33:19:@484.4]
  assign _GEN_94 = 4'he == select_5 ? io_inData_14 : _GEN_93; // @[Switch.scala 33:19:@484.4]
  assign _T_1952 = {valid_5_7,valid_5_6,valid_5_5,valid_5_4,valid_5_3,valid_5_2,valid_5_1,valid_5_0}; // @[Switch.scala 34:32:@491.4]
  assign _T_1960 = {valid_5_15,valid_5_14,valid_5_13,valid_5_12,valid_5_11,valid_5_10,valid_5_9,valid_5_8,_T_1952}; // @[Switch.scala 34:32:@499.4]
  assign _T_1964 = io_inAddr_0 == 4'h6; // @[Switch.scala 30:53:@502.4]
  assign valid_6_0 = io_inValid_0 & _T_1964; // @[Switch.scala 30:36:@503.4]
  assign _T_1967 = io_inAddr_1 == 4'h6; // @[Switch.scala 30:53:@505.4]
  assign valid_6_1 = io_inValid_1 & _T_1967; // @[Switch.scala 30:36:@506.4]
  assign _T_1970 = io_inAddr_2 == 4'h6; // @[Switch.scala 30:53:@508.4]
  assign valid_6_2 = io_inValid_2 & _T_1970; // @[Switch.scala 30:36:@509.4]
  assign _T_1973 = io_inAddr_3 == 4'h6; // @[Switch.scala 30:53:@511.4]
  assign valid_6_3 = io_inValid_3 & _T_1973; // @[Switch.scala 30:36:@512.4]
  assign _T_1976 = io_inAddr_4 == 4'h6; // @[Switch.scala 30:53:@514.4]
  assign valid_6_4 = io_inValid_4 & _T_1976; // @[Switch.scala 30:36:@515.4]
  assign _T_1979 = io_inAddr_5 == 4'h6; // @[Switch.scala 30:53:@517.4]
  assign valid_6_5 = io_inValid_5 & _T_1979; // @[Switch.scala 30:36:@518.4]
  assign _T_1982 = io_inAddr_6 == 4'h6; // @[Switch.scala 30:53:@520.4]
  assign valid_6_6 = io_inValid_6 & _T_1982; // @[Switch.scala 30:36:@521.4]
  assign _T_1985 = io_inAddr_7 == 4'h6; // @[Switch.scala 30:53:@523.4]
  assign valid_6_7 = io_inValid_7 & _T_1985; // @[Switch.scala 30:36:@524.4]
  assign _T_1988 = io_inAddr_8 == 4'h6; // @[Switch.scala 30:53:@526.4]
  assign valid_6_8 = io_inValid_8 & _T_1988; // @[Switch.scala 30:36:@527.4]
  assign _T_1991 = io_inAddr_9 == 4'h6; // @[Switch.scala 30:53:@529.4]
  assign valid_6_9 = io_inValid_9 & _T_1991; // @[Switch.scala 30:36:@530.4]
  assign _T_1994 = io_inAddr_10 == 4'h6; // @[Switch.scala 30:53:@532.4]
  assign valid_6_10 = io_inValid_10 & _T_1994; // @[Switch.scala 30:36:@533.4]
  assign _T_1997 = io_inAddr_11 == 4'h6; // @[Switch.scala 30:53:@535.4]
  assign valid_6_11 = io_inValid_11 & _T_1997; // @[Switch.scala 30:36:@536.4]
  assign _T_2000 = io_inAddr_12 == 4'h6; // @[Switch.scala 30:53:@538.4]
  assign valid_6_12 = io_inValid_12 & _T_2000; // @[Switch.scala 30:36:@539.4]
  assign _T_2003 = io_inAddr_13 == 4'h6; // @[Switch.scala 30:53:@541.4]
  assign valid_6_13 = io_inValid_13 & _T_2003; // @[Switch.scala 30:36:@542.4]
  assign _T_2006 = io_inAddr_14 == 4'h6; // @[Switch.scala 30:53:@544.4]
  assign valid_6_14 = io_inValid_14 & _T_2006; // @[Switch.scala 30:36:@545.4]
  assign _T_2009 = io_inAddr_15 == 4'h6; // @[Switch.scala 30:53:@547.4]
  assign valid_6_15 = io_inValid_15 & _T_2009; // @[Switch.scala 30:36:@548.4]
  assign _T_2027 = valid_6_14 ? 4'he : 4'hf; // @[Mux.scala 31:69:@550.4]
  assign _T_2028 = valid_6_13 ? 4'hd : _T_2027; // @[Mux.scala 31:69:@551.4]
  assign _T_2029 = valid_6_12 ? 4'hc : _T_2028; // @[Mux.scala 31:69:@552.4]
  assign _T_2030 = valid_6_11 ? 4'hb : _T_2029; // @[Mux.scala 31:69:@553.4]
  assign _T_2031 = valid_6_10 ? 4'ha : _T_2030; // @[Mux.scala 31:69:@554.4]
  assign _T_2032 = valid_6_9 ? 4'h9 : _T_2031; // @[Mux.scala 31:69:@555.4]
  assign _T_2033 = valid_6_8 ? 4'h8 : _T_2032; // @[Mux.scala 31:69:@556.4]
  assign _T_2034 = valid_6_7 ? 4'h7 : _T_2033; // @[Mux.scala 31:69:@557.4]
  assign _T_2035 = valid_6_6 ? 4'h6 : _T_2034; // @[Mux.scala 31:69:@558.4]
  assign _T_2036 = valid_6_5 ? 4'h5 : _T_2035; // @[Mux.scala 31:69:@559.4]
  assign _T_2037 = valid_6_4 ? 4'h4 : _T_2036; // @[Mux.scala 31:69:@560.4]
  assign _T_2038 = valid_6_3 ? 4'h3 : _T_2037; // @[Mux.scala 31:69:@561.4]
  assign _T_2039 = valid_6_2 ? 4'h2 : _T_2038; // @[Mux.scala 31:69:@562.4]
  assign _T_2040 = valid_6_1 ? 4'h1 : _T_2039; // @[Mux.scala 31:69:@563.4]
  assign select_6 = valid_6_0 ? 4'h0 : _T_2040; // @[Mux.scala 31:69:@564.4]
  assign _GEN_97 = 4'h1 == select_6 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@566.4]
  assign _GEN_98 = 4'h2 == select_6 ? io_inData_2 : _GEN_97; // @[Switch.scala 33:19:@566.4]
  assign _GEN_99 = 4'h3 == select_6 ? io_inData_3 : _GEN_98; // @[Switch.scala 33:19:@566.4]
  assign _GEN_100 = 4'h4 == select_6 ? io_inData_4 : _GEN_99; // @[Switch.scala 33:19:@566.4]
  assign _GEN_101 = 4'h5 == select_6 ? io_inData_5 : _GEN_100; // @[Switch.scala 33:19:@566.4]
  assign _GEN_102 = 4'h6 == select_6 ? io_inData_6 : _GEN_101; // @[Switch.scala 33:19:@566.4]
  assign _GEN_103 = 4'h7 == select_6 ? io_inData_7 : _GEN_102; // @[Switch.scala 33:19:@566.4]
  assign _GEN_104 = 4'h8 == select_6 ? io_inData_8 : _GEN_103; // @[Switch.scala 33:19:@566.4]
  assign _GEN_105 = 4'h9 == select_6 ? io_inData_9 : _GEN_104; // @[Switch.scala 33:19:@566.4]
  assign _GEN_106 = 4'ha == select_6 ? io_inData_10 : _GEN_105; // @[Switch.scala 33:19:@566.4]
  assign _GEN_107 = 4'hb == select_6 ? io_inData_11 : _GEN_106; // @[Switch.scala 33:19:@566.4]
  assign _GEN_108 = 4'hc == select_6 ? io_inData_12 : _GEN_107; // @[Switch.scala 33:19:@566.4]
  assign _GEN_109 = 4'hd == select_6 ? io_inData_13 : _GEN_108; // @[Switch.scala 33:19:@566.4]
  assign _GEN_110 = 4'he == select_6 ? io_inData_14 : _GEN_109; // @[Switch.scala 33:19:@566.4]
  assign _T_2049 = {valid_6_7,valid_6_6,valid_6_5,valid_6_4,valid_6_3,valid_6_2,valid_6_1,valid_6_0}; // @[Switch.scala 34:32:@573.4]
  assign _T_2057 = {valid_6_15,valid_6_14,valid_6_13,valid_6_12,valid_6_11,valid_6_10,valid_6_9,valid_6_8,_T_2049}; // @[Switch.scala 34:32:@581.4]
  assign _T_2061 = io_inAddr_0 == 4'h7; // @[Switch.scala 30:53:@584.4]
  assign valid_7_0 = io_inValid_0 & _T_2061; // @[Switch.scala 30:36:@585.4]
  assign _T_2064 = io_inAddr_1 == 4'h7; // @[Switch.scala 30:53:@587.4]
  assign valid_7_1 = io_inValid_1 & _T_2064; // @[Switch.scala 30:36:@588.4]
  assign _T_2067 = io_inAddr_2 == 4'h7; // @[Switch.scala 30:53:@590.4]
  assign valid_7_2 = io_inValid_2 & _T_2067; // @[Switch.scala 30:36:@591.4]
  assign _T_2070 = io_inAddr_3 == 4'h7; // @[Switch.scala 30:53:@593.4]
  assign valid_7_3 = io_inValid_3 & _T_2070; // @[Switch.scala 30:36:@594.4]
  assign _T_2073 = io_inAddr_4 == 4'h7; // @[Switch.scala 30:53:@596.4]
  assign valid_7_4 = io_inValid_4 & _T_2073; // @[Switch.scala 30:36:@597.4]
  assign _T_2076 = io_inAddr_5 == 4'h7; // @[Switch.scala 30:53:@599.4]
  assign valid_7_5 = io_inValid_5 & _T_2076; // @[Switch.scala 30:36:@600.4]
  assign _T_2079 = io_inAddr_6 == 4'h7; // @[Switch.scala 30:53:@602.4]
  assign valid_7_6 = io_inValid_6 & _T_2079; // @[Switch.scala 30:36:@603.4]
  assign _T_2082 = io_inAddr_7 == 4'h7; // @[Switch.scala 30:53:@605.4]
  assign valid_7_7 = io_inValid_7 & _T_2082; // @[Switch.scala 30:36:@606.4]
  assign _T_2085 = io_inAddr_8 == 4'h7; // @[Switch.scala 30:53:@608.4]
  assign valid_7_8 = io_inValid_8 & _T_2085; // @[Switch.scala 30:36:@609.4]
  assign _T_2088 = io_inAddr_9 == 4'h7; // @[Switch.scala 30:53:@611.4]
  assign valid_7_9 = io_inValid_9 & _T_2088; // @[Switch.scala 30:36:@612.4]
  assign _T_2091 = io_inAddr_10 == 4'h7; // @[Switch.scala 30:53:@614.4]
  assign valid_7_10 = io_inValid_10 & _T_2091; // @[Switch.scala 30:36:@615.4]
  assign _T_2094 = io_inAddr_11 == 4'h7; // @[Switch.scala 30:53:@617.4]
  assign valid_7_11 = io_inValid_11 & _T_2094; // @[Switch.scala 30:36:@618.4]
  assign _T_2097 = io_inAddr_12 == 4'h7; // @[Switch.scala 30:53:@620.4]
  assign valid_7_12 = io_inValid_12 & _T_2097; // @[Switch.scala 30:36:@621.4]
  assign _T_2100 = io_inAddr_13 == 4'h7; // @[Switch.scala 30:53:@623.4]
  assign valid_7_13 = io_inValid_13 & _T_2100; // @[Switch.scala 30:36:@624.4]
  assign _T_2103 = io_inAddr_14 == 4'h7; // @[Switch.scala 30:53:@626.4]
  assign valid_7_14 = io_inValid_14 & _T_2103; // @[Switch.scala 30:36:@627.4]
  assign _T_2106 = io_inAddr_15 == 4'h7; // @[Switch.scala 30:53:@629.4]
  assign valid_7_15 = io_inValid_15 & _T_2106; // @[Switch.scala 30:36:@630.4]
  assign _T_2124 = valid_7_14 ? 4'he : 4'hf; // @[Mux.scala 31:69:@632.4]
  assign _T_2125 = valid_7_13 ? 4'hd : _T_2124; // @[Mux.scala 31:69:@633.4]
  assign _T_2126 = valid_7_12 ? 4'hc : _T_2125; // @[Mux.scala 31:69:@634.4]
  assign _T_2127 = valid_7_11 ? 4'hb : _T_2126; // @[Mux.scala 31:69:@635.4]
  assign _T_2128 = valid_7_10 ? 4'ha : _T_2127; // @[Mux.scala 31:69:@636.4]
  assign _T_2129 = valid_7_9 ? 4'h9 : _T_2128; // @[Mux.scala 31:69:@637.4]
  assign _T_2130 = valid_7_8 ? 4'h8 : _T_2129; // @[Mux.scala 31:69:@638.4]
  assign _T_2131 = valid_7_7 ? 4'h7 : _T_2130; // @[Mux.scala 31:69:@639.4]
  assign _T_2132 = valid_7_6 ? 4'h6 : _T_2131; // @[Mux.scala 31:69:@640.4]
  assign _T_2133 = valid_7_5 ? 4'h5 : _T_2132; // @[Mux.scala 31:69:@641.4]
  assign _T_2134 = valid_7_4 ? 4'h4 : _T_2133; // @[Mux.scala 31:69:@642.4]
  assign _T_2135 = valid_7_3 ? 4'h3 : _T_2134; // @[Mux.scala 31:69:@643.4]
  assign _T_2136 = valid_7_2 ? 4'h2 : _T_2135; // @[Mux.scala 31:69:@644.4]
  assign _T_2137 = valid_7_1 ? 4'h1 : _T_2136; // @[Mux.scala 31:69:@645.4]
  assign select_7 = valid_7_0 ? 4'h0 : _T_2137; // @[Mux.scala 31:69:@646.4]
  assign _GEN_113 = 4'h1 == select_7 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@648.4]
  assign _GEN_114 = 4'h2 == select_7 ? io_inData_2 : _GEN_113; // @[Switch.scala 33:19:@648.4]
  assign _GEN_115 = 4'h3 == select_7 ? io_inData_3 : _GEN_114; // @[Switch.scala 33:19:@648.4]
  assign _GEN_116 = 4'h4 == select_7 ? io_inData_4 : _GEN_115; // @[Switch.scala 33:19:@648.4]
  assign _GEN_117 = 4'h5 == select_7 ? io_inData_5 : _GEN_116; // @[Switch.scala 33:19:@648.4]
  assign _GEN_118 = 4'h6 == select_7 ? io_inData_6 : _GEN_117; // @[Switch.scala 33:19:@648.4]
  assign _GEN_119 = 4'h7 == select_7 ? io_inData_7 : _GEN_118; // @[Switch.scala 33:19:@648.4]
  assign _GEN_120 = 4'h8 == select_7 ? io_inData_8 : _GEN_119; // @[Switch.scala 33:19:@648.4]
  assign _GEN_121 = 4'h9 == select_7 ? io_inData_9 : _GEN_120; // @[Switch.scala 33:19:@648.4]
  assign _GEN_122 = 4'ha == select_7 ? io_inData_10 : _GEN_121; // @[Switch.scala 33:19:@648.4]
  assign _GEN_123 = 4'hb == select_7 ? io_inData_11 : _GEN_122; // @[Switch.scala 33:19:@648.4]
  assign _GEN_124 = 4'hc == select_7 ? io_inData_12 : _GEN_123; // @[Switch.scala 33:19:@648.4]
  assign _GEN_125 = 4'hd == select_7 ? io_inData_13 : _GEN_124; // @[Switch.scala 33:19:@648.4]
  assign _GEN_126 = 4'he == select_7 ? io_inData_14 : _GEN_125; // @[Switch.scala 33:19:@648.4]
  assign _T_2146 = {valid_7_7,valid_7_6,valid_7_5,valid_7_4,valid_7_3,valid_7_2,valid_7_1,valid_7_0}; // @[Switch.scala 34:32:@655.4]
  assign _T_2154 = {valid_7_15,valid_7_14,valid_7_13,valid_7_12,valid_7_11,valid_7_10,valid_7_9,valid_7_8,_T_2146}; // @[Switch.scala 34:32:@663.4]
  assign _T_2158 = io_inAddr_0 == 4'h8; // @[Switch.scala 30:53:@666.4]
  assign valid_8_0 = io_inValid_0 & _T_2158; // @[Switch.scala 30:36:@667.4]
  assign _T_2161 = io_inAddr_1 == 4'h8; // @[Switch.scala 30:53:@669.4]
  assign valid_8_1 = io_inValid_1 & _T_2161; // @[Switch.scala 30:36:@670.4]
  assign _T_2164 = io_inAddr_2 == 4'h8; // @[Switch.scala 30:53:@672.4]
  assign valid_8_2 = io_inValid_2 & _T_2164; // @[Switch.scala 30:36:@673.4]
  assign _T_2167 = io_inAddr_3 == 4'h8; // @[Switch.scala 30:53:@675.4]
  assign valid_8_3 = io_inValid_3 & _T_2167; // @[Switch.scala 30:36:@676.4]
  assign _T_2170 = io_inAddr_4 == 4'h8; // @[Switch.scala 30:53:@678.4]
  assign valid_8_4 = io_inValid_4 & _T_2170; // @[Switch.scala 30:36:@679.4]
  assign _T_2173 = io_inAddr_5 == 4'h8; // @[Switch.scala 30:53:@681.4]
  assign valid_8_5 = io_inValid_5 & _T_2173; // @[Switch.scala 30:36:@682.4]
  assign _T_2176 = io_inAddr_6 == 4'h8; // @[Switch.scala 30:53:@684.4]
  assign valid_8_6 = io_inValid_6 & _T_2176; // @[Switch.scala 30:36:@685.4]
  assign _T_2179 = io_inAddr_7 == 4'h8; // @[Switch.scala 30:53:@687.4]
  assign valid_8_7 = io_inValid_7 & _T_2179; // @[Switch.scala 30:36:@688.4]
  assign _T_2182 = io_inAddr_8 == 4'h8; // @[Switch.scala 30:53:@690.4]
  assign valid_8_8 = io_inValid_8 & _T_2182; // @[Switch.scala 30:36:@691.4]
  assign _T_2185 = io_inAddr_9 == 4'h8; // @[Switch.scala 30:53:@693.4]
  assign valid_8_9 = io_inValid_9 & _T_2185; // @[Switch.scala 30:36:@694.4]
  assign _T_2188 = io_inAddr_10 == 4'h8; // @[Switch.scala 30:53:@696.4]
  assign valid_8_10 = io_inValid_10 & _T_2188; // @[Switch.scala 30:36:@697.4]
  assign _T_2191 = io_inAddr_11 == 4'h8; // @[Switch.scala 30:53:@699.4]
  assign valid_8_11 = io_inValid_11 & _T_2191; // @[Switch.scala 30:36:@700.4]
  assign _T_2194 = io_inAddr_12 == 4'h8; // @[Switch.scala 30:53:@702.4]
  assign valid_8_12 = io_inValid_12 & _T_2194; // @[Switch.scala 30:36:@703.4]
  assign _T_2197 = io_inAddr_13 == 4'h8; // @[Switch.scala 30:53:@705.4]
  assign valid_8_13 = io_inValid_13 & _T_2197; // @[Switch.scala 30:36:@706.4]
  assign _T_2200 = io_inAddr_14 == 4'h8; // @[Switch.scala 30:53:@708.4]
  assign valid_8_14 = io_inValid_14 & _T_2200; // @[Switch.scala 30:36:@709.4]
  assign _T_2203 = io_inAddr_15 == 4'h8; // @[Switch.scala 30:53:@711.4]
  assign valid_8_15 = io_inValid_15 & _T_2203; // @[Switch.scala 30:36:@712.4]
  assign _T_2221 = valid_8_14 ? 4'he : 4'hf; // @[Mux.scala 31:69:@714.4]
  assign _T_2222 = valid_8_13 ? 4'hd : _T_2221; // @[Mux.scala 31:69:@715.4]
  assign _T_2223 = valid_8_12 ? 4'hc : _T_2222; // @[Mux.scala 31:69:@716.4]
  assign _T_2224 = valid_8_11 ? 4'hb : _T_2223; // @[Mux.scala 31:69:@717.4]
  assign _T_2225 = valid_8_10 ? 4'ha : _T_2224; // @[Mux.scala 31:69:@718.4]
  assign _T_2226 = valid_8_9 ? 4'h9 : _T_2225; // @[Mux.scala 31:69:@719.4]
  assign _T_2227 = valid_8_8 ? 4'h8 : _T_2226; // @[Mux.scala 31:69:@720.4]
  assign _T_2228 = valid_8_7 ? 4'h7 : _T_2227; // @[Mux.scala 31:69:@721.4]
  assign _T_2229 = valid_8_6 ? 4'h6 : _T_2228; // @[Mux.scala 31:69:@722.4]
  assign _T_2230 = valid_8_5 ? 4'h5 : _T_2229; // @[Mux.scala 31:69:@723.4]
  assign _T_2231 = valid_8_4 ? 4'h4 : _T_2230; // @[Mux.scala 31:69:@724.4]
  assign _T_2232 = valid_8_3 ? 4'h3 : _T_2231; // @[Mux.scala 31:69:@725.4]
  assign _T_2233 = valid_8_2 ? 4'h2 : _T_2232; // @[Mux.scala 31:69:@726.4]
  assign _T_2234 = valid_8_1 ? 4'h1 : _T_2233; // @[Mux.scala 31:69:@727.4]
  assign select_8 = valid_8_0 ? 4'h0 : _T_2234; // @[Mux.scala 31:69:@728.4]
  assign _GEN_129 = 4'h1 == select_8 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@730.4]
  assign _GEN_130 = 4'h2 == select_8 ? io_inData_2 : _GEN_129; // @[Switch.scala 33:19:@730.4]
  assign _GEN_131 = 4'h3 == select_8 ? io_inData_3 : _GEN_130; // @[Switch.scala 33:19:@730.4]
  assign _GEN_132 = 4'h4 == select_8 ? io_inData_4 : _GEN_131; // @[Switch.scala 33:19:@730.4]
  assign _GEN_133 = 4'h5 == select_8 ? io_inData_5 : _GEN_132; // @[Switch.scala 33:19:@730.4]
  assign _GEN_134 = 4'h6 == select_8 ? io_inData_6 : _GEN_133; // @[Switch.scala 33:19:@730.4]
  assign _GEN_135 = 4'h7 == select_8 ? io_inData_7 : _GEN_134; // @[Switch.scala 33:19:@730.4]
  assign _GEN_136 = 4'h8 == select_8 ? io_inData_8 : _GEN_135; // @[Switch.scala 33:19:@730.4]
  assign _GEN_137 = 4'h9 == select_8 ? io_inData_9 : _GEN_136; // @[Switch.scala 33:19:@730.4]
  assign _GEN_138 = 4'ha == select_8 ? io_inData_10 : _GEN_137; // @[Switch.scala 33:19:@730.4]
  assign _GEN_139 = 4'hb == select_8 ? io_inData_11 : _GEN_138; // @[Switch.scala 33:19:@730.4]
  assign _GEN_140 = 4'hc == select_8 ? io_inData_12 : _GEN_139; // @[Switch.scala 33:19:@730.4]
  assign _GEN_141 = 4'hd == select_8 ? io_inData_13 : _GEN_140; // @[Switch.scala 33:19:@730.4]
  assign _GEN_142 = 4'he == select_8 ? io_inData_14 : _GEN_141; // @[Switch.scala 33:19:@730.4]
  assign _T_2243 = {valid_8_7,valid_8_6,valid_8_5,valid_8_4,valid_8_3,valid_8_2,valid_8_1,valid_8_0}; // @[Switch.scala 34:32:@737.4]
  assign _T_2251 = {valid_8_15,valid_8_14,valid_8_13,valid_8_12,valid_8_11,valid_8_10,valid_8_9,valid_8_8,_T_2243}; // @[Switch.scala 34:32:@745.4]
  assign _T_2255 = io_inAddr_0 == 4'h9; // @[Switch.scala 30:53:@748.4]
  assign valid_9_0 = io_inValid_0 & _T_2255; // @[Switch.scala 30:36:@749.4]
  assign _T_2258 = io_inAddr_1 == 4'h9; // @[Switch.scala 30:53:@751.4]
  assign valid_9_1 = io_inValid_1 & _T_2258; // @[Switch.scala 30:36:@752.4]
  assign _T_2261 = io_inAddr_2 == 4'h9; // @[Switch.scala 30:53:@754.4]
  assign valid_9_2 = io_inValid_2 & _T_2261; // @[Switch.scala 30:36:@755.4]
  assign _T_2264 = io_inAddr_3 == 4'h9; // @[Switch.scala 30:53:@757.4]
  assign valid_9_3 = io_inValid_3 & _T_2264; // @[Switch.scala 30:36:@758.4]
  assign _T_2267 = io_inAddr_4 == 4'h9; // @[Switch.scala 30:53:@760.4]
  assign valid_9_4 = io_inValid_4 & _T_2267; // @[Switch.scala 30:36:@761.4]
  assign _T_2270 = io_inAddr_5 == 4'h9; // @[Switch.scala 30:53:@763.4]
  assign valid_9_5 = io_inValid_5 & _T_2270; // @[Switch.scala 30:36:@764.4]
  assign _T_2273 = io_inAddr_6 == 4'h9; // @[Switch.scala 30:53:@766.4]
  assign valid_9_6 = io_inValid_6 & _T_2273; // @[Switch.scala 30:36:@767.4]
  assign _T_2276 = io_inAddr_7 == 4'h9; // @[Switch.scala 30:53:@769.4]
  assign valid_9_7 = io_inValid_7 & _T_2276; // @[Switch.scala 30:36:@770.4]
  assign _T_2279 = io_inAddr_8 == 4'h9; // @[Switch.scala 30:53:@772.4]
  assign valid_9_8 = io_inValid_8 & _T_2279; // @[Switch.scala 30:36:@773.4]
  assign _T_2282 = io_inAddr_9 == 4'h9; // @[Switch.scala 30:53:@775.4]
  assign valid_9_9 = io_inValid_9 & _T_2282; // @[Switch.scala 30:36:@776.4]
  assign _T_2285 = io_inAddr_10 == 4'h9; // @[Switch.scala 30:53:@778.4]
  assign valid_9_10 = io_inValid_10 & _T_2285; // @[Switch.scala 30:36:@779.4]
  assign _T_2288 = io_inAddr_11 == 4'h9; // @[Switch.scala 30:53:@781.4]
  assign valid_9_11 = io_inValid_11 & _T_2288; // @[Switch.scala 30:36:@782.4]
  assign _T_2291 = io_inAddr_12 == 4'h9; // @[Switch.scala 30:53:@784.4]
  assign valid_9_12 = io_inValid_12 & _T_2291; // @[Switch.scala 30:36:@785.4]
  assign _T_2294 = io_inAddr_13 == 4'h9; // @[Switch.scala 30:53:@787.4]
  assign valid_9_13 = io_inValid_13 & _T_2294; // @[Switch.scala 30:36:@788.4]
  assign _T_2297 = io_inAddr_14 == 4'h9; // @[Switch.scala 30:53:@790.4]
  assign valid_9_14 = io_inValid_14 & _T_2297; // @[Switch.scala 30:36:@791.4]
  assign _T_2300 = io_inAddr_15 == 4'h9; // @[Switch.scala 30:53:@793.4]
  assign valid_9_15 = io_inValid_15 & _T_2300; // @[Switch.scala 30:36:@794.4]
  assign _T_2318 = valid_9_14 ? 4'he : 4'hf; // @[Mux.scala 31:69:@796.4]
  assign _T_2319 = valid_9_13 ? 4'hd : _T_2318; // @[Mux.scala 31:69:@797.4]
  assign _T_2320 = valid_9_12 ? 4'hc : _T_2319; // @[Mux.scala 31:69:@798.4]
  assign _T_2321 = valid_9_11 ? 4'hb : _T_2320; // @[Mux.scala 31:69:@799.4]
  assign _T_2322 = valid_9_10 ? 4'ha : _T_2321; // @[Mux.scala 31:69:@800.4]
  assign _T_2323 = valid_9_9 ? 4'h9 : _T_2322; // @[Mux.scala 31:69:@801.4]
  assign _T_2324 = valid_9_8 ? 4'h8 : _T_2323; // @[Mux.scala 31:69:@802.4]
  assign _T_2325 = valid_9_7 ? 4'h7 : _T_2324; // @[Mux.scala 31:69:@803.4]
  assign _T_2326 = valid_9_6 ? 4'h6 : _T_2325; // @[Mux.scala 31:69:@804.4]
  assign _T_2327 = valid_9_5 ? 4'h5 : _T_2326; // @[Mux.scala 31:69:@805.4]
  assign _T_2328 = valid_9_4 ? 4'h4 : _T_2327; // @[Mux.scala 31:69:@806.4]
  assign _T_2329 = valid_9_3 ? 4'h3 : _T_2328; // @[Mux.scala 31:69:@807.4]
  assign _T_2330 = valid_9_2 ? 4'h2 : _T_2329; // @[Mux.scala 31:69:@808.4]
  assign _T_2331 = valid_9_1 ? 4'h1 : _T_2330; // @[Mux.scala 31:69:@809.4]
  assign select_9 = valid_9_0 ? 4'h0 : _T_2331; // @[Mux.scala 31:69:@810.4]
  assign _GEN_145 = 4'h1 == select_9 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@812.4]
  assign _GEN_146 = 4'h2 == select_9 ? io_inData_2 : _GEN_145; // @[Switch.scala 33:19:@812.4]
  assign _GEN_147 = 4'h3 == select_9 ? io_inData_3 : _GEN_146; // @[Switch.scala 33:19:@812.4]
  assign _GEN_148 = 4'h4 == select_9 ? io_inData_4 : _GEN_147; // @[Switch.scala 33:19:@812.4]
  assign _GEN_149 = 4'h5 == select_9 ? io_inData_5 : _GEN_148; // @[Switch.scala 33:19:@812.4]
  assign _GEN_150 = 4'h6 == select_9 ? io_inData_6 : _GEN_149; // @[Switch.scala 33:19:@812.4]
  assign _GEN_151 = 4'h7 == select_9 ? io_inData_7 : _GEN_150; // @[Switch.scala 33:19:@812.4]
  assign _GEN_152 = 4'h8 == select_9 ? io_inData_8 : _GEN_151; // @[Switch.scala 33:19:@812.4]
  assign _GEN_153 = 4'h9 == select_9 ? io_inData_9 : _GEN_152; // @[Switch.scala 33:19:@812.4]
  assign _GEN_154 = 4'ha == select_9 ? io_inData_10 : _GEN_153; // @[Switch.scala 33:19:@812.4]
  assign _GEN_155 = 4'hb == select_9 ? io_inData_11 : _GEN_154; // @[Switch.scala 33:19:@812.4]
  assign _GEN_156 = 4'hc == select_9 ? io_inData_12 : _GEN_155; // @[Switch.scala 33:19:@812.4]
  assign _GEN_157 = 4'hd == select_9 ? io_inData_13 : _GEN_156; // @[Switch.scala 33:19:@812.4]
  assign _GEN_158 = 4'he == select_9 ? io_inData_14 : _GEN_157; // @[Switch.scala 33:19:@812.4]
  assign _T_2340 = {valid_9_7,valid_9_6,valid_9_5,valid_9_4,valid_9_3,valid_9_2,valid_9_1,valid_9_0}; // @[Switch.scala 34:32:@819.4]
  assign _T_2348 = {valid_9_15,valid_9_14,valid_9_13,valid_9_12,valid_9_11,valid_9_10,valid_9_9,valid_9_8,_T_2340}; // @[Switch.scala 34:32:@827.4]
  assign _T_2352 = io_inAddr_0 == 4'ha; // @[Switch.scala 30:53:@830.4]
  assign valid_10_0 = io_inValid_0 & _T_2352; // @[Switch.scala 30:36:@831.4]
  assign _T_2355 = io_inAddr_1 == 4'ha; // @[Switch.scala 30:53:@833.4]
  assign valid_10_1 = io_inValid_1 & _T_2355; // @[Switch.scala 30:36:@834.4]
  assign _T_2358 = io_inAddr_2 == 4'ha; // @[Switch.scala 30:53:@836.4]
  assign valid_10_2 = io_inValid_2 & _T_2358; // @[Switch.scala 30:36:@837.4]
  assign _T_2361 = io_inAddr_3 == 4'ha; // @[Switch.scala 30:53:@839.4]
  assign valid_10_3 = io_inValid_3 & _T_2361; // @[Switch.scala 30:36:@840.4]
  assign _T_2364 = io_inAddr_4 == 4'ha; // @[Switch.scala 30:53:@842.4]
  assign valid_10_4 = io_inValid_4 & _T_2364; // @[Switch.scala 30:36:@843.4]
  assign _T_2367 = io_inAddr_5 == 4'ha; // @[Switch.scala 30:53:@845.4]
  assign valid_10_5 = io_inValid_5 & _T_2367; // @[Switch.scala 30:36:@846.4]
  assign _T_2370 = io_inAddr_6 == 4'ha; // @[Switch.scala 30:53:@848.4]
  assign valid_10_6 = io_inValid_6 & _T_2370; // @[Switch.scala 30:36:@849.4]
  assign _T_2373 = io_inAddr_7 == 4'ha; // @[Switch.scala 30:53:@851.4]
  assign valid_10_7 = io_inValid_7 & _T_2373; // @[Switch.scala 30:36:@852.4]
  assign _T_2376 = io_inAddr_8 == 4'ha; // @[Switch.scala 30:53:@854.4]
  assign valid_10_8 = io_inValid_8 & _T_2376; // @[Switch.scala 30:36:@855.4]
  assign _T_2379 = io_inAddr_9 == 4'ha; // @[Switch.scala 30:53:@857.4]
  assign valid_10_9 = io_inValid_9 & _T_2379; // @[Switch.scala 30:36:@858.4]
  assign _T_2382 = io_inAddr_10 == 4'ha; // @[Switch.scala 30:53:@860.4]
  assign valid_10_10 = io_inValid_10 & _T_2382; // @[Switch.scala 30:36:@861.4]
  assign _T_2385 = io_inAddr_11 == 4'ha; // @[Switch.scala 30:53:@863.4]
  assign valid_10_11 = io_inValid_11 & _T_2385; // @[Switch.scala 30:36:@864.4]
  assign _T_2388 = io_inAddr_12 == 4'ha; // @[Switch.scala 30:53:@866.4]
  assign valid_10_12 = io_inValid_12 & _T_2388; // @[Switch.scala 30:36:@867.4]
  assign _T_2391 = io_inAddr_13 == 4'ha; // @[Switch.scala 30:53:@869.4]
  assign valid_10_13 = io_inValid_13 & _T_2391; // @[Switch.scala 30:36:@870.4]
  assign _T_2394 = io_inAddr_14 == 4'ha; // @[Switch.scala 30:53:@872.4]
  assign valid_10_14 = io_inValid_14 & _T_2394; // @[Switch.scala 30:36:@873.4]
  assign _T_2397 = io_inAddr_15 == 4'ha; // @[Switch.scala 30:53:@875.4]
  assign valid_10_15 = io_inValid_15 & _T_2397; // @[Switch.scala 30:36:@876.4]
  assign _T_2415 = valid_10_14 ? 4'he : 4'hf; // @[Mux.scala 31:69:@878.4]
  assign _T_2416 = valid_10_13 ? 4'hd : _T_2415; // @[Mux.scala 31:69:@879.4]
  assign _T_2417 = valid_10_12 ? 4'hc : _T_2416; // @[Mux.scala 31:69:@880.4]
  assign _T_2418 = valid_10_11 ? 4'hb : _T_2417; // @[Mux.scala 31:69:@881.4]
  assign _T_2419 = valid_10_10 ? 4'ha : _T_2418; // @[Mux.scala 31:69:@882.4]
  assign _T_2420 = valid_10_9 ? 4'h9 : _T_2419; // @[Mux.scala 31:69:@883.4]
  assign _T_2421 = valid_10_8 ? 4'h8 : _T_2420; // @[Mux.scala 31:69:@884.4]
  assign _T_2422 = valid_10_7 ? 4'h7 : _T_2421; // @[Mux.scala 31:69:@885.4]
  assign _T_2423 = valid_10_6 ? 4'h6 : _T_2422; // @[Mux.scala 31:69:@886.4]
  assign _T_2424 = valid_10_5 ? 4'h5 : _T_2423; // @[Mux.scala 31:69:@887.4]
  assign _T_2425 = valid_10_4 ? 4'h4 : _T_2424; // @[Mux.scala 31:69:@888.4]
  assign _T_2426 = valid_10_3 ? 4'h3 : _T_2425; // @[Mux.scala 31:69:@889.4]
  assign _T_2427 = valid_10_2 ? 4'h2 : _T_2426; // @[Mux.scala 31:69:@890.4]
  assign _T_2428 = valid_10_1 ? 4'h1 : _T_2427; // @[Mux.scala 31:69:@891.4]
  assign select_10 = valid_10_0 ? 4'h0 : _T_2428; // @[Mux.scala 31:69:@892.4]
  assign _GEN_161 = 4'h1 == select_10 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@894.4]
  assign _GEN_162 = 4'h2 == select_10 ? io_inData_2 : _GEN_161; // @[Switch.scala 33:19:@894.4]
  assign _GEN_163 = 4'h3 == select_10 ? io_inData_3 : _GEN_162; // @[Switch.scala 33:19:@894.4]
  assign _GEN_164 = 4'h4 == select_10 ? io_inData_4 : _GEN_163; // @[Switch.scala 33:19:@894.4]
  assign _GEN_165 = 4'h5 == select_10 ? io_inData_5 : _GEN_164; // @[Switch.scala 33:19:@894.4]
  assign _GEN_166 = 4'h6 == select_10 ? io_inData_6 : _GEN_165; // @[Switch.scala 33:19:@894.4]
  assign _GEN_167 = 4'h7 == select_10 ? io_inData_7 : _GEN_166; // @[Switch.scala 33:19:@894.4]
  assign _GEN_168 = 4'h8 == select_10 ? io_inData_8 : _GEN_167; // @[Switch.scala 33:19:@894.4]
  assign _GEN_169 = 4'h9 == select_10 ? io_inData_9 : _GEN_168; // @[Switch.scala 33:19:@894.4]
  assign _GEN_170 = 4'ha == select_10 ? io_inData_10 : _GEN_169; // @[Switch.scala 33:19:@894.4]
  assign _GEN_171 = 4'hb == select_10 ? io_inData_11 : _GEN_170; // @[Switch.scala 33:19:@894.4]
  assign _GEN_172 = 4'hc == select_10 ? io_inData_12 : _GEN_171; // @[Switch.scala 33:19:@894.4]
  assign _GEN_173 = 4'hd == select_10 ? io_inData_13 : _GEN_172; // @[Switch.scala 33:19:@894.4]
  assign _GEN_174 = 4'he == select_10 ? io_inData_14 : _GEN_173; // @[Switch.scala 33:19:@894.4]
  assign _T_2437 = {valid_10_7,valid_10_6,valid_10_5,valid_10_4,valid_10_3,valid_10_2,valid_10_1,valid_10_0}; // @[Switch.scala 34:32:@901.4]
  assign _T_2445 = {valid_10_15,valid_10_14,valid_10_13,valid_10_12,valid_10_11,valid_10_10,valid_10_9,valid_10_8,_T_2437}; // @[Switch.scala 34:32:@909.4]
  assign _T_2449 = io_inAddr_0 == 4'hb; // @[Switch.scala 30:53:@912.4]
  assign valid_11_0 = io_inValid_0 & _T_2449; // @[Switch.scala 30:36:@913.4]
  assign _T_2452 = io_inAddr_1 == 4'hb; // @[Switch.scala 30:53:@915.4]
  assign valid_11_1 = io_inValid_1 & _T_2452; // @[Switch.scala 30:36:@916.4]
  assign _T_2455 = io_inAddr_2 == 4'hb; // @[Switch.scala 30:53:@918.4]
  assign valid_11_2 = io_inValid_2 & _T_2455; // @[Switch.scala 30:36:@919.4]
  assign _T_2458 = io_inAddr_3 == 4'hb; // @[Switch.scala 30:53:@921.4]
  assign valid_11_3 = io_inValid_3 & _T_2458; // @[Switch.scala 30:36:@922.4]
  assign _T_2461 = io_inAddr_4 == 4'hb; // @[Switch.scala 30:53:@924.4]
  assign valid_11_4 = io_inValid_4 & _T_2461; // @[Switch.scala 30:36:@925.4]
  assign _T_2464 = io_inAddr_5 == 4'hb; // @[Switch.scala 30:53:@927.4]
  assign valid_11_5 = io_inValid_5 & _T_2464; // @[Switch.scala 30:36:@928.4]
  assign _T_2467 = io_inAddr_6 == 4'hb; // @[Switch.scala 30:53:@930.4]
  assign valid_11_6 = io_inValid_6 & _T_2467; // @[Switch.scala 30:36:@931.4]
  assign _T_2470 = io_inAddr_7 == 4'hb; // @[Switch.scala 30:53:@933.4]
  assign valid_11_7 = io_inValid_7 & _T_2470; // @[Switch.scala 30:36:@934.4]
  assign _T_2473 = io_inAddr_8 == 4'hb; // @[Switch.scala 30:53:@936.4]
  assign valid_11_8 = io_inValid_8 & _T_2473; // @[Switch.scala 30:36:@937.4]
  assign _T_2476 = io_inAddr_9 == 4'hb; // @[Switch.scala 30:53:@939.4]
  assign valid_11_9 = io_inValid_9 & _T_2476; // @[Switch.scala 30:36:@940.4]
  assign _T_2479 = io_inAddr_10 == 4'hb; // @[Switch.scala 30:53:@942.4]
  assign valid_11_10 = io_inValid_10 & _T_2479; // @[Switch.scala 30:36:@943.4]
  assign _T_2482 = io_inAddr_11 == 4'hb; // @[Switch.scala 30:53:@945.4]
  assign valid_11_11 = io_inValid_11 & _T_2482; // @[Switch.scala 30:36:@946.4]
  assign _T_2485 = io_inAddr_12 == 4'hb; // @[Switch.scala 30:53:@948.4]
  assign valid_11_12 = io_inValid_12 & _T_2485; // @[Switch.scala 30:36:@949.4]
  assign _T_2488 = io_inAddr_13 == 4'hb; // @[Switch.scala 30:53:@951.4]
  assign valid_11_13 = io_inValid_13 & _T_2488; // @[Switch.scala 30:36:@952.4]
  assign _T_2491 = io_inAddr_14 == 4'hb; // @[Switch.scala 30:53:@954.4]
  assign valid_11_14 = io_inValid_14 & _T_2491; // @[Switch.scala 30:36:@955.4]
  assign _T_2494 = io_inAddr_15 == 4'hb; // @[Switch.scala 30:53:@957.4]
  assign valid_11_15 = io_inValid_15 & _T_2494; // @[Switch.scala 30:36:@958.4]
  assign _T_2512 = valid_11_14 ? 4'he : 4'hf; // @[Mux.scala 31:69:@960.4]
  assign _T_2513 = valid_11_13 ? 4'hd : _T_2512; // @[Mux.scala 31:69:@961.4]
  assign _T_2514 = valid_11_12 ? 4'hc : _T_2513; // @[Mux.scala 31:69:@962.4]
  assign _T_2515 = valid_11_11 ? 4'hb : _T_2514; // @[Mux.scala 31:69:@963.4]
  assign _T_2516 = valid_11_10 ? 4'ha : _T_2515; // @[Mux.scala 31:69:@964.4]
  assign _T_2517 = valid_11_9 ? 4'h9 : _T_2516; // @[Mux.scala 31:69:@965.4]
  assign _T_2518 = valid_11_8 ? 4'h8 : _T_2517; // @[Mux.scala 31:69:@966.4]
  assign _T_2519 = valid_11_7 ? 4'h7 : _T_2518; // @[Mux.scala 31:69:@967.4]
  assign _T_2520 = valid_11_6 ? 4'h6 : _T_2519; // @[Mux.scala 31:69:@968.4]
  assign _T_2521 = valid_11_5 ? 4'h5 : _T_2520; // @[Mux.scala 31:69:@969.4]
  assign _T_2522 = valid_11_4 ? 4'h4 : _T_2521; // @[Mux.scala 31:69:@970.4]
  assign _T_2523 = valid_11_3 ? 4'h3 : _T_2522; // @[Mux.scala 31:69:@971.4]
  assign _T_2524 = valid_11_2 ? 4'h2 : _T_2523; // @[Mux.scala 31:69:@972.4]
  assign _T_2525 = valid_11_1 ? 4'h1 : _T_2524; // @[Mux.scala 31:69:@973.4]
  assign select_11 = valid_11_0 ? 4'h0 : _T_2525; // @[Mux.scala 31:69:@974.4]
  assign _GEN_177 = 4'h1 == select_11 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@976.4]
  assign _GEN_178 = 4'h2 == select_11 ? io_inData_2 : _GEN_177; // @[Switch.scala 33:19:@976.4]
  assign _GEN_179 = 4'h3 == select_11 ? io_inData_3 : _GEN_178; // @[Switch.scala 33:19:@976.4]
  assign _GEN_180 = 4'h4 == select_11 ? io_inData_4 : _GEN_179; // @[Switch.scala 33:19:@976.4]
  assign _GEN_181 = 4'h5 == select_11 ? io_inData_5 : _GEN_180; // @[Switch.scala 33:19:@976.4]
  assign _GEN_182 = 4'h6 == select_11 ? io_inData_6 : _GEN_181; // @[Switch.scala 33:19:@976.4]
  assign _GEN_183 = 4'h7 == select_11 ? io_inData_7 : _GEN_182; // @[Switch.scala 33:19:@976.4]
  assign _GEN_184 = 4'h8 == select_11 ? io_inData_8 : _GEN_183; // @[Switch.scala 33:19:@976.4]
  assign _GEN_185 = 4'h9 == select_11 ? io_inData_9 : _GEN_184; // @[Switch.scala 33:19:@976.4]
  assign _GEN_186 = 4'ha == select_11 ? io_inData_10 : _GEN_185; // @[Switch.scala 33:19:@976.4]
  assign _GEN_187 = 4'hb == select_11 ? io_inData_11 : _GEN_186; // @[Switch.scala 33:19:@976.4]
  assign _GEN_188 = 4'hc == select_11 ? io_inData_12 : _GEN_187; // @[Switch.scala 33:19:@976.4]
  assign _GEN_189 = 4'hd == select_11 ? io_inData_13 : _GEN_188; // @[Switch.scala 33:19:@976.4]
  assign _GEN_190 = 4'he == select_11 ? io_inData_14 : _GEN_189; // @[Switch.scala 33:19:@976.4]
  assign _T_2534 = {valid_11_7,valid_11_6,valid_11_5,valid_11_4,valid_11_3,valid_11_2,valid_11_1,valid_11_0}; // @[Switch.scala 34:32:@983.4]
  assign _T_2542 = {valid_11_15,valid_11_14,valid_11_13,valid_11_12,valid_11_11,valid_11_10,valid_11_9,valid_11_8,_T_2534}; // @[Switch.scala 34:32:@991.4]
  assign _T_2546 = io_inAddr_0 == 4'hc; // @[Switch.scala 30:53:@994.4]
  assign valid_12_0 = io_inValid_0 & _T_2546; // @[Switch.scala 30:36:@995.4]
  assign _T_2549 = io_inAddr_1 == 4'hc; // @[Switch.scala 30:53:@997.4]
  assign valid_12_1 = io_inValid_1 & _T_2549; // @[Switch.scala 30:36:@998.4]
  assign _T_2552 = io_inAddr_2 == 4'hc; // @[Switch.scala 30:53:@1000.4]
  assign valid_12_2 = io_inValid_2 & _T_2552; // @[Switch.scala 30:36:@1001.4]
  assign _T_2555 = io_inAddr_3 == 4'hc; // @[Switch.scala 30:53:@1003.4]
  assign valid_12_3 = io_inValid_3 & _T_2555; // @[Switch.scala 30:36:@1004.4]
  assign _T_2558 = io_inAddr_4 == 4'hc; // @[Switch.scala 30:53:@1006.4]
  assign valid_12_4 = io_inValid_4 & _T_2558; // @[Switch.scala 30:36:@1007.4]
  assign _T_2561 = io_inAddr_5 == 4'hc; // @[Switch.scala 30:53:@1009.4]
  assign valid_12_5 = io_inValid_5 & _T_2561; // @[Switch.scala 30:36:@1010.4]
  assign _T_2564 = io_inAddr_6 == 4'hc; // @[Switch.scala 30:53:@1012.4]
  assign valid_12_6 = io_inValid_6 & _T_2564; // @[Switch.scala 30:36:@1013.4]
  assign _T_2567 = io_inAddr_7 == 4'hc; // @[Switch.scala 30:53:@1015.4]
  assign valid_12_7 = io_inValid_7 & _T_2567; // @[Switch.scala 30:36:@1016.4]
  assign _T_2570 = io_inAddr_8 == 4'hc; // @[Switch.scala 30:53:@1018.4]
  assign valid_12_8 = io_inValid_8 & _T_2570; // @[Switch.scala 30:36:@1019.4]
  assign _T_2573 = io_inAddr_9 == 4'hc; // @[Switch.scala 30:53:@1021.4]
  assign valid_12_9 = io_inValid_9 & _T_2573; // @[Switch.scala 30:36:@1022.4]
  assign _T_2576 = io_inAddr_10 == 4'hc; // @[Switch.scala 30:53:@1024.4]
  assign valid_12_10 = io_inValid_10 & _T_2576; // @[Switch.scala 30:36:@1025.4]
  assign _T_2579 = io_inAddr_11 == 4'hc; // @[Switch.scala 30:53:@1027.4]
  assign valid_12_11 = io_inValid_11 & _T_2579; // @[Switch.scala 30:36:@1028.4]
  assign _T_2582 = io_inAddr_12 == 4'hc; // @[Switch.scala 30:53:@1030.4]
  assign valid_12_12 = io_inValid_12 & _T_2582; // @[Switch.scala 30:36:@1031.4]
  assign _T_2585 = io_inAddr_13 == 4'hc; // @[Switch.scala 30:53:@1033.4]
  assign valid_12_13 = io_inValid_13 & _T_2585; // @[Switch.scala 30:36:@1034.4]
  assign _T_2588 = io_inAddr_14 == 4'hc; // @[Switch.scala 30:53:@1036.4]
  assign valid_12_14 = io_inValid_14 & _T_2588; // @[Switch.scala 30:36:@1037.4]
  assign _T_2591 = io_inAddr_15 == 4'hc; // @[Switch.scala 30:53:@1039.4]
  assign valid_12_15 = io_inValid_15 & _T_2591; // @[Switch.scala 30:36:@1040.4]
  assign _T_2609 = valid_12_14 ? 4'he : 4'hf; // @[Mux.scala 31:69:@1042.4]
  assign _T_2610 = valid_12_13 ? 4'hd : _T_2609; // @[Mux.scala 31:69:@1043.4]
  assign _T_2611 = valid_12_12 ? 4'hc : _T_2610; // @[Mux.scala 31:69:@1044.4]
  assign _T_2612 = valid_12_11 ? 4'hb : _T_2611; // @[Mux.scala 31:69:@1045.4]
  assign _T_2613 = valid_12_10 ? 4'ha : _T_2612; // @[Mux.scala 31:69:@1046.4]
  assign _T_2614 = valid_12_9 ? 4'h9 : _T_2613; // @[Mux.scala 31:69:@1047.4]
  assign _T_2615 = valid_12_8 ? 4'h8 : _T_2614; // @[Mux.scala 31:69:@1048.4]
  assign _T_2616 = valid_12_7 ? 4'h7 : _T_2615; // @[Mux.scala 31:69:@1049.4]
  assign _T_2617 = valid_12_6 ? 4'h6 : _T_2616; // @[Mux.scala 31:69:@1050.4]
  assign _T_2618 = valid_12_5 ? 4'h5 : _T_2617; // @[Mux.scala 31:69:@1051.4]
  assign _T_2619 = valid_12_4 ? 4'h4 : _T_2618; // @[Mux.scala 31:69:@1052.4]
  assign _T_2620 = valid_12_3 ? 4'h3 : _T_2619; // @[Mux.scala 31:69:@1053.4]
  assign _T_2621 = valid_12_2 ? 4'h2 : _T_2620; // @[Mux.scala 31:69:@1054.4]
  assign _T_2622 = valid_12_1 ? 4'h1 : _T_2621; // @[Mux.scala 31:69:@1055.4]
  assign select_12 = valid_12_0 ? 4'h0 : _T_2622; // @[Mux.scala 31:69:@1056.4]
  assign _GEN_193 = 4'h1 == select_12 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@1058.4]
  assign _GEN_194 = 4'h2 == select_12 ? io_inData_2 : _GEN_193; // @[Switch.scala 33:19:@1058.4]
  assign _GEN_195 = 4'h3 == select_12 ? io_inData_3 : _GEN_194; // @[Switch.scala 33:19:@1058.4]
  assign _GEN_196 = 4'h4 == select_12 ? io_inData_4 : _GEN_195; // @[Switch.scala 33:19:@1058.4]
  assign _GEN_197 = 4'h5 == select_12 ? io_inData_5 : _GEN_196; // @[Switch.scala 33:19:@1058.4]
  assign _GEN_198 = 4'h6 == select_12 ? io_inData_6 : _GEN_197; // @[Switch.scala 33:19:@1058.4]
  assign _GEN_199 = 4'h7 == select_12 ? io_inData_7 : _GEN_198; // @[Switch.scala 33:19:@1058.4]
  assign _GEN_200 = 4'h8 == select_12 ? io_inData_8 : _GEN_199; // @[Switch.scala 33:19:@1058.4]
  assign _GEN_201 = 4'h9 == select_12 ? io_inData_9 : _GEN_200; // @[Switch.scala 33:19:@1058.4]
  assign _GEN_202 = 4'ha == select_12 ? io_inData_10 : _GEN_201; // @[Switch.scala 33:19:@1058.4]
  assign _GEN_203 = 4'hb == select_12 ? io_inData_11 : _GEN_202; // @[Switch.scala 33:19:@1058.4]
  assign _GEN_204 = 4'hc == select_12 ? io_inData_12 : _GEN_203; // @[Switch.scala 33:19:@1058.4]
  assign _GEN_205 = 4'hd == select_12 ? io_inData_13 : _GEN_204; // @[Switch.scala 33:19:@1058.4]
  assign _GEN_206 = 4'he == select_12 ? io_inData_14 : _GEN_205; // @[Switch.scala 33:19:@1058.4]
  assign _T_2631 = {valid_12_7,valid_12_6,valid_12_5,valid_12_4,valid_12_3,valid_12_2,valid_12_1,valid_12_0}; // @[Switch.scala 34:32:@1065.4]
  assign _T_2639 = {valid_12_15,valid_12_14,valid_12_13,valid_12_12,valid_12_11,valid_12_10,valid_12_9,valid_12_8,_T_2631}; // @[Switch.scala 34:32:@1073.4]
  assign _T_2643 = io_inAddr_0 == 4'hd; // @[Switch.scala 30:53:@1076.4]
  assign valid_13_0 = io_inValid_0 & _T_2643; // @[Switch.scala 30:36:@1077.4]
  assign _T_2646 = io_inAddr_1 == 4'hd; // @[Switch.scala 30:53:@1079.4]
  assign valid_13_1 = io_inValid_1 & _T_2646; // @[Switch.scala 30:36:@1080.4]
  assign _T_2649 = io_inAddr_2 == 4'hd; // @[Switch.scala 30:53:@1082.4]
  assign valid_13_2 = io_inValid_2 & _T_2649; // @[Switch.scala 30:36:@1083.4]
  assign _T_2652 = io_inAddr_3 == 4'hd; // @[Switch.scala 30:53:@1085.4]
  assign valid_13_3 = io_inValid_3 & _T_2652; // @[Switch.scala 30:36:@1086.4]
  assign _T_2655 = io_inAddr_4 == 4'hd; // @[Switch.scala 30:53:@1088.4]
  assign valid_13_4 = io_inValid_4 & _T_2655; // @[Switch.scala 30:36:@1089.4]
  assign _T_2658 = io_inAddr_5 == 4'hd; // @[Switch.scala 30:53:@1091.4]
  assign valid_13_5 = io_inValid_5 & _T_2658; // @[Switch.scala 30:36:@1092.4]
  assign _T_2661 = io_inAddr_6 == 4'hd; // @[Switch.scala 30:53:@1094.4]
  assign valid_13_6 = io_inValid_6 & _T_2661; // @[Switch.scala 30:36:@1095.4]
  assign _T_2664 = io_inAddr_7 == 4'hd; // @[Switch.scala 30:53:@1097.4]
  assign valid_13_7 = io_inValid_7 & _T_2664; // @[Switch.scala 30:36:@1098.4]
  assign _T_2667 = io_inAddr_8 == 4'hd; // @[Switch.scala 30:53:@1100.4]
  assign valid_13_8 = io_inValid_8 & _T_2667; // @[Switch.scala 30:36:@1101.4]
  assign _T_2670 = io_inAddr_9 == 4'hd; // @[Switch.scala 30:53:@1103.4]
  assign valid_13_9 = io_inValid_9 & _T_2670; // @[Switch.scala 30:36:@1104.4]
  assign _T_2673 = io_inAddr_10 == 4'hd; // @[Switch.scala 30:53:@1106.4]
  assign valid_13_10 = io_inValid_10 & _T_2673; // @[Switch.scala 30:36:@1107.4]
  assign _T_2676 = io_inAddr_11 == 4'hd; // @[Switch.scala 30:53:@1109.4]
  assign valid_13_11 = io_inValid_11 & _T_2676; // @[Switch.scala 30:36:@1110.4]
  assign _T_2679 = io_inAddr_12 == 4'hd; // @[Switch.scala 30:53:@1112.4]
  assign valid_13_12 = io_inValid_12 & _T_2679; // @[Switch.scala 30:36:@1113.4]
  assign _T_2682 = io_inAddr_13 == 4'hd; // @[Switch.scala 30:53:@1115.4]
  assign valid_13_13 = io_inValid_13 & _T_2682; // @[Switch.scala 30:36:@1116.4]
  assign _T_2685 = io_inAddr_14 == 4'hd; // @[Switch.scala 30:53:@1118.4]
  assign valid_13_14 = io_inValid_14 & _T_2685; // @[Switch.scala 30:36:@1119.4]
  assign _T_2688 = io_inAddr_15 == 4'hd; // @[Switch.scala 30:53:@1121.4]
  assign valid_13_15 = io_inValid_15 & _T_2688; // @[Switch.scala 30:36:@1122.4]
  assign _T_2706 = valid_13_14 ? 4'he : 4'hf; // @[Mux.scala 31:69:@1124.4]
  assign _T_2707 = valid_13_13 ? 4'hd : _T_2706; // @[Mux.scala 31:69:@1125.4]
  assign _T_2708 = valid_13_12 ? 4'hc : _T_2707; // @[Mux.scala 31:69:@1126.4]
  assign _T_2709 = valid_13_11 ? 4'hb : _T_2708; // @[Mux.scala 31:69:@1127.4]
  assign _T_2710 = valid_13_10 ? 4'ha : _T_2709; // @[Mux.scala 31:69:@1128.4]
  assign _T_2711 = valid_13_9 ? 4'h9 : _T_2710; // @[Mux.scala 31:69:@1129.4]
  assign _T_2712 = valid_13_8 ? 4'h8 : _T_2711; // @[Mux.scala 31:69:@1130.4]
  assign _T_2713 = valid_13_7 ? 4'h7 : _T_2712; // @[Mux.scala 31:69:@1131.4]
  assign _T_2714 = valid_13_6 ? 4'h6 : _T_2713; // @[Mux.scala 31:69:@1132.4]
  assign _T_2715 = valid_13_5 ? 4'h5 : _T_2714; // @[Mux.scala 31:69:@1133.4]
  assign _T_2716 = valid_13_4 ? 4'h4 : _T_2715; // @[Mux.scala 31:69:@1134.4]
  assign _T_2717 = valid_13_3 ? 4'h3 : _T_2716; // @[Mux.scala 31:69:@1135.4]
  assign _T_2718 = valid_13_2 ? 4'h2 : _T_2717; // @[Mux.scala 31:69:@1136.4]
  assign _T_2719 = valid_13_1 ? 4'h1 : _T_2718; // @[Mux.scala 31:69:@1137.4]
  assign select_13 = valid_13_0 ? 4'h0 : _T_2719; // @[Mux.scala 31:69:@1138.4]
  assign _GEN_209 = 4'h1 == select_13 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@1140.4]
  assign _GEN_210 = 4'h2 == select_13 ? io_inData_2 : _GEN_209; // @[Switch.scala 33:19:@1140.4]
  assign _GEN_211 = 4'h3 == select_13 ? io_inData_3 : _GEN_210; // @[Switch.scala 33:19:@1140.4]
  assign _GEN_212 = 4'h4 == select_13 ? io_inData_4 : _GEN_211; // @[Switch.scala 33:19:@1140.4]
  assign _GEN_213 = 4'h5 == select_13 ? io_inData_5 : _GEN_212; // @[Switch.scala 33:19:@1140.4]
  assign _GEN_214 = 4'h6 == select_13 ? io_inData_6 : _GEN_213; // @[Switch.scala 33:19:@1140.4]
  assign _GEN_215 = 4'h7 == select_13 ? io_inData_7 : _GEN_214; // @[Switch.scala 33:19:@1140.4]
  assign _GEN_216 = 4'h8 == select_13 ? io_inData_8 : _GEN_215; // @[Switch.scala 33:19:@1140.4]
  assign _GEN_217 = 4'h9 == select_13 ? io_inData_9 : _GEN_216; // @[Switch.scala 33:19:@1140.4]
  assign _GEN_218 = 4'ha == select_13 ? io_inData_10 : _GEN_217; // @[Switch.scala 33:19:@1140.4]
  assign _GEN_219 = 4'hb == select_13 ? io_inData_11 : _GEN_218; // @[Switch.scala 33:19:@1140.4]
  assign _GEN_220 = 4'hc == select_13 ? io_inData_12 : _GEN_219; // @[Switch.scala 33:19:@1140.4]
  assign _GEN_221 = 4'hd == select_13 ? io_inData_13 : _GEN_220; // @[Switch.scala 33:19:@1140.4]
  assign _GEN_222 = 4'he == select_13 ? io_inData_14 : _GEN_221; // @[Switch.scala 33:19:@1140.4]
  assign _T_2728 = {valid_13_7,valid_13_6,valid_13_5,valid_13_4,valid_13_3,valid_13_2,valid_13_1,valid_13_0}; // @[Switch.scala 34:32:@1147.4]
  assign _T_2736 = {valid_13_15,valid_13_14,valid_13_13,valid_13_12,valid_13_11,valid_13_10,valid_13_9,valid_13_8,_T_2728}; // @[Switch.scala 34:32:@1155.4]
  assign _T_2740 = io_inAddr_0 == 4'he; // @[Switch.scala 30:53:@1158.4]
  assign valid_14_0 = io_inValid_0 & _T_2740; // @[Switch.scala 30:36:@1159.4]
  assign _T_2743 = io_inAddr_1 == 4'he; // @[Switch.scala 30:53:@1161.4]
  assign valid_14_1 = io_inValid_1 & _T_2743; // @[Switch.scala 30:36:@1162.4]
  assign _T_2746 = io_inAddr_2 == 4'he; // @[Switch.scala 30:53:@1164.4]
  assign valid_14_2 = io_inValid_2 & _T_2746; // @[Switch.scala 30:36:@1165.4]
  assign _T_2749 = io_inAddr_3 == 4'he; // @[Switch.scala 30:53:@1167.4]
  assign valid_14_3 = io_inValid_3 & _T_2749; // @[Switch.scala 30:36:@1168.4]
  assign _T_2752 = io_inAddr_4 == 4'he; // @[Switch.scala 30:53:@1170.4]
  assign valid_14_4 = io_inValid_4 & _T_2752; // @[Switch.scala 30:36:@1171.4]
  assign _T_2755 = io_inAddr_5 == 4'he; // @[Switch.scala 30:53:@1173.4]
  assign valid_14_5 = io_inValid_5 & _T_2755; // @[Switch.scala 30:36:@1174.4]
  assign _T_2758 = io_inAddr_6 == 4'he; // @[Switch.scala 30:53:@1176.4]
  assign valid_14_6 = io_inValid_6 & _T_2758; // @[Switch.scala 30:36:@1177.4]
  assign _T_2761 = io_inAddr_7 == 4'he; // @[Switch.scala 30:53:@1179.4]
  assign valid_14_7 = io_inValid_7 & _T_2761; // @[Switch.scala 30:36:@1180.4]
  assign _T_2764 = io_inAddr_8 == 4'he; // @[Switch.scala 30:53:@1182.4]
  assign valid_14_8 = io_inValid_8 & _T_2764; // @[Switch.scala 30:36:@1183.4]
  assign _T_2767 = io_inAddr_9 == 4'he; // @[Switch.scala 30:53:@1185.4]
  assign valid_14_9 = io_inValid_9 & _T_2767; // @[Switch.scala 30:36:@1186.4]
  assign _T_2770 = io_inAddr_10 == 4'he; // @[Switch.scala 30:53:@1188.4]
  assign valid_14_10 = io_inValid_10 & _T_2770; // @[Switch.scala 30:36:@1189.4]
  assign _T_2773 = io_inAddr_11 == 4'he; // @[Switch.scala 30:53:@1191.4]
  assign valid_14_11 = io_inValid_11 & _T_2773; // @[Switch.scala 30:36:@1192.4]
  assign _T_2776 = io_inAddr_12 == 4'he; // @[Switch.scala 30:53:@1194.4]
  assign valid_14_12 = io_inValid_12 & _T_2776; // @[Switch.scala 30:36:@1195.4]
  assign _T_2779 = io_inAddr_13 == 4'he; // @[Switch.scala 30:53:@1197.4]
  assign valid_14_13 = io_inValid_13 & _T_2779; // @[Switch.scala 30:36:@1198.4]
  assign _T_2782 = io_inAddr_14 == 4'he; // @[Switch.scala 30:53:@1200.4]
  assign valid_14_14 = io_inValid_14 & _T_2782; // @[Switch.scala 30:36:@1201.4]
  assign _T_2785 = io_inAddr_15 == 4'he; // @[Switch.scala 30:53:@1203.4]
  assign valid_14_15 = io_inValid_15 & _T_2785; // @[Switch.scala 30:36:@1204.4]
  assign _T_2803 = valid_14_14 ? 4'he : 4'hf; // @[Mux.scala 31:69:@1206.4]
  assign _T_2804 = valid_14_13 ? 4'hd : _T_2803; // @[Mux.scala 31:69:@1207.4]
  assign _T_2805 = valid_14_12 ? 4'hc : _T_2804; // @[Mux.scala 31:69:@1208.4]
  assign _T_2806 = valid_14_11 ? 4'hb : _T_2805; // @[Mux.scala 31:69:@1209.4]
  assign _T_2807 = valid_14_10 ? 4'ha : _T_2806; // @[Mux.scala 31:69:@1210.4]
  assign _T_2808 = valid_14_9 ? 4'h9 : _T_2807; // @[Mux.scala 31:69:@1211.4]
  assign _T_2809 = valid_14_8 ? 4'h8 : _T_2808; // @[Mux.scala 31:69:@1212.4]
  assign _T_2810 = valid_14_7 ? 4'h7 : _T_2809; // @[Mux.scala 31:69:@1213.4]
  assign _T_2811 = valid_14_6 ? 4'h6 : _T_2810; // @[Mux.scala 31:69:@1214.4]
  assign _T_2812 = valid_14_5 ? 4'h5 : _T_2811; // @[Mux.scala 31:69:@1215.4]
  assign _T_2813 = valid_14_4 ? 4'h4 : _T_2812; // @[Mux.scala 31:69:@1216.4]
  assign _T_2814 = valid_14_3 ? 4'h3 : _T_2813; // @[Mux.scala 31:69:@1217.4]
  assign _T_2815 = valid_14_2 ? 4'h2 : _T_2814; // @[Mux.scala 31:69:@1218.4]
  assign _T_2816 = valid_14_1 ? 4'h1 : _T_2815; // @[Mux.scala 31:69:@1219.4]
  assign select_14 = valid_14_0 ? 4'h0 : _T_2816; // @[Mux.scala 31:69:@1220.4]
  assign _GEN_225 = 4'h1 == select_14 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@1222.4]
  assign _GEN_226 = 4'h2 == select_14 ? io_inData_2 : _GEN_225; // @[Switch.scala 33:19:@1222.4]
  assign _GEN_227 = 4'h3 == select_14 ? io_inData_3 : _GEN_226; // @[Switch.scala 33:19:@1222.4]
  assign _GEN_228 = 4'h4 == select_14 ? io_inData_4 : _GEN_227; // @[Switch.scala 33:19:@1222.4]
  assign _GEN_229 = 4'h5 == select_14 ? io_inData_5 : _GEN_228; // @[Switch.scala 33:19:@1222.4]
  assign _GEN_230 = 4'h6 == select_14 ? io_inData_6 : _GEN_229; // @[Switch.scala 33:19:@1222.4]
  assign _GEN_231 = 4'h7 == select_14 ? io_inData_7 : _GEN_230; // @[Switch.scala 33:19:@1222.4]
  assign _GEN_232 = 4'h8 == select_14 ? io_inData_8 : _GEN_231; // @[Switch.scala 33:19:@1222.4]
  assign _GEN_233 = 4'h9 == select_14 ? io_inData_9 : _GEN_232; // @[Switch.scala 33:19:@1222.4]
  assign _GEN_234 = 4'ha == select_14 ? io_inData_10 : _GEN_233; // @[Switch.scala 33:19:@1222.4]
  assign _GEN_235 = 4'hb == select_14 ? io_inData_11 : _GEN_234; // @[Switch.scala 33:19:@1222.4]
  assign _GEN_236 = 4'hc == select_14 ? io_inData_12 : _GEN_235; // @[Switch.scala 33:19:@1222.4]
  assign _GEN_237 = 4'hd == select_14 ? io_inData_13 : _GEN_236; // @[Switch.scala 33:19:@1222.4]
  assign _GEN_238 = 4'he == select_14 ? io_inData_14 : _GEN_237; // @[Switch.scala 33:19:@1222.4]
  assign _T_2825 = {valid_14_7,valid_14_6,valid_14_5,valid_14_4,valid_14_3,valid_14_2,valid_14_1,valid_14_0}; // @[Switch.scala 34:32:@1229.4]
  assign _T_2833 = {valid_14_15,valid_14_14,valid_14_13,valid_14_12,valid_14_11,valid_14_10,valid_14_9,valid_14_8,_T_2825}; // @[Switch.scala 34:32:@1237.4]
  assign _T_2837 = io_inAddr_0 == 4'hf; // @[Switch.scala 30:53:@1240.4]
  assign valid_15_0 = io_inValid_0 & _T_2837; // @[Switch.scala 30:36:@1241.4]
  assign _T_2840 = io_inAddr_1 == 4'hf; // @[Switch.scala 30:53:@1243.4]
  assign valid_15_1 = io_inValid_1 & _T_2840; // @[Switch.scala 30:36:@1244.4]
  assign _T_2843 = io_inAddr_2 == 4'hf; // @[Switch.scala 30:53:@1246.4]
  assign valid_15_2 = io_inValid_2 & _T_2843; // @[Switch.scala 30:36:@1247.4]
  assign _T_2846 = io_inAddr_3 == 4'hf; // @[Switch.scala 30:53:@1249.4]
  assign valid_15_3 = io_inValid_3 & _T_2846; // @[Switch.scala 30:36:@1250.4]
  assign _T_2849 = io_inAddr_4 == 4'hf; // @[Switch.scala 30:53:@1252.4]
  assign valid_15_4 = io_inValid_4 & _T_2849; // @[Switch.scala 30:36:@1253.4]
  assign _T_2852 = io_inAddr_5 == 4'hf; // @[Switch.scala 30:53:@1255.4]
  assign valid_15_5 = io_inValid_5 & _T_2852; // @[Switch.scala 30:36:@1256.4]
  assign _T_2855 = io_inAddr_6 == 4'hf; // @[Switch.scala 30:53:@1258.4]
  assign valid_15_6 = io_inValid_6 & _T_2855; // @[Switch.scala 30:36:@1259.4]
  assign _T_2858 = io_inAddr_7 == 4'hf; // @[Switch.scala 30:53:@1261.4]
  assign valid_15_7 = io_inValid_7 & _T_2858; // @[Switch.scala 30:36:@1262.4]
  assign _T_2861 = io_inAddr_8 == 4'hf; // @[Switch.scala 30:53:@1264.4]
  assign valid_15_8 = io_inValid_8 & _T_2861; // @[Switch.scala 30:36:@1265.4]
  assign _T_2864 = io_inAddr_9 == 4'hf; // @[Switch.scala 30:53:@1267.4]
  assign valid_15_9 = io_inValid_9 & _T_2864; // @[Switch.scala 30:36:@1268.4]
  assign _T_2867 = io_inAddr_10 == 4'hf; // @[Switch.scala 30:53:@1270.4]
  assign valid_15_10 = io_inValid_10 & _T_2867; // @[Switch.scala 30:36:@1271.4]
  assign _T_2870 = io_inAddr_11 == 4'hf; // @[Switch.scala 30:53:@1273.4]
  assign valid_15_11 = io_inValid_11 & _T_2870; // @[Switch.scala 30:36:@1274.4]
  assign _T_2873 = io_inAddr_12 == 4'hf; // @[Switch.scala 30:53:@1276.4]
  assign valid_15_12 = io_inValid_12 & _T_2873; // @[Switch.scala 30:36:@1277.4]
  assign _T_2876 = io_inAddr_13 == 4'hf; // @[Switch.scala 30:53:@1279.4]
  assign valid_15_13 = io_inValid_13 & _T_2876; // @[Switch.scala 30:36:@1280.4]
  assign _T_2879 = io_inAddr_14 == 4'hf; // @[Switch.scala 30:53:@1282.4]
  assign valid_15_14 = io_inValid_14 & _T_2879; // @[Switch.scala 30:36:@1283.4]
  assign _T_2882 = io_inAddr_15 == 4'hf; // @[Switch.scala 30:53:@1285.4]
  assign valid_15_15 = io_inValid_15 & _T_2882; // @[Switch.scala 30:36:@1286.4]
  assign _T_2900 = valid_15_14 ? 4'he : 4'hf; // @[Mux.scala 31:69:@1288.4]
  assign _T_2901 = valid_15_13 ? 4'hd : _T_2900; // @[Mux.scala 31:69:@1289.4]
  assign _T_2902 = valid_15_12 ? 4'hc : _T_2901; // @[Mux.scala 31:69:@1290.4]
  assign _T_2903 = valid_15_11 ? 4'hb : _T_2902; // @[Mux.scala 31:69:@1291.4]
  assign _T_2904 = valid_15_10 ? 4'ha : _T_2903; // @[Mux.scala 31:69:@1292.4]
  assign _T_2905 = valid_15_9 ? 4'h9 : _T_2904; // @[Mux.scala 31:69:@1293.4]
  assign _T_2906 = valid_15_8 ? 4'h8 : _T_2905; // @[Mux.scala 31:69:@1294.4]
  assign _T_2907 = valid_15_7 ? 4'h7 : _T_2906; // @[Mux.scala 31:69:@1295.4]
  assign _T_2908 = valid_15_6 ? 4'h6 : _T_2907; // @[Mux.scala 31:69:@1296.4]
  assign _T_2909 = valid_15_5 ? 4'h5 : _T_2908; // @[Mux.scala 31:69:@1297.4]
  assign _T_2910 = valid_15_4 ? 4'h4 : _T_2909; // @[Mux.scala 31:69:@1298.4]
  assign _T_2911 = valid_15_3 ? 4'h3 : _T_2910; // @[Mux.scala 31:69:@1299.4]
  assign _T_2912 = valid_15_2 ? 4'h2 : _T_2911; // @[Mux.scala 31:69:@1300.4]
  assign _T_2913 = valid_15_1 ? 4'h1 : _T_2912; // @[Mux.scala 31:69:@1301.4]
  assign select_15 = valid_15_0 ? 4'h0 : _T_2913; // @[Mux.scala 31:69:@1302.4]
  assign _GEN_241 = 4'h1 == select_15 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@1304.4]
  assign _GEN_242 = 4'h2 == select_15 ? io_inData_2 : _GEN_241; // @[Switch.scala 33:19:@1304.4]
  assign _GEN_243 = 4'h3 == select_15 ? io_inData_3 : _GEN_242; // @[Switch.scala 33:19:@1304.4]
  assign _GEN_244 = 4'h4 == select_15 ? io_inData_4 : _GEN_243; // @[Switch.scala 33:19:@1304.4]
  assign _GEN_245 = 4'h5 == select_15 ? io_inData_5 : _GEN_244; // @[Switch.scala 33:19:@1304.4]
  assign _GEN_246 = 4'h6 == select_15 ? io_inData_6 : _GEN_245; // @[Switch.scala 33:19:@1304.4]
  assign _GEN_247 = 4'h7 == select_15 ? io_inData_7 : _GEN_246; // @[Switch.scala 33:19:@1304.4]
  assign _GEN_248 = 4'h8 == select_15 ? io_inData_8 : _GEN_247; // @[Switch.scala 33:19:@1304.4]
  assign _GEN_249 = 4'h9 == select_15 ? io_inData_9 : _GEN_248; // @[Switch.scala 33:19:@1304.4]
  assign _GEN_250 = 4'ha == select_15 ? io_inData_10 : _GEN_249; // @[Switch.scala 33:19:@1304.4]
  assign _GEN_251 = 4'hb == select_15 ? io_inData_11 : _GEN_250; // @[Switch.scala 33:19:@1304.4]
  assign _GEN_252 = 4'hc == select_15 ? io_inData_12 : _GEN_251; // @[Switch.scala 33:19:@1304.4]
  assign _GEN_253 = 4'hd == select_15 ? io_inData_13 : _GEN_252; // @[Switch.scala 33:19:@1304.4]
  assign _GEN_254 = 4'he == select_15 ? io_inData_14 : _GEN_253; // @[Switch.scala 33:19:@1304.4]
  assign _T_2922 = {valid_15_7,valid_15_6,valid_15_5,valid_15_4,valid_15_3,valid_15_2,valid_15_1,valid_15_0}; // @[Switch.scala 34:32:@1311.4]
  assign _T_2930 = {valid_15_15,valid_15_14,valid_15_13,valid_15_12,valid_15_11,valid_15_10,valid_15_9,valid_15_8,_T_2922}; // @[Switch.scala 34:32:@1319.4]
  assign _T_4164 = select_0 == 4'h0; // @[Switch.scala 41:52:@1323.4]
  assign output_0_0 = io_outValid_0 & _T_4164; // @[Switch.scala 41:38:@1324.4]
  assign _T_4167 = select_1 == 4'h0; // @[Switch.scala 41:52:@1326.4]
  assign output_0_1 = io_outValid_1 & _T_4167; // @[Switch.scala 41:38:@1327.4]
  assign _T_4170 = select_2 == 4'h0; // @[Switch.scala 41:52:@1329.4]
  assign output_0_2 = io_outValid_2 & _T_4170; // @[Switch.scala 41:38:@1330.4]
  assign _T_4173 = select_3 == 4'h0; // @[Switch.scala 41:52:@1332.4]
  assign output_0_3 = io_outValid_3 & _T_4173; // @[Switch.scala 41:38:@1333.4]
  assign _T_4176 = select_4 == 4'h0; // @[Switch.scala 41:52:@1335.4]
  assign output_0_4 = io_outValid_4 & _T_4176; // @[Switch.scala 41:38:@1336.4]
  assign _T_4179 = select_5 == 4'h0; // @[Switch.scala 41:52:@1338.4]
  assign output_0_5 = io_outValid_5 & _T_4179; // @[Switch.scala 41:38:@1339.4]
  assign _T_4182 = select_6 == 4'h0; // @[Switch.scala 41:52:@1341.4]
  assign output_0_6 = io_outValid_6 & _T_4182; // @[Switch.scala 41:38:@1342.4]
  assign _T_4185 = select_7 == 4'h0; // @[Switch.scala 41:52:@1344.4]
  assign output_0_7 = io_outValid_7 & _T_4185; // @[Switch.scala 41:38:@1345.4]
  assign _T_4188 = select_8 == 4'h0; // @[Switch.scala 41:52:@1347.4]
  assign output_0_8 = io_outValid_8 & _T_4188; // @[Switch.scala 41:38:@1348.4]
  assign _T_4191 = select_9 == 4'h0; // @[Switch.scala 41:52:@1350.4]
  assign output_0_9 = io_outValid_9 & _T_4191; // @[Switch.scala 41:38:@1351.4]
  assign _T_4194 = select_10 == 4'h0; // @[Switch.scala 41:52:@1353.4]
  assign output_0_10 = io_outValid_10 & _T_4194; // @[Switch.scala 41:38:@1354.4]
  assign _T_4197 = select_11 == 4'h0; // @[Switch.scala 41:52:@1356.4]
  assign output_0_11 = io_outValid_11 & _T_4197; // @[Switch.scala 41:38:@1357.4]
  assign _T_4200 = select_12 == 4'h0; // @[Switch.scala 41:52:@1359.4]
  assign output_0_12 = io_outValid_12 & _T_4200; // @[Switch.scala 41:38:@1360.4]
  assign _T_4203 = select_13 == 4'h0; // @[Switch.scala 41:52:@1362.4]
  assign output_0_13 = io_outValid_13 & _T_4203; // @[Switch.scala 41:38:@1363.4]
  assign _T_4206 = select_14 == 4'h0; // @[Switch.scala 41:52:@1365.4]
  assign output_0_14 = io_outValid_14 & _T_4206; // @[Switch.scala 41:38:@1366.4]
  assign _T_4209 = select_15 == 4'h0; // @[Switch.scala 41:52:@1368.4]
  assign output_0_15 = io_outValid_15 & _T_4209; // @[Switch.scala 41:38:@1369.4]
  assign _T_4217 = {output_0_7,output_0_6,output_0_5,output_0_4,output_0_3,output_0_2,output_0_1,output_0_0}; // @[Switch.scala 43:31:@1377.4]
  assign _T_4225 = {output_0_15,output_0_14,output_0_13,output_0_12,output_0_11,output_0_10,output_0_9,output_0_8,_T_4217}; // @[Switch.scala 43:31:@1385.4]
  assign _T_4229 = select_0 == 4'h1; // @[Switch.scala 41:52:@1388.4]
  assign output_1_0 = io_outValid_0 & _T_4229; // @[Switch.scala 41:38:@1389.4]
  assign _T_4232 = select_1 == 4'h1; // @[Switch.scala 41:52:@1391.4]
  assign output_1_1 = io_outValid_1 & _T_4232; // @[Switch.scala 41:38:@1392.4]
  assign _T_4235 = select_2 == 4'h1; // @[Switch.scala 41:52:@1394.4]
  assign output_1_2 = io_outValid_2 & _T_4235; // @[Switch.scala 41:38:@1395.4]
  assign _T_4238 = select_3 == 4'h1; // @[Switch.scala 41:52:@1397.4]
  assign output_1_3 = io_outValid_3 & _T_4238; // @[Switch.scala 41:38:@1398.4]
  assign _T_4241 = select_4 == 4'h1; // @[Switch.scala 41:52:@1400.4]
  assign output_1_4 = io_outValid_4 & _T_4241; // @[Switch.scala 41:38:@1401.4]
  assign _T_4244 = select_5 == 4'h1; // @[Switch.scala 41:52:@1403.4]
  assign output_1_5 = io_outValid_5 & _T_4244; // @[Switch.scala 41:38:@1404.4]
  assign _T_4247 = select_6 == 4'h1; // @[Switch.scala 41:52:@1406.4]
  assign output_1_6 = io_outValid_6 & _T_4247; // @[Switch.scala 41:38:@1407.4]
  assign _T_4250 = select_7 == 4'h1; // @[Switch.scala 41:52:@1409.4]
  assign output_1_7 = io_outValid_7 & _T_4250; // @[Switch.scala 41:38:@1410.4]
  assign _T_4253 = select_8 == 4'h1; // @[Switch.scala 41:52:@1412.4]
  assign output_1_8 = io_outValid_8 & _T_4253; // @[Switch.scala 41:38:@1413.4]
  assign _T_4256 = select_9 == 4'h1; // @[Switch.scala 41:52:@1415.4]
  assign output_1_9 = io_outValid_9 & _T_4256; // @[Switch.scala 41:38:@1416.4]
  assign _T_4259 = select_10 == 4'h1; // @[Switch.scala 41:52:@1418.4]
  assign output_1_10 = io_outValid_10 & _T_4259; // @[Switch.scala 41:38:@1419.4]
  assign _T_4262 = select_11 == 4'h1; // @[Switch.scala 41:52:@1421.4]
  assign output_1_11 = io_outValid_11 & _T_4262; // @[Switch.scala 41:38:@1422.4]
  assign _T_4265 = select_12 == 4'h1; // @[Switch.scala 41:52:@1424.4]
  assign output_1_12 = io_outValid_12 & _T_4265; // @[Switch.scala 41:38:@1425.4]
  assign _T_4268 = select_13 == 4'h1; // @[Switch.scala 41:52:@1427.4]
  assign output_1_13 = io_outValid_13 & _T_4268; // @[Switch.scala 41:38:@1428.4]
  assign _T_4271 = select_14 == 4'h1; // @[Switch.scala 41:52:@1430.4]
  assign output_1_14 = io_outValid_14 & _T_4271; // @[Switch.scala 41:38:@1431.4]
  assign _T_4274 = select_15 == 4'h1; // @[Switch.scala 41:52:@1433.4]
  assign output_1_15 = io_outValid_15 & _T_4274; // @[Switch.scala 41:38:@1434.4]
  assign _T_4282 = {output_1_7,output_1_6,output_1_5,output_1_4,output_1_3,output_1_2,output_1_1,output_1_0}; // @[Switch.scala 43:31:@1442.4]
  assign _T_4290 = {output_1_15,output_1_14,output_1_13,output_1_12,output_1_11,output_1_10,output_1_9,output_1_8,_T_4282}; // @[Switch.scala 43:31:@1450.4]
  assign _T_4294 = select_0 == 4'h2; // @[Switch.scala 41:52:@1453.4]
  assign output_2_0 = io_outValid_0 & _T_4294; // @[Switch.scala 41:38:@1454.4]
  assign _T_4297 = select_1 == 4'h2; // @[Switch.scala 41:52:@1456.4]
  assign output_2_1 = io_outValid_1 & _T_4297; // @[Switch.scala 41:38:@1457.4]
  assign _T_4300 = select_2 == 4'h2; // @[Switch.scala 41:52:@1459.4]
  assign output_2_2 = io_outValid_2 & _T_4300; // @[Switch.scala 41:38:@1460.4]
  assign _T_4303 = select_3 == 4'h2; // @[Switch.scala 41:52:@1462.4]
  assign output_2_3 = io_outValid_3 & _T_4303; // @[Switch.scala 41:38:@1463.4]
  assign _T_4306 = select_4 == 4'h2; // @[Switch.scala 41:52:@1465.4]
  assign output_2_4 = io_outValid_4 & _T_4306; // @[Switch.scala 41:38:@1466.4]
  assign _T_4309 = select_5 == 4'h2; // @[Switch.scala 41:52:@1468.4]
  assign output_2_5 = io_outValid_5 & _T_4309; // @[Switch.scala 41:38:@1469.4]
  assign _T_4312 = select_6 == 4'h2; // @[Switch.scala 41:52:@1471.4]
  assign output_2_6 = io_outValid_6 & _T_4312; // @[Switch.scala 41:38:@1472.4]
  assign _T_4315 = select_7 == 4'h2; // @[Switch.scala 41:52:@1474.4]
  assign output_2_7 = io_outValid_7 & _T_4315; // @[Switch.scala 41:38:@1475.4]
  assign _T_4318 = select_8 == 4'h2; // @[Switch.scala 41:52:@1477.4]
  assign output_2_8 = io_outValid_8 & _T_4318; // @[Switch.scala 41:38:@1478.4]
  assign _T_4321 = select_9 == 4'h2; // @[Switch.scala 41:52:@1480.4]
  assign output_2_9 = io_outValid_9 & _T_4321; // @[Switch.scala 41:38:@1481.4]
  assign _T_4324 = select_10 == 4'h2; // @[Switch.scala 41:52:@1483.4]
  assign output_2_10 = io_outValid_10 & _T_4324; // @[Switch.scala 41:38:@1484.4]
  assign _T_4327 = select_11 == 4'h2; // @[Switch.scala 41:52:@1486.4]
  assign output_2_11 = io_outValid_11 & _T_4327; // @[Switch.scala 41:38:@1487.4]
  assign _T_4330 = select_12 == 4'h2; // @[Switch.scala 41:52:@1489.4]
  assign output_2_12 = io_outValid_12 & _T_4330; // @[Switch.scala 41:38:@1490.4]
  assign _T_4333 = select_13 == 4'h2; // @[Switch.scala 41:52:@1492.4]
  assign output_2_13 = io_outValid_13 & _T_4333; // @[Switch.scala 41:38:@1493.4]
  assign _T_4336 = select_14 == 4'h2; // @[Switch.scala 41:52:@1495.4]
  assign output_2_14 = io_outValid_14 & _T_4336; // @[Switch.scala 41:38:@1496.4]
  assign _T_4339 = select_15 == 4'h2; // @[Switch.scala 41:52:@1498.4]
  assign output_2_15 = io_outValid_15 & _T_4339; // @[Switch.scala 41:38:@1499.4]
  assign _T_4347 = {output_2_7,output_2_6,output_2_5,output_2_4,output_2_3,output_2_2,output_2_1,output_2_0}; // @[Switch.scala 43:31:@1507.4]
  assign _T_4355 = {output_2_15,output_2_14,output_2_13,output_2_12,output_2_11,output_2_10,output_2_9,output_2_8,_T_4347}; // @[Switch.scala 43:31:@1515.4]
  assign _T_4359 = select_0 == 4'h3; // @[Switch.scala 41:52:@1518.4]
  assign output_3_0 = io_outValid_0 & _T_4359; // @[Switch.scala 41:38:@1519.4]
  assign _T_4362 = select_1 == 4'h3; // @[Switch.scala 41:52:@1521.4]
  assign output_3_1 = io_outValid_1 & _T_4362; // @[Switch.scala 41:38:@1522.4]
  assign _T_4365 = select_2 == 4'h3; // @[Switch.scala 41:52:@1524.4]
  assign output_3_2 = io_outValid_2 & _T_4365; // @[Switch.scala 41:38:@1525.4]
  assign _T_4368 = select_3 == 4'h3; // @[Switch.scala 41:52:@1527.4]
  assign output_3_3 = io_outValid_3 & _T_4368; // @[Switch.scala 41:38:@1528.4]
  assign _T_4371 = select_4 == 4'h3; // @[Switch.scala 41:52:@1530.4]
  assign output_3_4 = io_outValid_4 & _T_4371; // @[Switch.scala 41:38:@1531.4]
  assign _T_4374 = select_5 == 4'h3; // @[Switch.scala 41:52:@1533.4]
  assign output_3_5 = io_outValid_5 & _T_4374; // @[Switch.scala 41:38:@1534.4]
  assign _T_4377 = select_6 == 4'h3; // @[Switch.scala 41:52:@1536.4]
  assign output_3_6 = io_outValid_6 & _T_4377; // @[Switch.scala 41:38:@1537.4]
  assign _T_4380 = select_7 == 4'h3; // @[Switch.scala 41:52:@1539.4]
  assign output_3_7 = io_outValid_7 & _T_4380; // @[Switch.scala 41:38:@1540.4]
  assign _T_4383 = select_8 == 4'h3; // @[Switch.scala 41:52:@1542.4]
  assign output_3_8 = io_outValid_8 & _T_4383; // @[Switch.scala 41:38:@1543.4]
  assign _T_4386 = select_9 == 4'h3; // @[Switch.scala 41:52:@1545.4]
  assign output_3_9 = io_outValid_9 & _T_4386; // @[Switch.scala 41:38:@1546.4]
  assign _T_4389 = select_10 == 4'h3; // @[Switch.scala 41:52:@1548.4]
  assign output_3_10 = io_outValid_10 & _T_4389; // @[Switch.scala 41:38:@1549.4]
  assign _T_4392 = select_11 == 4'h3; // @[Switch.scala 41:52:@1551.4]
  assign output_3_11 = io_outValid_11 & _T_4392; // @[Switch.scala 41:38:@1552.4]
  assign _T_4395 = select_12 == 4'h3; // @[Switch.scala 41:52:@1554.4]
  assign output_3_12 = io_outValid_12 & _T_4395; // @[Switch.scala 41:38:@1555.4]
  assign _T_4398 = select_13 == 4'h3; // @[Switch.scala 41:52:@1557.4]
  assign output_3_13 = io_outValid_13 & _T_4398; // @[Switch.scala 41:38:@1558.4]
  assign _T_4401 = select_14 == 4'h3; // @[Switch.scala 41:52:@1560.4]
  assign output_3_14 = io_outValid_14 & _T_4401; // @[Switch.scala 41:38:@1561.4]
  assign _T_4404 = select_15 == 4'h3; // @[Switch.scala 41:52:@1563.4]
  assign output_3_15 = io_outValid_15 & _T_4404; // @[Switch.scala 41:38:@1564.4]
  assign _T_4412 = {output_3_7,output_3_6,output_3_5,output_3_4,output_3_3,output_3_2,output_3_1,output_3_0}; // @[Switch.scala 43:31:@1572.4]
  assign _T_4420 = {output_3_15,output_3_14,output_3_13,output_3_12,output_3_11,output_3_10,output_3_9,output_3_8,_T_4412}; // @[Switch.scala 43:31:@1580.4]
  assign _T_4424 = select_0 == 4'h4; // @[Switch.scala 41:52:@1583.4]
  assign output_4_0 = io_outValid_0 & _T_4424; // @[Switch.scala 41:38:@1584.4]
  assign _T_4427 = select_1 == 4'h4; // @[Switch.scala 41:52:@1586.4]
  assign output_4_1 = io_outValid_1 & _T_4427; // @[Switch.scala 41:38:@1587.4]
  assign _T_4430 = select_2 == 4'h4; // @[Switch.scala 41:52:@1589.4]
  assign output_4_2 = io_outValid_2 & _T_4430; // @[Switch.scala 41:38:@1590.4]
  assign _T_4433 = select_3 == 4'h4; // @[Switch.scala 41:52:@1592.4]
  assign output_4_3 = io_outValid_3 & _T_4433; // @[Switch.scala 41:38:@1593.4]
  assign _T_4436 = select_4 == 4'h4; // @[Switch.scala 41:52:@1595.4]
  assign output_4_4 = io_outValid_4 & _T_4436; // @[Switch.scala 41:38:@1596.4]
  assign _T_4439 = select_5 == 4'h4; // @[Switch.scala 41:52:@1598.4]
  assign output_4_5 = io_outValid_5 & _T_4439; // @[Switch.scala 41:38:@1599.4]
  assign _T_4442 = select_6 == 4'h4; // @[Switch.scala 41:52:@1601.4]
  assign output_4_6 = io_outValid_6 & _T_4442; // @[Switch.scala 41:38:@1602.4]
  assign _T_4445 = select_7 == 4'h4; // @[Switch.scala 41:52:@1604.4]
  assign output_4_7 = io_outValid_7 & _T_4445; // @[Switch.scala 41:38:@1605.4]
  assign _T_4448 = select_8 == 4'h4; // @[Switch.scala 41:52:@1607.4]
  assign output_4_8 = io_outValid_8 & _T_4448; // @[Switch.scala 41:38:@1608.4]
  assign _T_4451 = select_9 == 4'h4; // @[Switch.scala 41:52:@1610.4]
  assign output_4_9 = io_outValid_9 & _T_4451; // @[Switch.scala 41:38:@1611.4]
  assign _T_4454 = select_10 == 4'h4; // @[Switch.scala 41:52:@1613.4]
  assign output_4_10 = io_outValid_10 & _T_4454; // @[Switch.scala 41:38:@1614.4]
  assign _T_4457 = select_11 == 4'h4; // @[Switch.scala 41:52:@1616.4]
  assign output_4_11 = io_outValid_11 & _T_4457; // @[Switch.scala 41:38:@1617.4]
  assign _T_4460 = select_12 == 4'h4; // @[Switch.scala 41:52:@1619.4]
  assign output_4_12 = io_outValid_12 & _T_4460; // @[Switch.scala 41:38:@1620.4]
  assign _T_4463 = select_13 == 4'h4; // @[Switch.scala 41:52:@1622.4]
  assign output_4_13 = io_outValid_13 & _T_4463; // @[Switch.scala 41:38:@1623.4]
  assign _T_4466 = select_14 == 4'h4; // @[Switch.scala 41:52:@1625.4]
  assign output_4_14 = io_outValid_14 & _T_4466; // @[Switch.scala 41:38:@1626.4]
  assign _T_4469 = select_15 == 4'h4; // @[Switch.scala 41:52:@1628.4]
  assign output_4_15 = io_outValid_15 & _T_4469; // @[Switch.scala 41:38:@1629.4]
  assign _T_4477 = {output_4_7,output_4_6,output_4_5,output_4_4,output_4_3,output_4_2,output_4_1,output_4_0}; // @[Switch.scala 43:31:@1637.4]
  assign _T_4485 = {output_4_15,output_4_14,output_4_13,output_4_12,output_4_11,output_4_10,output_4_9,output_4_8,_T_4477}; // @[Switch.scala 43:31:@1645.4]
  assign _T_4489 = select_0 == 4'h5; // @[Switch.scala 41:52:@1648.4]
  assign output_5_0 = io_outValid_0 & _T_4489; // @[Switch.scala 41:38:@1649.4]
  assign _T_4492 = select_1 == 4'h5; // @[Switch.scala 41:52:@1651.4]
  assign output_5_1 = io_outValid_1 & _T_4492; // @[Switch.scala 41:38:@1652.4]
  assign _T_4495 = select_2 == 4'h5; // @[Switch.scala 41:52:@1654.4]
  assign output_5_2 = io_outValid_2 & _T_4495; // @[Switch.scala 41:38:@1655.4]
  assign _T_4498 = select_3 == 4'h5; // @[Switch.scala 41:52:@1657.4]
  assign output_5_3 = io_outValid_3 & _T_4498; // @[Switch.scala 41:38:@1658.4]
  assign _T_4501 = select_4 == 4'h5; // @[Switch.scala 41:52:@1660.4]
  assign output_5_4 = io_outValid_4 & _T_4501; // @[Switch.scala 41:38:@1661.4]
  assign _T_4504 = select_5 == 4'h5; // @[Switch.scala 41:52:@1663.4]
  assign output_5_5 = io_outValid_5 & _T_4504; // @[Switch.scala 41:38:@1664.4]
  assign _T_4507 = select_6 == 4'h5; // @[Switch.scala 41:52:@1666.4]
  assign output_5_6 = io_outValid_6 & _T_4507; // @[Switch.scala 41:38:@1667.4]
  assign _T_4510 = select_7 == 4'h5; // @[Switch.scala 41:52:@1669.4]
  assign output_5_7 = io_outValid_7 & _T_4510; // @[Switch.scala 41:38:@1670.4]
  assign _T_4513 = select_8 == 4'h5; // @[Switch.scala 41:52:@1672.4]
  assign output_5_8 = io_outValid_8 & _T_4513; // @[Switch.scala 41:38:@1673.4]
  assign _T_4516 = select_9 == 4'h5; // @[Switch.scala 41:52:@1675.4]
  assign output_5_9 = io_outValid_9 & _T_4516; // @[Switch.scala 41:38:@1676.4]
  assign _T_4519 = select_10 == 4'h5; // @[Switch.scala 41:52:@1678.4]
  assign output_5_10 = io_outValid_10 & _T_4519; // @[Switch.scala 41:38:@1679.4]
  assign _T_4522 = select_11 == 4'h5; // @[Switch.scala 41:52:@1681.4]
  assign output_5_11 = io_outValid_11 & _T_4522; // @[Switch.scala 41:38:@1682.4]
  assign _T_4525 = select_12 == 4'h5; // @[Switch.scala 41:52:@1684.4]
  assign output_5_12 = io_outValid_12 & _T_4525; // @[Switch.scala 41:38:@1685.4]
  assign _T_4528 = select_13 == 4'h5; // @[Switch.scala 41:52:@1687.4]
  assign output_5_13 = io_outValid_13 & _T_4528; // @[Switch.scala 41:38:@1688.4]
  assign _T_4531 = select_14 == 4'h5; // @[Switch.scala 41:52:@1690.4]
  assign output_5_14 = io_outValid_14 & _T_4531; // @[Switch.scala 41:38:@1691.4]
  assign _T_4534 = select_15 == 4'h5; // @[Switch.scala 41:52:@1693.4]
  assign output_5_15 = io_outValid_15 & _T_4534; // @[Switch.scala 41:38:@1694.4]
  assign _T_4542 = {output_5_7,output_5_6,output_5_5,output_5_4,output_5_3,output_5_2,output_5_1,output_5_0}; // @[Switch.scala 43:31:@1702.4]
  assign _T_4550 = {output_5_15,output_5_14,output_5_13,output_5_12,output_5_11,output_5_10,output_5_9,output_5_8,_T_4542}; // @[Switch.scala 43:31:@1710.4]
  assign _T_4554 = select_0 == 4'h6; // @[Switch.scala 41:52:@1713.4]
  assign output_6_0 = io_outValid_0 & _T_4554; // @[Switch.scala 41:38:@1714.4]
  assign _T_4557 = select_1 == 4'h6; // @[Switch.scala 41:52:@1716.4]
  assign output_6_1 = io_outValid_1 & _T_4557; // @[Switch.scala 41:38:@1717.4]
  assign _T_4560 = select_2 == 4'h6; // @[Switch.scala 41:52:@1719.4]
  assign output_6_2 = io_outValid_2 & _T_4560; // @[Switch.scala 41:38:@1720.4]
  assign _T_4563 = select_3 == 4'h6; // @[Switch.scala 41:52:@1722.4]
  assign output_6_3 = io_outValid_3 & _T_4563; // @[Switch.scala 41:38:@1723.4]
  assign _T_4566 = select_4 == 4'h6; // @[Switch.scala 41:52:@1725.4]
  assign output_6_4 = io_outValid_4 & _T_4566; // @[Switch.scala 41:38:@1726.4]
  assign _T_4569 = select_5 == 4'h6; // @[Switch.scala 41:52:@1728.4]
  assign output_6_5 = io_outValid_5 & _T_4569; // @[Switch.scala 41:38:@1729.4]
  assign _T_4572 = select_6 == 4'h6; // @[Switch.scala 41:52:@1731.4]
  assign output_6_6 = io_outValid_6 & _T_4572; // @[Switch.scala 41:38:@1732.4]
  assign _T_4575 = select_7 == 4'h6; // @[Switch.scala 41:52:@1734.4]
  assign output_6_7 = io_outValid_7 & _T_4575; // @[Switch.scala 41:38:@1735.4]
  assign _T_4578 = select_8 == 4'h6; // @[Switch.scala 41:52:@1737.4]
  assign output_6_8 = io_outValid_8 & _T_4578; // @[Switch.scala 41:38:@1738.4]
  assign _T_4581 = select_9 == 4'h6; // @[Switch.scala 41:52:@1740.4]
  assign output_6_9 = io_outValid_9 & _T_4581; // @[Switch.scala 41:38:@1741.4]
  assign _T_4584 = select_10 == 4'h6; // @[Switch.scala 41:52:@1743.4]
  assign output_6_10 = io_outValid_10 & _T_4584; // @[Switch.scala 41:38:@1744.4]
  assign _T_4587 = select_11 == 4'h6; // @[Switch.scala 41:52:@1746.4]
  assign output_6_11 = io_outValid_11 & _T_4587; // @[Switch.scala 41:38:@1747.4]
  assign _T_4590 = select_12 == 4'h6; // @[Switch.scala 41:52:@1749.4]
  assign output_6_12 = io_outValid_12 & _T_4590; // @[Switch.scala 41:38:@1750.4]
  assign _T_4593 = select_13 == 4'h6; // @[Switch.scala 41:52:@1752.4]
  assign output_6_13 = io_outValid_13 & _T_4593; // @[Switch.scala 41:38:@1753.4]
  assign _T_4596 = select_14 == 4'h6; // @[Switch.scala 41:52:@1755.4]
  assign output_6_14 = io_outValid_14 & _T_4596; // @[Switch.scala 41:38:@1756.4]
  assign _T_4599 = select_15 == 4'h6; // @[Switch.scala 41:52:@1758.4]
  assign output_6_15 = io_outValid_15 & _T_4599; // @[Switch.scala 41:38:@1759.4]
  assign _T_4607 = {output_6_7,output_6_6,output_6_5,output_6_4,output_6_3,output_6_2,output_6_1,output_6_0}; // @[Switch.scala 43:31:@1767.4]
  assign _T_4615 = {output_6_15,output_6_14,output_6_13,output_6_12,output_6_11,output_6_10,output_6_9,output_6_8,_T_4607}; // @[Switch.scala 43:31:@1775.4]
  assign _T_4619 = select_0 == 4'h7; // @[Switch.scala 41:52:@1778.4]
  assign output_7_0 = io_outValid_0 & _T_4619; // @[Switch.scala 41:38:@1779.4]
  assign _T_4622 = select_1 == 4'h7; // @[Switch.scala 41:52:@1781.4]
  assign output_7_1 = io_outValid_1 & _T_4622; // @[Switch.scala 41:38:@1782.4]
  assign _T_4625 = select_2 == 4'h7; // @[Switch.scala 41:52:@1784.4]
  assign output_7_2 = io_outValid_2 & _T_4625; // @[Switch.scala 41:38:@1785.4]
  assign _T_4628 = select_3 == 4'h7; // @[Switch.scala 41:52:@1787.4]
  assign output_7_3 = io_outValid_3 & _T_4628; // @[Switch.scala 41:38:@1788.4]
  assign _T_4631 = select_4 == 4'h7; // @[Switch.scala 41:52:@1790.4]
  assign output_7_4 = io_outValid_4 & _T_4631; // @[Switch.scala 41:38:@1791.4]
  assign _T_4634 = select_5 == 4'h7; // @[Switch.scala 41:52:@1793.4]
  assign output_7_5 = io_outValid_5 & _T_4634; // @[Switch.scala 41:38:@1794.4]
  assign _T_4637 = select_6 == 4'h7; // @[Switch.scala 41:52:@1796.4]
  assign output_7_6 = io_outValid_6 & _T_4637; // @[Switch.scala 41:38:@1797.4]
  assign _T_4640 = select_7 == 4'h7; // @[Switch.scala 41:52:@1799.4]
  assign output_7_7 = io_outValid_7 & _T_4640; // @[Switch.scala 41:38:@1800.4]
  assign _T_4643 = select_8 == 4'h7; // @[Switch.scala 41:52:@1802.4]
  assign output_7_8 = io_outValid_8 & _T_4643; // @[Switch.scala 41:38:@1803.4]
  assign _T_4646 = select_9 == 4'h7; // @[Switch.scala 41:52:@1805.4]
  assign output_7_9 = io_outValid_9 & _T_4646; // @[Switch.scala 41:38:@1806.4]
  assign _T_4649 = select_10 == 4'h7; // @[Switch.scala 41:52:@1808.4]
  assign output_7_10 = io_outValid_10 & _T_4649; // @[Switch.scala 41:38:@1809.4]
  assign _T_4652 = select_11 == 4'h7; // @[Switch.scala 41:52:@1811.4]
  assign output_7_11 = io_outValid_11 & _T_4652; // @[Switch.scala 41:38:@1812.4]
  assign _T_4655 = select_12 == 4'h7; // @[Switch.scala 41:52:@1814.4]
  assign output_7_12 = io_outValid_12 & _T_4655; // @[Switch.scala 41:38:@1815.4]
  assign _T_4658 = select_13 == 4'h7; // @[Switch.scala 41:52:@1817.4]
  assign output_7_13 = io_outValid_13 & _T_4658; // @[Switch.scala 41:38:@1818.4]
  assign _T_4661 = select_14 == 4'h7; // @[Switch.scala 41:52:@1820.4]
  assign output_7_14 = io_outValid_14 & _T_4661; // @[Switch.scala 41:38:@1821.4]
  assign _T_4664 = select_15 == 4'h7; // @[Switch.scala 41:52:@1823.4]
  assign output_7_15 = io_outValid_15 & _T_4664; // @[Switch.scala 41:38:@1824.4]
  assign _T_4672 = {output_7_7,output_7_6,output_7_5,output_7_4,output_7_3,output_7_2,output_7_1,output_7_0}; // @[Switch.scala 43:31:@1832.4]
  assign _T_4680 = {output_7_15,output_7_14,output_7_13,output_7_12,output_7_11,output_7_10,output_7_9,output_7_8,_T_4672}; // @[Switch.scala 43:31:@1840.4]
  assign _T_4684 = select_0 == 4'h8; // @[Switch.scala 41:52:@1843.4]
  assign output_8_0 = io_outValid_0 & _T_4684; // @[Switch.scala 41:38:@1844.4]
  assign _T_4687 = select_1 == 4'h8; // @[Switch.scala 41:52:@1846.4]
  assign output_8_1 = io_outValid_1 & _T_4687; // @[Switch.scala 41:38:@1847.4]
  assign _T_4690 = select_2 == 4'h8; // @[Switch.scala 41:52:@1849.4]
  assign output_8_2 = io_outValid_2 & _T_4690; // @[Switch.scala 41:38:@1850.4]
  assign _T_4693 = select_3 == 4'h8; // @[Switch.scala 41:52:@1852.4]
  assign output_8_3 = io_outValid_3 & _T_4693; // @[Switch.scala 41:38:@1853.4]
  assign _T_4696 = select_4 == 4'h8; // @[Switch.scala 41:52:@1855.4]
  assign output_8_4 = io_outValid_4 & _T_4696; // @[Switch.scala 41:38:@1856.4]
  assign _T_4699 = select_5 == 4'h8; // @[Switch.scala 41:52:@1858.4]
  assign output_8_5 = io_outValid_5 & _T_4699; // @[Switch.scala 41:38:@1859.4]
  assign _T_4702 = select_6 == 4'h8; // @[Switch.scala 41:52:@1861.4]
  assign output_8_6 = io_outValid_6 & _T_4702; // @[Switch.scala 41:38:@1862.4]
  assign _T_4705 = select_7 == 4'h8; // @[Switch.scala 41:52:@1864.4]
  assign output_8_7 = io_outValid_7 & _T_4705; // @[Switch.scala 41:38:@1865.4]
  assign _T_4708 = select_8 == 4'h8; // @[Switch.scala 41:52:@1867.4]
  assign output_8_8 = io_outValid_8 & _T_4708; // @[Switch.scala 41:38:@1868.4]
  assign _T_4711 = select_9 == 4'h8; // @[Switch.scala 41:52:@1870.4]
  assign output_8_9 = io_outValid_9 & _T_4711; // @[Switch.scala 41:38:@1871.4]
  assign _T_4714 = select_10 == 4'h8; // @[Switch.scala 41:52:@1873.4]
  assign output_8_10 = io_outValid_10 & _T_4714; // @[Switch.scala 41:38:@1874.4]
  assign _T_4717 = select_11 == 4'h8; // @[Switch.scala 41:52:@1876.4]
  assign output_8_11 = io_outValid_11 & _T_4717; // @[Switch.scala 41:38:@1877.4]
  assign _T_4720 = select_12 == 4'h8; // @[Switch.scala 41:52:@1879.4]
  assign output_8_12 = io_outValid_12 & _T_4720; // @[Switch.scala 41:38:@1880.4]
  assign _T_4723 = select_13 == 4'h8; // @[Switch.scala 41:52:@1882.4]
  assign output_8_13 = io_outValid_13 & _T_4723; // @[Switch.scala 41:38:@1883.4]
  assign _T_4726 = select_14 == 4'h8; // @[Switch.scala 41:52:@1885.4]
  assign output_8_14 = io_outValid_14 & _T_4726; // @[Switch.scala 41:38:@1886.4]
  assign _T_4729 = select_15 == 4'h8; // @[Switch.scala 41:52:@1888.4]
  assign output_8_15 = io_outValid_15 & _T_4729; // @[Switch.scala 41:38:@1889.4]
  assign _T_4737 = {output_8_7,output_8_6,output_8_5,output_8_4,output_8_3,output_8_2,output_8_1,output_8_0}; // @[Switch.scala 43:31:@1897.4]
  assign _T_4745 = {output_8_15,output_8_14,output_8_13,output_8_12,output_8_11,output_8_10,output_8_9,output_8_8,_T_4737}; // @[Switch.scala 43:31:@1905.4]
  assign _T_4749 = select_0 == 4'h9; // @[Switch.scala 41:52:@1908.4]
  assign output_9_0 = io_outValid_0 & _T_4749; // @[Switch.scala 41:38:@1909.4]
  assign _T_4752 = select_1 == 4'h9; // @[Switch.scala 41:52:@1911.4]
  assign output_9_1 = io_outValid_1 & _T_4752; // @[Switch.scala 41:38:@1912.4]
  assign _T_4755 = select_2 == 4'h9; // @[Switch.scala 41:52:@1914.4]
  assign output_9_2 = io_outValid_2 & _T_4755; // @[Switch.scala 41:38:@1915.4]
  assign _T_4758 = select_3 == 4'h9; // @[Switch.scala 41:52:@1917.4]
  assign output_9_3 = io_outValid_3 & _T_4758; // @[Switch.scala 41:38:@1918.4]
  assign _T_4761 = select_4 == 4'h9; // @[Switch.scala 41:52:@1920.4]
  assign output_9_4 = io_outValid_4 & _T_4761; // @[Switch.scala 41:38:@1921.4]
  assign _T_4764 = select_5 == 4'h9; // @[Switch.scala 41:52:@1923.4]
  assign output_9_5 = io_outValid_5 & _T_4764; // @[Switch.scala 41:38:@1924.4]
  assign _T_4767 = select_6 == 4'h9; // @[Switch.scala 41:52:@1926.4]
  assign output_9_6 = io_outValid_6 & _T_4767; // @[Switch.scala 41:38:@1927.4]
  assign _T_4770 = select_7 == 4'h9; // @[Switch.scala 41:52:@1929.4]
  assign output_9_7 = io_outValid_7 & _T_4770; // @[Switch.scala 41:38:@1930.4]
  assign _T_4773 = select_8 == 4'h9; // @[Switch.scala 41:52:@1932.4]
  assign output_9_8 = io_outValid_8 & _T_4773; // @[Switch.scala 41:38:@1933.4]
  assign _T_4776 = select_9 == 4'h9; // @[Switch.scala 41:52:@1935.4]
  assign output_9_9 = io_outValid_9 & _T_4776; // @[Switch.scala 41:38:@1936.4]
  assign _T_4779 = select_10 == 4'h9; // @[Switch.scala 41:52:@1938.4]
  assign output_9_10 = io_outValid_10 & _T_4779; // @[Switch.scala 41:38:@1939.4]
  assign _T_4782 = select_11 == 4'h9; // @[Switch.scala 41:52:@1941.4]
  assign output_9_11 = io_outValid_11 & _T_4782; // @[Switch.scala 41:38:@1942.4]
  assign _T_4785 = select_12 == 4'h9; // @[Switch.scala 41:52:@1944.4]
  assign output_9_12 = io_outValid_12 & _T_4785; // @[Switch.scala 41:38:@1945.4]
  assign _T_4788 = select_13 == 4'h9; // @[Switch.scala 41:52:@1947.4]
  assign output_9_13 = io_outValid_13 & _T_4788; // @[Switch.scala 41:38:@1948.4]
  assign _T_4791 = select_14 == 4'h9; // @[Switch.scala 41:52:@1950.4]
  assign output_9_14 = io_outValid_14 & _T_4791; // @[Switch.scala 41:38:@1951.4]
  assign _T_4794 = select_15 == 4'h9; // @[Switch.scala 41:52:@1953.4]
  assign output_9_15 = io_outValid_15 & _T_4794; // @[Switch.scala 41:38:@1954.4]
  assign _T_4802 = {output_9_7,output_9_6,output_9_5,output_9_4,output_9_3,output_9_2,output_9_1,output_9_0}; // @[Switch.scala 43:31:@1962.4]
  assign _T_4810 = {output_9_15,output_9_14,output_9_13,output_9_12,output_9_11,output_9_10,output_9_9,output_9_8,_T_4802}; // @[Switch.scala 43:31:@1970.4]
  assign _T_4814 = select_0 == 4'ha; // @[Switch.scala 41:52:@1973.4]
  assign output_10_0 = io_outValid_0 & _T_4814; // @[Switch.scala 41:38:@1974.4]
  assign _T_4817 = select_1 == 4'ha; // @[Switch.scala 41:52:@1976.4]
  assign output_10_1 = io_outValid_1 & _T_4817; // @[Switch.scala 41:38:@1977.4]
  assign _T_4820 = select_2 == 4'ha; // @[Switch.scala 41:52:@1979.4]
  assign output_10_2 = io_outValid_2 & _T_4820; // @[Switch.scala 41:38:@1980.4]
  assign _T_4823 = select_3 == 4'ha; // @[Switch.scala 41:52:@1982.4]
  assign output_10_3 = io_outValid_3 & _T_4823; // @[Switch.scala 41:38:@1983.4]
  assign _T_4826 = select_4 == 4'ha; // @[Switch.scala 41:52:@1985.4]
  assign output_10_4 = io_outValid_4 & _T_4826; // @[Switch.scala 41:38:@1986.4]
  assign _T_4829 = select_5 == 4'ha; // @[Switch.scala 41:52:@1988.4]
  assign output_10_5 = io_outValid_5 & _T_4829; // @[Switch.scala 41:38:@1989.4]
  assign _T_4832 = select_6 == 4'ha; // @[Switch.scala 41:52:@1991.4]
  assign output_10_6 = io_outValid_6 & _T_4832; // @[Switch.scala 41:38:@1992.4]
  assign _T_4835 = select_7 == 4'ha; // @[Switch.scala 41:52:@1994.4]
  assign output_10_7 = io_outValid_7 & _T_4835; // @[Switch.scala 41:38:@1995.4]
  assign _T_4838 = select_8 == 4'ha; // @[Switch.scala 41:52:@1997.4]
  assign output_10_8 = io_outValid_8 & _T_4838; // @[Switch.scala 41:38:@1998.4]
  assign _T_4841 = select_9 == 4'ha; // @[Switch.scala 41:52:@2000.4]
  assign output_10_9 = io_outValid_9 & _T_4841; // @[Switch.scala 41:38:@2001.4]
  assign _T_4844 = select_10 == 4'ha; // @[Switch.scala 41:52:@2003.4]
  assign output_10_10 = io_outValid_10 & _T_4844; // @[Switch.scala 41:38:@2004.4]
  assign _T_4847 = select_11 == 4'ha; // @[Switch.scala 41:52:@2006.4]
  assign output_10_11 = io_outValid_11 & _T_4847; // @[Switch.scala 41:38:@2007.4]
  assign _T_4850 = select_12 == 4'ha; // @[Switch.scala 41:52:@2009.4]
  assign output_10_12 = io_outValid_12 & _T_4850; // @[Switch.scala 41:38:@2010.4]
  assign _T_4853 = select_13 == 4'ha; // @[Switch.scala 41:52:@2012.4]
  assign output_10_13 = io_outValid_13 & _T_4853; // @[Switch.scala 41:38:@2013.4]
  assign _T_4856 = select_14 == 4'ha; // @[Switch.scala 41:52:@2015.4]
  assign output_10_14 = io_outValid_14 & _T_4856; // @[Switch.scala 41:38:@2016.4]
  assign _T_4859 = select_15 == 4'ha; // @[Switch.scala 41:52:@2018.4]
  assign output_10_15 = io_outValid_15 & _T_4859; // @[Switch.scala 41:38:@2019.4]
  assign _T_4867 = {output_10_7,output_10_6,output_10_5,output_10_4,output_10_3,output_10_2,output_10_1,output_10_0}; // @[Switch.scala 43:31:@2027.4]
  assign _T_4875 = {output_10_15,output_10_14,output_10_13,output_10_12,output_10_11,output_10_10,output_10_9,output_10_8,_T_4867}; // @[Switch.scala 43:31:@2035.4]
  assign _T_4879 = select_0 == 4'hb; // @[Switch.scala 41:52:@2038.4]
  assign output_11_0 = io_outValid_0 & _T_4879; // @[Switch.scala 41:38:@2039.4]
  assign _T_4882 = select_1 == 4'hb; // @[Switch.scala 41:52:@2041.4]
  assign output_11_1 = io_outValid_1 & _T_4882; // @[Switch.scala 41:38:@2042.4]
  assign _T_4885 = select_2 == 4'hb; // @[Switch.scala 41:52:@2044.4]
  assign output_11_2 = io_outValid_2 & _T_4885; // @[Switch.scala 41:38:@2045.4]
  assign _T_4888 = select_3 == 4'hb; // @[Switch.scala 41:52:@2047.4]
  assign output_11_3 = io_outValid_3 & _T_4888; // @[Switch.scala 41:38:@2048.4]
  assign _T_4891 = select_4 == 4'hb; // @[Switch.scala 41:52:@2050.4]
  assign output_11_4 = io_outValid_4 & _T_4891; // @[Switch.scala 41:38:@2051.4]
  assign _T_4894 = select_5 == 4'hb; // @[Switch.scala 41:52:@2053.4]
  assign output_11_5 = io_outValid_5 & _T_4894; // @[Switch.scala 41:38:@2054.4]
  assign _T_4897 = select_6 == 4'hb; // @[Switch.scala 41:52:@2056.4]
  assign output_11_6 = io_outValid_6 & _T_4897; // @[Switch.scala 41:38:@2057.4]
  assign _T_4900 = select_7 == 4'hb; // @[Switch.scala 41:52:@2059.4]
  assign output_11_7 = io_outValid_7 & _T_4900; // @[Switch.scala 41:38:@2060.4]
  assign _T_4903 = select_8 == 4'hb; // @[Switch.scala 41:52:@2062.4]
  assign output_11_8 = io_outValid_8 & _T_4903; // @[Switch.scala 41:38:@2063.4]
  assign _T_4906 = select_9 == 4'hb; // @[Switch.scala 41:52:@2065.4]
  assign output_11_9 = io_outValid_9 & _T_4906; // @[Switch.scala 41:38:@2066.4]
  assign _T_4909 = select_10 == 4'hb; // @[Switch.scala 41:52:@2068.4]
  assign output_11_10 = io_outValid_10 & _T_4909; // @[Switch.scala 41:38:@2069.4]
  assign _T_4912 = select_11 == 4'hb; // @[Switch.scala 41:52:@2071.4]
  assign output_11_11 = io_outValid_11 & _T_4912; // @[Switch.scala 41:38:@2072.4]
  assign _T_4915 = select_12 == 4'hb; // @[Switch.scala 41:52:@2074.4]
  assign output_11_12 = io_outValid_12 & _T_4915; // @[Switch.scala 41:38:@2075.4]
  assign _T_4918 = select_13 == 4'hb; // @[Switch.scala 41:52:@2077.4]
  assign output_11_13 = io_outValid_13 & _T_4918; // @[Switch.scala 41:38:@2078.4]
  assign _T_4921 = select_14 == 4'hb; // @[Switch.scala 41:52:@2080.4]
  assign output_11_14 = io_outValid_14 & _T_4921; // @[Switch.scala 41:38:@2081.4]
  assign _T_4924 = select_15 == 4'hb; // @[Switch.scala 41:52:@2083.4]
  assign output_11_15 = io_outValid_15 & _T_4924; // @[Switch.scala 41:38:@2084.4]
  assign _T_4932 = {output_11_7,output_11_6,output_11_5,output_11_4,output_11_3,output_11_2,output_11_1,output_11_0}; // @[Switch.scala 43:31:@2092.4]
  assign _T_4940 = {output_11_15,output_11_14,output_11_13,output_11_12,output_11_11,output_11_10,output_11_9,output_11_8,_T_4932}; // @[Switch.scala 43:31:@2100.4]
  assign _T_4944 = select_0 == 4'hc; // @[Switch.scala 41:52:@2103.4]
  assign output_12_0 = io_outValid_0 & _T_4944; // @[Switch.scala 41:38:@2104.4]
  assign _T_4947 = select_1 == 4'hc; // @[Switch.scala 41:52:@2106.4]
  assign output_12_1 = io_outValid_1 & _T_4947; // @[Switch.scala 41:38:@2107.4]
  assign _T_4950 = select_2 == 4'hc; // @[Switch.scala 41:52:@2109.4]
  assign output_12_2 = io_outValid_2 & _T_4950; // @[Switch.scala 41:38:@2110.4]
  assign _T_4953 = select_3 == 4'hc; // @[Switch.scala 41:52:@2112.4]
  assign output_12_3 = io_outValid_3 & _T_4953; // @[Switch.scala 41:38:@2113.4]
  assign _T_4956 = select_4 == 4'hc; // @[Switch.scala 41:52:@2115.4]
  assign output_12_4 = io_outValid_4 & _T_4956; // @[Switch.scala 41:38:@2116.4]
  assign _T_4959 = select_5 == 4'hc; // @[Switch.scala 41:52:@2118.4]
  assign output_12_5 = io_outValid_5 & _T_4959; // @[Switch.scala 41:38:@2119.4]
  assign _T_4962 = select_6 == 4'hc; // @[Switch.scala 41:52:@2121.4]
  assign output_12_6 = io_outValid_6 & _T_4962; // @[Switch.scala 41:38:@2122.4]
  assign _T_4965 = select_7 == 4'hc; // @[Switch.scala 41:52:@2124.4]
  assign output_12_7 = io_outValid_7 & _T_4965; // @[Switch.scala 41:38:@2125.4]
  assign _T_4968 = select_8 == 4'hc; // @[Switch.scala 41:52:@2127.4]
  assign output_12_8 = io_outValid_8 & _T_4968; // @[Switch.scala 41:38:@2128.4]
  assign _T_4971 = select_9 == 4'hc; // @[Switch.scala 41:52:@2130.4]
  assign output_12_9 = io_outValid_9 & _T_4971; // @[Switch.scala 41:38:@2131.4]
  assign _T_4974 = select_10 == 4'hc; // @[Switch.scala 41:52:@2133.4]
  assign output_12_10 = io_outValid_10 & _T_4974; // @[Switch.scala 41:38:@2134.4]
  assign _T_4977 = select_11 == 4'hc; // @[Switch.scala 41:52:@2136.4]
  assign output_12_11 = io_outValid_11 & _T_4977; // @[Switch.scala 41:38:@2137.4]
  assign _T_4980 = select_12 == 4'hc; // @[Switch.scala 41:52:@2139.4]
  assign output_12_12 = io_outValid_12 & _T_4980; // @[Switch.scala 41:38:@2140.4]
  assign _T_4983 = select_13 == 4'hc; // @[Switch.scala 41:52:@2142.4]
  assign output_12_13 = io_outValid_13 & _T_4983; // @[Switch.scala 41:38:@2143.4]
  assign _T_4986 = select_14 == 4'hc; // @[Switch.scala 41:52:@2145.4]
  assign output_12_14 = io_outValid_14 & _T_4986; // @[Switch.scala 41:38:@2146.4]
  assign _T_4989 = select_15 == 4'hc; // @[Switch.scala 41:52:@2148.4]
  assign output_12_15 = io_outValid_15 & _T_4989; // @[Switch.scala 41:38:@2149.4]
  assign _T_4997 = {output_12_7,output_12_6,output_12_5,output_12_4,output_12_3,output_12_2,output_12_1,output_12_0}; // @[Switch.scala 43:31:@2157.4]
  assign _T_5005 = {output_12_15,output_12_14,output_12_13,output_12_12,output_12_11,output_12_10,output_12_9,output_12_8,_T_4997}; // @[Switch.scala 43:31:@2165.4]
  assign _T_5009 = select_0 == 4'hd; // @[Switch.scala 41:52:@2168.4]
  assign output_13_0 = io_outValid_0 & _T_5009; // @[Switch.scala 41:38:@2169.4]
  assign _T_5012 = select_1 == 4'hd; // @[Switch.scala 41:52:@2171.4]
  assign output_13_1 = io_outValid_1 & _T_5012; // @[Switch.scala 41:38:@2172.4]
  assign _T_5015 = select_2 == 4'hd; // @[Switch.scala 41:52:@2174.4]
  assign output_13_2 = io_outValid_2 & _T_5015; // @[Switch.scala 41:38:@2175.4]
  assign _T_5018 = select_3 == 4'hd; // @[Switch.scala 41:52:@2177.4]
  assign output_13_3 = io_outValid_3 & _T_5018; // @[Switch.scala 41:38:@2178.4]
  assign _T_5021 = select_4 == 4'hd; // @[Switch.scala 41:52:@2180.4]
  assign output_13_4 = io_outValid_4 & _T_5021; // @[Switch.scala 41:38:@2181.4]
  assign _T_5024 = select_5 == 4'hd; // @[Switch.scala 41:52:@2183.4]
  assign output_13_5 = io_outValid_5 & _T_5024; // @[Switch.scala 41:38:@2184.4]
  assign _T_5027 = select_6 == 4'hd; // @[Switch.scala 41:52:@2186.4]
  assign output_13_6 = io_outValid_6 & _T_5027; // @[Switch.scala 41:38:@2187.4]
  assign _T_5030 = select_7 == 4'hd; // @[Switch.scala 41:52:@2189.4]
  assign output_13_7 = io_outValid_7 & _T_5030; // @[Switch.scala 41:38:@2190.4]
  assign _T_5033 = select_8 == 4'hd; // @[Switch.scala 41:52:@2192.4]
  assign output_13_8 = io_outValid_8 & _T_5033; // @[Switch.scala 41:38:@2193.4]
  assign _T_5036 = select_9 == 4'hd; // @[Switch.scala 41:52:@2195.4]
  assign output_13_9 = io_outValid_9 & _T_5036; // @[Switch.scala 41:38:@2196.4]
  assign _T_5039 = select_10 == 4'hd; // @[Switch.scala 41:52:@2198.4]
  assign output_13_10 = io_outValid_10 & _T_5039; // @[Switch.scala 41:38:@2199.4]
  assign _T_5042 = select_11 == 4'hd; // @[Switch.scala 41:52:@2201.4]
  assign output_13_11 = io_outValid_11 & _T_5042; // @[Switch.scala 41:38:@2202.4]
  assign _T_5045 = select_12 == 4'hd; // @[Switch.scala 41:52:@2204.4]
  assign output_13_12 = io_outValid_12 & _T_5045; // @[Switch.scala 41:38:@2205.4]
  assign _T_5048 = select_13 == 4'hd; // @[Switch.scala 41:52:@2207.4]
  assign output_13_13 = io_outValid_13 & _T_5048; // @[Switch.scala 41:38:@2208.4]
  assign _T_5051 = select_14 == 4'hd; // @[Switch.scala 41:52:@2210.4]
  assign output_13_14 = io_outValid_14 & _T_5051; // @[Switch.scala 41:38:@2211.4]
  assign _T_5054 = select_15 == 4'hd; // @[Switch.scala 41:52:@2213.4]
  assign output_13_15 = io_outValid_15 & _T_5054; // @[Switch.scala 41:38:@2214.4]
  assign _T_5062 = {output_13_7,output_13_6,output_13_5,output_13_4,output_13_3,output_13_2,output_13_1,output_13_0}; // @[Switch.scala 43:31:@2222.4]
  assign _T_5070 = {output_13_15,output_13_14,output_13_13,output_13_12,output_13_11,output_13_10,output_13_9,output_13_8,_T_5062}; // @[Switch.scala 43:31:@2230.4]
  assign _T_5074 = select_0 == 4'he; // @[Switch.scala 41:52:@2233.4]
  assign output_14_0 = io_outValid_0 & _T_5074; // @[Switch.scala 41:38:@2234.4]
  assign _T_5077 = select_1 == 4'he; // @[Switch.scala 41:52:@2236.4]
  assign output_14_1 = io_outValid_1 & _T_5077; // @[Switch.scala 41:38:@2237.4]
  assign _T_5080 = select_2 == 4'he; // @[Switch.scala 41:52:@2239.4]
  assign output_14_2 = io_outValid_2 & _T_5080; // @[Switch.scala 41:38:@2240.4]
  assign _T_5083 = select_3 == 4'he; // @[Switch.scala 41:52:@2242.4]
  assign output_14_3 = io_outValid_3 & _T_5083; // @[Switch.scala 41:38:@2243.4]
  assign _T_5086 = select_4 == 4'he; // @[Switch.scala 41:52:@2245.4]
  assign output_14_4 = io_outValid_4 & _T_5086; // @[Switch.scala 41:38:@2246.4]
  assign _T_5089 = select_5 == 4'he; // @[Switch.scala 41:52:@2248.4]
  assign output_14_5 = io_outValid_5 & _T_5089; // @[Switch.scala 41:38:@2249.4]
  assign _T_5092 = select_6 == 4'he; // @[Switch.scala 41:52:@2251.4]
  assign output_14_6 = io_outValid_6 & _T_5092; // @[Switch.scala 41:38:@2252.4]
  assign _T_5095 = select_7 == 4'he; // @[Switch.scala 41:52:@2254.4]
  assign output_14_7 = io_outValid_7 & _T_5095; // @[Switch.scala 41:38:@2255.4]
  assign _T_5098 = select_8 == 4'he; // @[Switch.scala 41:52:@2257.4]
  assign output_14_8 = io_outValid_8 & _T_5098; // @[Switch.scala 41:38:@2258.4]
  assign _T_5101 = select_9 == 4'he; // @[Switch.scala 41:52:@2260.4]
  assign output_14_9 = io_outValid_9 & _T_5101; // @[Switch.scala 41:38:@2261.4]
  assign _T_5104 = select_10 == 4'he; // @[Switch.scala 41:52:@2263.4]
  assign output_14_10 = io_outValid_10 & _T_5104; // @[Switch.scala 41:38:@2264.4]
  assign _T_5107 = select_11 == 4'he; // @[Switch.scala 41:52:@2266.4]
  assign output_14_11 = io_outValid_11 & _T_5107; // @[Switch.scala 41:38:@2267.4]
  assign _T_5110 = select_12 == 4'he; // @[Switch.scala 41:52:@2269.4]
  assign output_14_12 = io_outValid_12 & _T_5110; // @[Switch.scala 41:38:@2270.4]
  assign _T_5113 = select_13 == 4'he; // @[Switch.scala 41:52:@2272.4]
  assign output_14_13 = io_outValid_13 & _T_5113; // @[Switch.scala 41:38:@2273.4]
  assign _T_5116 = select_14 == 4'he; // @[Switch.scala 41:52:@2275.4]
  assign output_14_14 = io_outValid_14 & _T_5116; // @[Switch.scala 41:38:@2276.4]
  assign _T_5119 = select_15 == 4'he; // @[Switch.scala 41:52:@2278.4]
  assign output_14_15 = io_outValid_15 & _T_5119; // @[Switch.scala 41:38:@2279.4]
  assign _T_5127 = {output_14_7,output_14_6,output_14_5,output_14_4,output_14_3,output_14_2,output_14_1,output_14_0}; // @[Switch.scala 43:31:@2287.4]
  assign _T_5135 = {output_14_15,output_14_14,output_14_13,output_14_12,output_14_11,output_14_10,output_14_9,output_14_8,_T_5127}; // @[Switch.scala 43:31:@2295.4]
  assign _T_5139 = select_0 == 4'hf; // @[Switch.scala 41:52:@2298.4]
  assign output_15_0 = io_outValid_0 & _T_5139; // @[Switch.scala 41:38:@2299.4]
  assign _T_5142 = select_1 == 4'hf; // @[Switch.scala 41:52:@2301.4]
  assign output_15_1 = io_outValid_1 & _T_5142; // @[Switch.scala 41:38:@2302.4]
  assign _T_5145 = select_2 == 4'hf; // @[Switch.scala 41:52:@2304.4]
  assign output_15_2 = io_outValid_2 & _T_5145; // @[Switch.scala 41:38:@2305.4]
  assign _T_5148 = select_3 == 4'hf; // @[Switch.scala 41:52:@2307.4]
  assign output_15_3 = io_outValid_3 & _T_5148; // @[Switch.scala 41:38:@2308.4]
  assign _T_5151 = select_4 == 4'hf; // @[Switch.scala 41:52:@2310.4]
  assign output_15_4 = io_outValid_4 & _T_5151; // @[Switch.scala 41:38:@2311.4]
  assign _T_5154 = select_5 == 4'hf; // @[Switch.scala 41:52:@2313.4]
  assign output_15_5 = io_outValid_5 & _T_5154; // @[Switch.scala 41:38:@2314.4]
  assign _T_5157 = select_6 == 4'hf; // @[Switch.scala 41:52:@2316.4]
  assign output_15_6 = io_outValid_6 & _T_5157; // @[Switch.scala 41:38:@2317.4]
  assign _T_5160 = select_7 == 4'hf; // @[Switch.scala 41:52:@2319.4]
  assign output_15_7 = io_outValid_7 & _T_5160; // @[Switch.scala 41:38:@2320.4]
  assign _T_5163 = select_8 == 4'hf; // @[Switch.scala 41:52:@2322.4]
  assign output_15_8 = io_outValid_8 & _T_5163; // @[Switch.scala 41:38:@2323.4]
  assign _T_5166 = select_9 == 4'hf; // @[Switch.scala 41:52:@2325.4]
  assign output_15_9 = io_outValid_9 & _T_5166; // @[Switch.scala 41:38:@2326.4]
  assign _T_5169 = select_10 == 4'hf; // @[Switch.scala 41:52:@2328.4]
  assign output_15_10 = io_outValid_10 & _T_5169; // @[Switch.scala 41:38:@2329.4]
  assign _T_5172 = select_11 == 4'hf; // @[Switch.scala 41:52:@2331.4]
  assign output_15_11 = io_outValid_11 & _T_5172; // @[Switch.scala 41:38:@2332.4]
  assign _T_5175 = select_12 == 4'hf; // @[Switch.scala 41:52:@2334.4]
  assign output_15_12 = io_outValid_12 & _T_5175; // @[Switch.scala 41:38:@2335.4]
  assign _T_5178 = select_13 == 4'hf; // @[Switch.scala 41:52:@2337.4]
  assign output_15_13 = io_outValid_13 & _T_5178; // @[Switch.scala 41:38:@2338.4]
  assign _T_5181 = select_14 == 4'hf; // @[Switch.scala 41:52:@2340.4]
  assign output_15_14 = io_outValid_14 & _T_5181; // @[Switch.scala 41:38:@2341.4]
  assign _T_5184 = select_15 == 4'hf; // @[Switch.scala 41:52:@2343.4]
  assign output_15_15 = io_outValid_15 & _T_5184; // @[Switch.scala 41:38:@2344.4]
  assign _T_5192 = {output_15_7,output_15_6,output_15_5,output_15_4,output_15_3,output_15_2,output_15_1,output_15_0}; // @[Switch.scala 43:31:@2352.4]
  assign _T_5200 = {output_15_15,output_15_14,output_15_13,output_15_12,output_15_11,output_15_10,output_15_9,output_15_8,_T_5192}; // @[Switch.scala 43:31:@2360.4]
  assign io_outAck_0 = _T_4225 != 16'h0; // @[Switch.scala 43:18:@1387.4]
  assign io_outAck_1 = _T_4290 != 16'h0; // @[Switch.scala 43:18:@1452.4]
  assign io_outAck_2 = _T_4355 != 16'h0; // @[Switch.scala 43:18:@1517.4]
  assign io_outAck_3 = _T_4420 != 16'h0; // @[Switch.scala 43:18:@1582.4]
  assign io_outAck_4 = _T_4485 != 16'h0; // @[Switch.scala 43:18:@1647.4]
  assign io_outAck_5 = _T_4550 != 16'h0; // @[Switch.scala 43:18:@1712.4]
  assign io_outAck_6 = _T_4615 != 16'h0; // @[Switch.scala 43:18:@1777.4]
  assign io_outAck_7 = _T_4680 != 16'h0; // @[Switch.scala 43:18:@1842.4]
  assign io_outAck_8 = _T_4745 != 16'h0; // @[Switch.scala 43:18:@1907.4]
  assign io_outAck_9 = _T_4810 != 16'h0; // @[Switch.scala 43:18:@1972.4]
  assign io_outAck_10 = _T_4875 != 16'h0; // @[Switch.scala 43:18:@2037.4]
  assign io_outAck_11 = _T_4940 != 16'h0; // @[Switch.scala 43:18:@2102.4]
  assign io_outAck_12 = _T_5005 != 16'h0; // @[Switch.scala 43:18:@2167.4]
  assign io_outAck_13 = _T_5070 != 16'h0; // @[Switch.scala 43:18:@2232.4]
  assign io_outAck_14 = _T_5135 != 16'h0; // @[Switch.scala 43:18:@2297.4]
  assign io_outAck_15 = _T_5200 != 16'h0; // @[Switch.scala 43:18:@2362.4]
  assign io_outData_0 = 4'hf == select_0 ? io_inData_15 : _GEN_14; // @[Switch.scala 33:19:@74.4]
  assign io_outData_1 = 4'hf == select_1 ? io_inData_15 : _GEN_30; // @[Switch.scala 33:19:@156.4]
  assign io_outData_2 = 4'hf == select_2 ? io_inData_15 : _GEN_46; // @[Switch.scala 33:19:@238.4]
  assign io_outData_3 = 4'hf == select_3 ? io_inData_15 : _GEN_62; // @[Switch.scala 33:19:@320.4]
  assign io_outData_4 = 4'hf == select_4 ? io_inData_15 : _GEN_78; // @[Switch.scala 33:19:@402.4]
  assign io_outData_5 = 4'hf == select_5 ? io_inData_15 : _GEN_94; // @[Switch.scala 33:19:@484.4]
  assign io_outData_6 = 4'hf == select_6 ? io_inData_15 : _GEN_110; // @[Switch.scala 33:19:@566.4]
  assign io_outData_7 = 4'hf == select_7 ? io_inData_15 : _GEN_126; // @[Switch.scala 33:19:@648.4]
  assign io_outData_8 = 4'hf == select_8 ? io_inData_15 : _GEN_142; // @[Switch.scala 33:19:@730.4]
  assign io_outData_9 = 4'hf == select_9 ? io_inData_15 : _GEN_158; // @[Switch.scala 33:19:@812.4]
  assign io_outData_10 = 4'hf == select_10 ? io_inData_15 : _GEN_174; // @[Switch.scala 33:19:@894.4]
  assign io_outData_11 = 4'hf == select_11 ? io_inData_15 : _GEN_190; // @[Switch.scala 33:19:@976.4]
  assign io_outData_12 = 4'hf == select_12 ? io_inData_15 : _GEN_206; // @[Switch.scala 33:19:@1058.4]
  assign io_outData_13 = 4'hf == select_13 ? io_inData_15 : _GEN_222; // @[Switch.scala 33:19:@1140.4]
  assign io_outData_14 = 4'hf == select_14 ? io_inData_15 : _GEN_238; // @[Switch.scala 33:19:@1222.4]
  assign io_outData_15 = 4'hf == select_15 ? io_inData_15 : _GEN_254; // @[Switch.scala 33:19:@1304.4]
  assign io_outValid_0 = _T_1475 != 16'h0; // @[Switch.scala 34:20:@91.4]
  assign io_outValid_1 = _T_1572 != 16'h0; // @[Switch.scala 34:20:@173.4]
  assign io_outValid_2 = _T_1669 != 16'h0; // @[Switch.scala 34:20:@255.4]
  assign io_outValid_3 = _T_1766 != 16'h0; // @[Switch.scala 34:20:@337.4]
  assign io_outValid_4 = _T_1863 != 16'h0; // @[Switch.scala 34:20:@419.4]
  assign io_outValid_5 = _T_1960 != 16'h0; // @[Switch.scala 34:20:@501.4]
  assign io_outValid_6 = _T_2057 != 16'h0; // @[Switch.scala 34:20:@583.4]
  assign io_outValid_7 = _T_2154 != 16'h0; // @[Switch.scala 34:20:@665.4]
  assign io_outValid_8 = _T_2251 != 16'h0; // @[Switch.scala 34:20:@747.4]
  assign io_outValid_9 = _T_2348 != 16'h0; // @[Switch.scala 34:20:@829.4]
  assign io_outValid_10 = _T_2445 != 16'h0; // @[Switch.scala 34:20:@911.4]
  assign io_outValid_11 = _T_2542 != 16'h0; // @[Switch.scala 34:20:@993.4]
  assign io_outValid_12 = _T_2639 != 16'h0; // @[Switch.scala 34:20:@1075.4]
  assign io_outValid_13 = _T_2736 != 16'h0; // @[Switch.scala 34:20:@1157.4]
  assign io_outValid_14 = _T_2833 != 16'h0; // @[Switch.scala 34:20:@1239.4]
  assign io_outValid_15 = _T_2930 != 16'h0; // @[Switch.scala 34:20:@1321.4]
endmodule
module SwitchWrapper( // @[:@2364.2]
  input         clock, // @[:@2365.4]
  input         reset, // @[:@2366.4]
  input  [3:0]  io_inAddr_0, // @[:@2367.4]
  input  [3:0]  io_inAddr_1, // @[:@2367.4]
  input  [3:0]  io_inAddr_2, // @[:@2367.4]
  input  [3:0]  io_inAddr_3, // @[:@2367.4]
  input  [3:0]  io_inAddr_4, // @[:@2367.4]
  input  [3:0]  io_inAddr_5, // @[:@2367.4]
  input  [3:0]  io_inAddr_6, // @[:@2367.4]
  input  [3:0]  io_inAddr_7, // @[:@2367.4]
  input  [3:0]  io_inAddr_8, // @[:@2367.4]
  input  [3:0]  io_inAddr_9, // @[:@2367.4]
  input  [3:0]  io_inAddr_10, // @[:@2367.4]
  input  [3:0]  io_inAddr_11, // @[:@2367.4]
  input  [3:0]  io_inAddr_12, // @[:@2367.4]
  input  [3:0]  io_inAddr_13, // @[:@2367.4]
  input  [3:0]  io_inAddr_14, // @[:@2367.4]
  input  [3:0]  io_inAddr_15, // @[:@2367.4]
  input  [47:0] io_inData_0, // @[:@2367.4]
  input  [47:0] io_inData_1, // @[:@2367.4]
  input  [47:0] io_inData_2, // @[:@2367.4]
  input  [47:0] io_inData_3, // @[:@2367.4]
  input  [47:0] io_inData_4, // @[:@2367.4]
  input  [47:0] io_inData_5, // @[:@2367.4]
  input  [47:0] io_inData_6, // @[:@2367.4]
  input  [47:0] io_inData_7, // @[:@2367.4]
  input  [47:0] io_inData_8, // @[:@2367.4]
  input  [47:0] io_inData_9, // @[:@2367.4]
  input  [47:0] io_inData_10, // @[:@2367.4]
  input  [47:0] io_inData_11, // @[:@2367.4]
  input  [47:0] io_inData_12, // @[:@2367.4]
  input  [47:0] io_inData_13, // @[:@2367.4]
  input  [47:0] io_inData_14, // @[:@2367.4]
  input  [47:0] io_inData_15, // @[:@2367.4]
  input         io_inValid_0, // @[:@2367.4]
  input         io_inValid_1, // @[:@2367.4]
  input         io_inValid_2, // @[:@2367.4]
  input         io_inValid_3, // @[:@2367.4]
  input         io_inValid_4, // @[:@2367.4]
  input         io_inValid_5, // @[:@2367.4]
  input         io_inValid_6, // @[:@2367.4]
  input         io_inValid_7, // @[:@2367.4]
  input         io_inValid_8, // @[:@2367.4]
  input         io_inValid_9, // @[:@2367.4]
  input         io_inValid_10, // @[:@2367.4]
  input         io_inValid_11, // @[:@2367.4]
  input         io_inValid_12, // @[:@2367.4]
  input         io_inValid_13, // @[:@2367.4]
  input         io_inValid_14, // @[:@2367.4]
  input         io_inValid_15, // @[:@2367.4]
  output        io_outAck_0, // @[:@2367.4]
  output        io_outAck_1, // @[:@2367.4]
  output        io_outAck_2, // @[:@2367.4]
  output        io_outAck_3, // @[:@2367.4]
  output        io_outAck_4, // @[:@2367.4]
  output        io_outAck_5, // @[:@2367.4]
  output        io_outAck_6, // @[:@2367.4]
  output        io_outAck_7, // @[:@2367.4]
  output        io_outAck_8, // @[:@2367.4]
  output        io_outAck_9, // @[:@2367.4]
  output        io_outAck_10, // @[:@2367.4]
  output        io_outAck_11, // @[:@2367.4]
  output        io_outAck_12, // @[:@2367.4]
  output        io_outAck_13, // @[:@2367.4]
  output        io_outAck_14, // @[:@2367.4]
  output        io_outAck_15, // @[:@2367.4]
  output [47:0] io_outData_0, // @[:@2367.4]
  output [47:0] io_outData_1, // @[:@2367.4]
  output [47:0] io_outData_2, // @[:@2367.4]
  output [47:0] io_outData_3, // @[:@2367.4]
  output [47:0] io_outData_4, // @[:@2367.4]
  output [47:0] io_outData_5, // @[:@2367.4]
  output [47:0] io_outData_6, // @[:@2367.4]
  output [47:0] io_outData_7, // @[:@2367.4]
  output [47:0] io_outData_8, // @[:@2367.4]
  output [47:0] io_outData_9, // @[:@2367.4]
  output [47:0] io_outData_10, // @[:@2367.4]
  output [47:0] io_outData_11, // @[:@2367.4]
  output [47:0] io_outData_12, // @[:@2367.4]
  output [47:0] io_outData_13, // @[:@2367.4]
  output [47:0] io_outData_14, // @[:@2367.4]
  output [47:0] io_outData_15, // @[:@2367.4]
  output        io_outValid_0, // @[:@2367.4]
  output        io_outValid_1, // @[:@2367.4]
  output        io_outValid_2, // @[:@2367.4]
  output        io_outValid_3, // @[:@2367.4]
  output        io_outValid_4, // @[:@2367.4]
  output        io_outValid_5, // @[:@2367.4]
  output        io_outValid_6, // @[:@2367.4]
  output        io_outValid_7, // @[:@2367.4]
  output        io_outValid_8, // @[:@2367.4]
  output        io_outValid_9, // @[:@2367.4]
  output        io_outValid_10, // @[:@2367.4]
  output        io_outValid_11, // @[:@2367.4]
  output        io_outValid_12, // @[:@2367.4]
  output        io_outValid_13, // @[:@2367.4]
  output        io_outValid_14, // @[:@2367.4]
  output        io_outValid_15 // @[:@2367.4]
);
  wire [3:0] switch_io_inAddr_0; // @[Switch.scala 50:22:@2369.4]
  wire [3:0] switch_io_inAddr_1; // @[Switch.scala 50:22:@2369.4]
  wire [3:0] switch_io_inAddr_2; // @[Switch.scala 50:22:@2369.4]
  wire [3:0] switch_io_inAddr_3; // @[Switch.scala 50:22:@2369.4]
  wire [3:0] switch_io_inAddr_4; // @[Switch.scala 50:22:@2369.4]
  wire [3:0] switch_io_inAddr_5; // @[Switch.scala 50:22:@2369.4]
  wire [3:0] switch_io_inAddr_6; // @[Switch.scala 50:22:@2369.4]
  wire [3:0] switch_io_inAddr_7; // @[Switch.scala 50:22:@2369.4]
  wire [3:0] switch_io_inAddr_8; // @[Switch.scala 50:22:@2369.4]
  wire [3:0] switch_io_inAddr_9; // @[Switch.scala 50:22:@2369.4]
  wire [3:0] switch_io_inAddr_10; // @[Switch.scala 50:22:@2369.4]
  wire [3:0] switch_io_inAddr_11; // @[Switch.scala 50:22:@2369.4]
  wire [3:0] switch_io_inAddr_12; // @[Switch.scala 50:22:@2369.4]
  wire [3:0] switch_io_inAddr_13; // @[Switch.scala 50:22:@2369.4]
  wire [3:0] switch_io_inAddr_14; // @[Switch.scala 50:22:@2369.4]
  wire [3:0] switch_io_inAddr_15; // @[Switch.scala 50:22:@2369.4]
  wire [47:0] switch_io_inData_0; // @[Switch.scala 50:22:@2369.4]
  wire [47:0] switch_io_inData_1; // @[Switch.scala 50:22:@2369.4]
  wire [47:0] switch_io_inData_2; // @[Switch.scala 50:22:@2369.4]
  wire [47:0] switch_io_inData_3; // @[Switch.scala 50:22:@2369.4]
  wire [47:0] switch_io_inData_4; // @[Switch.scala 50:22:@2369.4]
  wire [47:0] switch_io_inData_5; // @[Switch.scala 50:22:@2369.4]
  wire [47:0] switch_io_inData_6; // @[Switch.scala 50:22:@2369.4]
  wire [47:0] switch_io_inData_7; // @[Switch.scala 50:22:@2369.4]
  wire [47:0] switch_io_inData_8; // @[Switch.scala 50:22:@2369.4]
  wire [47:0] switch_io_inData_9; // @[Switch.scala 50:22:@2369.4]
  wire [47:0] switch_io_inData_10; // @[Switch.scala 50:22:@2369.4]
  wire [47:0] switch_io_inData_11; // @[Switch.scala 50:22:@2369.4]
  wire [47:0] switch_io_inData_12; // @[Switch.scala 50:22:@2369.4]
  wire [47:0] switch_io_inData_13; // @[Switch.scala 50:22:@2369.4]
  wire [47:0] switch_io_inData_14; // @[Switch.scala 50:22:@2369.4]
  wire [47:0] switch_io_inData_15; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_inValid_0; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_inValid_1; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_inValid_2; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_inValid_3; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_inValid_4; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_inValid_5; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_inValid_6; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_inValid_7; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_inValid_8; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_inValid_9; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_inValid_10; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_inValid_11; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_inValid_12; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_inValid_13; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_inValid_14; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_inValid_15; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_outAck_0; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_outAck_1; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_outAck_2; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_outAck_3; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_outAck_4; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_outAck_5; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_outAck_6; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_outAck_7; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_outAck_8; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_outAck_9; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_outAck_10; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_outAck_11; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_outAck_12; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_outAck_13; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_outAck_14; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_outAck_15; // @[Switch.scala 50:22:@2369.4]
  wire [47:0] switch_io_outData_0; // @[Switch.scala 50:22:@2369.4]
  wire [47:0] switch_io_outData_1; // @[Switch.scala 50:22:@2369.4]
  wire [47:0] switch_io_outData_2; // @[Switch.scala 50:22:@2369.4]
  wire [47:0] switch_io_outData_3; // @[Switch.scala 50:22:@2369.4]
  wire [47:0] switch_io_outData_4; // @[Switch.scala 50:22:@2369.4]
  wire [47:0] switch_io_outData_5; // @[Switch.scala 50:22:@2369.4]
  wire [47:0] switch_io_outData_6; // @[Switch.scala 50:22:@2369.4]
  wire [47:0] switch_io_outData_7; // @[Switch.scala 50:22:@2369.4]
  wire [47:0] switch_io_outData_8; // @[Switch.scala 50:22:@2369.4]
  wire [47:0] switch_io_outData_9; // @[Switch.scala 50:22:@2369.4]
  wire [47:0] switch_io_outData_10; // @[Switch.scala 50:22:@2369.4]
  wire [47:0] switch_io_outData_11; // @[Switch.scala 50:22:@2369.4]
  wire [47:0] switch_io_outData_12; // @[Switch.scala 50:22:@2369.4]
  wire [47:0] switch_io_outData_13; // @[Switch.scala 50:22:@2369.4]
  wire [47:0] switch_io_outData_14; // @[Switch.scala 50:22:@2369.4]
  wire [47:0] switch_io_outData_15; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_outValid_0; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_outValid_1; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_outValid_2; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_outValid_3; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_outValid_4; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_outValid_5; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_outValid_6; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_outValid_7; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_outValid_8; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_outValid_9; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_outValid_10; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_outValid_11; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_outValid_12; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_outValid_13; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_outValid_14; // @[Switch.scala 50:22:@2369.4]
  wire  switch_io_outValid_15; // @[Switch.scala 50:22:@2369.4]
  reg [3:0] _T_166_0; // @[Switch.scala 51:30:@2372.4]
  reg [31:0] _RAND_0;
  reg [3:0] _T_166_1; // @[Switch.scala 51:30:@2372.4]
  reg [31:0] _RAND_1;
  reg [3:0] _T_166_2; // @[Switch.scala 51:30:@2372.4]
  reg [31:0] _RAND_2;
  reg [3:0] _T_166_3; // @[Switch.scala 51:30:@2372.4]
  reg [31:0] _RAND_3;
  reg [3:0] _T_166_4; // @[Switch.scala 51:30:@2372.4]
  reg [31:0] _RAND_4;
  reg [3:0] _T_166_5; // @[Switch.scala 51:30:@2372.4]
  reg [31:0] _RAND_5;
  reg [3:0] _T_166_6; // @[Switch.scala 51:30:@2372.4]
  reg [31:0] _RAND_6;
  reg [3:0] _T_166_7; // @[Switch.scala 51:30:@2372.4]
  reg [31:0] _RAND_7;
  reg [3:0] _T_166_8; // @[Switch.scala 51:30:@2372.4]
  reg [31:0] _RAND_8;
  reg [3:0] _T_166_9; // @[Switch.scala 51:30:@2372.4]
  reg [31:0] _RAND_9;
  reg [3:0] _T_166_10; // @[Switch.scala 51:30:@2372.4]
  reg [31:0] _RAND_10;
  reg [3:0] _T_166_11; // @[Switch.scala 51:30:@2372.4]
  reg [31:0] _RAND_11;
  reg [3:0] _T_166_12; // @[Switch.scala 51:30:@2372.4]
  reg [31:0] _RAND_12;
  reg [3:0] _T_166_13; // @[Switch.scala 51:30:@2372.4]
  reg [31:0] _RAND_13;
  reg [3:0] _T_166_14; // @[Switch.scala 51:30:@2372.4]
  reg [31:0] _RAND_14;
  reg [3:0] _T_166_15; // @[Switch.scala 51:30:@2372.4]
  reg [31:0] _RAND_15;
  reg [47:0] _T_255_0; // @[Switch.scala 52:30:@2405.4]
  reg [63:0] _RAND_16;
  reg [47:0] _T_255_1; // @[Switch.scala 52:30:@2405.4]
  reg [63:0] _RAND_17;
  reg [47:0] _T_255_2; // @[Switch.scala 52:30:@2405.4]
  reg [63:0] _RAND_18;
  reg [47:0] _T_255_3; // @[Switch.scala 52:30:@2405.4]
  reg [63:0] _RAND_19;
  reg [47:0] _T_255_4; // @[Switch.scala 52:30:@2405.4]
  reg [63:0] _RAND_20;
  reg [47:0] _T_255_5; // @[Switch.scala 52:30:@2405.4]
  reg [63:0] _RAND_21;
  reg [47:0] _T_255_6; // @[Switch.scala 52:30:@2405.4]
  reg [63:0] _RAND_22;
  reg [47:0] _T_255_7; // @[Switch.scala 52:30:@2405.4]
  reg [63:0] _RAND_23;
  reg [47:0] _T_255_8; // @[Switch.scala 52:30:@2405.4]
  reg [63:0] _RAND_24;
  reg [47:0] _T_255_9; // @[Switch.scala 52:30:@2405.4]
  reg [63:0] _RAND_25;
  reg [47:0] _T_255_10; // @[Switch.scala 52:30:@2405.4]
  reg [63:0] _RAND_26;
  reg [47:0] _T_255_11; // @[Switch.scala 52:30:@2405.4]
  reg [63:0] _RAND_27;
  reg [47:0] _T_255_12; // @[Switch.scala 52:30:@2405.4]
  reg [63:0] _RAND_28;
  reg [47:0] _T_255_13; // @[Switch.scala 52:30:@2405.4]
  reg [63:0] _RAND_29;
  reg [47:0] _T_255_14; // @[Switch.scala 52:30:@2405.4]
  reg [63:0] _RAND_30;
  reg [47:0] _T_255_15; // @[Switch.scala 52:30:@2405.4]
  reg [63:0] _RAND_31;
  reg  _T_344_0; // @[Switch.scala 53:31:@2438.4]
  reg [31:0] _RAND_32;
  reg  _T_344_1; // @[Switch.scala 53:31:@2438.4]
  reg [31:0] _RAND_33;
  reg  _T_344_2; // @[Switch.scala 53:31:@2438.4]
  reg [31:0] _RAND_34;
  reg  _T_344_3; // @[Switch.scala 53:31:@2438.4]
  reg [31:0] _RAND_35;
  reg  _T_344_4; // @[Switch.scala 53:31:@2438.4]
  reg [31:0] _RAND_36;
  reg  _T_344_5; // @[Switch.scala 53:31:@2438.4]
  reg [31:0] _RAND_37;
  reg  _T_344_6; // @[Switch.scala 53:31:@2438.4]
  reg [31:0] _RAND_38;
  reg  _T_344_7; // @[Switch.scala 53:31:@2438.4]
  reg [31:0] _RAND_39;
  reg  _T_344_8; // @[Switch.scala 53:31:@2438.4]
  reg [31:0] _RAND_40;
  reg  _T_344_9; // @[Switch.scala 53:31:@2438.4]
  reg [31:0] _RAND_41;
  reg  _T_344_10; // @[Switch.scala 53:31:@2438.4]
  reg [31:0] _RAND_42;
  reg  _T_344_11; // @[Switch.scala 53:31:@2438.4]
  reg [31:0] _RAND_43;
  reg  _T_344_12; // @[Switch.scala 53:31:@2438.4]
  reg [31:0] _RAND_44;
  reg  _T_344_13; // @[Switch.scala 53:31:@2438.4]
  reg [31:0] _RAND_45;
  reg  _T_344_14; // @[Switch.scala 53:31:@2438.4]
  reg [31:0] _RAND_46;
  reg  _T_344_15; // @[Switch.scala 53:31:@2438.4]
  reg [31:0] _RAND_47;
  reg  _T_433_0; // @[Switch.scala 54:23:@2471.4]
  reg [31:0] _RAND_48;
  reg  _T_433_1; // @[Switch.scala 54:23:@2471.4]
  reg [31:0] _RAND_49;
  reg  _T_433_2; // @[Switch.scala 54:23:@2471.4]
  reg [31:0] _RAND_50;
  reg  _T_433_3; // @[Switch.scala 54:23:@2471.4]
  reg [31:0] _RAND_51;
  reg  _T_433_4; // @[Switch.scala 54:23:@2471.4]
  reg [31:0] _RAND_52;
  reg  _T_433_5; // @[Switch.scala 54:23:@2471.4]
  reg [31:0] _RAND_53;
  reg  _T_433_6; // @[Switch.scala 54:23:@2471.4]
  reg [31:0] _RAND_54;
  reg  _T_433_7; // @[Switch.scala 54:23:@2471.4]
  reg [31:0] _RAND_55;
  reg  _T_433_8; // @[Switch.scala 54:23:@2471.4]
  reg [31:0] _RAND_56;
  reg  _T_433_9; // @[Switch.scala 54:23:@2471.4]
  reg [31:0] _RAND_57;
  reg  _T_433_10; // @[Switch.scala 54:23:@2471.4]
  reg [31:0] _RAND_58;
  reg  _T_433_11; // @[Switch.scala 54:23:@2471.4]
  reg [31:0] _RAND_59;
  reg  _T_433_12; // @[Switch.scala 54:23:@2471.4]
  reg [31:0] _RAND_60;
  reg  _T_433_13; // @[Switch.scala 54:23:@2471.4]
  reg [31:0] _RAND_61;
  reg  _T_433_14; // @[Switch.scala 54:23:@2471.4]
  reg [31:0] _RAND_62;
  reg  _T_433_15; // @[Switch.scala 54:23:@2471.4]
  reg [31:0] _RAND_63;
  reg [47:0] _T_522_0; // @[Switch.scala 55:24:@2504.4]
  reg [63:0] _RAND_64;
  reg [47:0] _T_522_1; // @[Switch.scala 55:24:@2504.4]
  reg [63:0] _RAND_65;
  reg [47:0] _T_522_2; // @[Switch.scala 55:24:@2504.4]
  reg [63:0] _RAND_66;
  reg [47:0] _T_522_3; // @[Switch.scala 55:24:@2504.4]
  reg [63:0] _RAND_67;
  reg [47:0] _T_522_4; // @[Switch.scala 55:24:@2504.4]
  reg [63:0] _RAND_68;
  reg [47:0] _T_522_5; // @[Switch.scala 55:24:@2504.4]
  reg [63:0] _RAND_69;
  reg [47:0] _T_522_6; // @[Switch.scala 55:24:@2504.4]
  reg [63:0] _RAND_70;
  reg [47:0] _T_522_7; // @[Switch.scala 55:24:@2504.4]
  reg [63:0] _RAND_71;
  reg [47:0] _T_522_8; // @[Switch.scala 55:24:@2504.4]
  reg [63:0] _RAND_72;
  reg [47:0] _T_522_9; // @[Switch.scala 55:24:@2504.4]
  reg [63:0] _RAND_73;
  reg [47:0] _T_522_10; // @[Switch.scala 55:24:@2504.4]
  reg [63:0] _RAND_74;
  reg [47:0] _T_522_11; // @[Switch.scala 55:24:@2504.4]
  reg [63:0] _RAND_75;
  reg [47:0] _T_522_12; // @[Switch.scala 55:24:@2504.4]
  reg [63:0] _RAND_76;
  reg [47:0] _T_522_13; // @[Switch.scala 55:24:@2504.4]
  reg [63:0] _RAND_77;
  reg [47:0] _T_522_14; // @[Switch.scala 55:24:@2504.4]
  reg [63:0] _RAND_78;
  reg [47:0] _T_522_15; // @[Switch.scala 55:24:@2504.4]
  reg [63:0] _RAND_79;
  reg  _T_611_0; // @[Switch.scala 56:25:@2537.4]
  reg [31:0] _RAND_80;
  reg  _T_611_1; // @[Switch.scala 56:25:@2537.4]
  reg [31:0] _RAND_81;
  reg  _T_611_2; // @[Switch.scala 56:25:@2537.4]
  reg [31:0] _RAND_82;
  reg  _T_611_3; // @[Switch.scala 56:25:@2537.4]
  reg [31:0] _RAND_83;
  reg  _T_611_4; // @[Switch.scala 56:25:@2537.4]
  reg [31:0] _RAND_84;
  reg  _T_611_5; // @[Switch.scala 56:25:@2537.4]
  reg [31:0] _RAND_85;
  reg  _T_611_6; // @[Switch.scala 56:25:@2537.4]
  reg [31:0] _RAND_86;
  reg  _T_611_7; // @[Switch.scala 56:25:@2537.4]
  reg [31:0] _RAND_87;
  reg  _T_611_8; // @[Switch.scala 56:25:@2537.4]
  reg [31:0] _RAND_88;
  reg  _T_611_9; // @[Switch.scala 56:25:@2537.4]
  reg [31:0] _RAND_89;
  reg  _T_611_10; // @[Switch.scala 56:25:@2537.4]
  reg [31:0] _RAND_90;
  reg  _T_611_11; // @[Switch.scala 56:25:@2537.4]
  reg [31:0] _RAND_91;
  reg  _T_611_12; // @[Switch.scala 56:25:@2537.4]
  reg [31:0] _RAND_92;
  reg  _T_611_13; // @[Switch.scala 56:25:@2537.4]
  reg [31:0] _RAND_93;
  reg  _T_611_14; // @[Switch.scala 56:25:@2537.4]
  reg [31:0] _RAND_94;
  reg  _T_611_15; // @[Switch.scala 56:25:@2537.4]
  reg [31:0] _RAND_95;
  Switch switch ( // @[Switch.scala 50:22:@2369.4]
    .io_inAddr_0(switch_io_inAddr_0),
    .io_inAddr_1(switch_io_inAddr_1),
    .io_inAddr_2(switch_io_inAddr_2),
    .io_inAddr_3(switch_io_inAddr_3),
    .io_inAddr_4(switch_io_inAddr_4),
    .io_inAddr_5(switch_io_inAddr_5),
    .io_inAddr_6(switch_io_inAddr_6),
    .io_inAddr_7(switch_io_inAddr_7),
    .io_inAddr_8(switch_io_inAddr_8),
    .io_inAddr_9(switch_io_inAddr_9),
    .io_inAddr_10(switch_io_inAddr_10),
    .io_inAddr_11(switch_io_inAddr_11),
    .io_inAddr_12(switch_io_inAddr_12),
    .io_inAddr_13(switch_io_inAddr_13),
    .io_inAddr_14(switch_io_inAddr_14),
    .io_inAddr_15(switch_io_inAddr_15),
    .io_inData_0(switch_io_inData_0),
    .io_inData_1(switch_io_inData_1),
    .io_inData_2(switch_io_inData_2),
    .io_inData_3(switch_io_inData_3),
    .io_inData_4(switch_io_inData_4),
    .io_inData_5(switch_io_inData_5),
    .io_inData_6(switch_io_inData_6),
    .io_inData_7(switch_io_inData_7),
    .io_inData_8(switch_io_inData_8),
    .io_inData_9(switch_io_inData_9),
    .io_inData_10(switch_io_inData_10),
    .io_inData_11(switch_io_inData_11),
    .io_inData_12(switch_io_inData_12),
    .io_inData_13(switch_io_inData_13),
    .io_inData_14(switch_io_inData_14),
    .io_inData_15(switch_io_inData_15),
    .io_inValid_0(switch_io_inValid_0),
    .io_inValid_1(switch_io_inValid_1),
    .io_inValid_2(switch_io_inValid_2),
    .io_inValid_3(switch_io_inValid_3),
    .io_inValid_4(switch_io_inValid_4),
    .io_inValid_5(switch_io_inValid_5),
    .io_inValid_6(switch_io_inValid_6),
    .io_inValid_7(switch_io_inValid_7),
    .io_inValid_8(switch_io_inValid_8),
    .io_inValid_9(switch_io_inValid_9),
    .io_inValid_10(switch_io_inValid_10),
    .io_inValid_11(switch_io_inValid_11),
    .io_inValid_12(switch_io_inValid_12),
    .io_inValid_13(switch_io_inValid_13),
    .io_inValid_14(switch_io_inValid_14),
    .io_inValid_15(switch_io_inValid_15),
    .io_outAck_0(switch_io_outAck_0),
    .io_outAck_1(switch_io_outAck_1),
    .io_outAck_2(switch_io_outAck_2),
    .io_outAck_3(switch_io_outAck_3),
    .io_outAck_4(switch_io_outAck_4),
    .io_outAck_5(switch_io_outAck_5),
    .io_outAck_6(switch_io_outAck_6),
    .io_outAck_7(switch_io_outAck_7),
    .io_outAck_8(switch_io_outAck_8),
    .io_outAck_9(switch_io_outAck_9),
    .io_outAck_10(switch_io_outAck_10),
    .io_outAck_11(switch_io_outAck_11),
    .io_outAck_12(switch_io_outAck_12),
    .io_outAck_13(switch_io_outAck_13),
    .io_outAck_14(switch_io_outAck_14),
    .io_outAck_15(switch_io_outAck_15),
    .io_outData_0(switch_io_outData_0),
    .io_outData_1(switch_io_outData_1),
    .io_outData_2(switch_io_outData_2),
    .io_outData_3(switch_io_outData_3),
    .io_outData_4(switch_io_outData_4),
    .io_outData_5(switch_io_outData_5),
    .io_outData_6(switch_io_outData_6),
    .io_outData_7(switch_io_outData_7),
    .io_outData_8(switch_io_outData_8),
    .io_outData_9(switch_io_outData_9),
    .io_outData_10(switch_io_outData_10),
    .io_outData_11(switch_io_outData_11),
    .io_outData_12(switch_io_outData_12),
    .io_outData_13(switch_io_outData_13),
    .io_outData_14(switch_io_outData_14),
    .io_outData_15(switch_io_outData_15),
    .io_outValid_0(switch_io_outValid_0),
    .io_outValid_1(switch_io_outValid_1),
    .io_outValid_2(switch_io_outValid_2),
    .io_outValid_3(switch_io_outValid_3),
    .io_outValid_4(switch_io_outValid_4),
    .io_outValid_5(switch_io_outValid_5),
    .io_outValid_6(switch_io_outValid_6),
    .io_outValid_7(switch_io_outValid_7),
    .io_outValid_8(switch_io_outValid_8),
    .io_outValid_9(switch_io_outValid_9),
    .io_outValid_10(switch_io_outValid_10),
    .io_outValid_11(switch_io_outValid_11),
    .io_outValid_12(switch_io_outValid_12),
    .io_outValid_13(switch_io_outValid_13),
    .io_outValid_14(switch_io_outValid_14),
    .io_outValid_15(switch_io_outValid_15)
  );
  assign io_outAck_0 = _T_433_0; // @[Switch.scala 54:13:@2488.4]
  assign io_outAck_1 = _T_433_1; // @[Switch.scala 54:13:@2489.4]
  assign io_outAck_2 = _T_433_2; // @[Switch.scala 54:13:@2490.4]
  assign io_outAck_3 = _T_433_3; // @[Switch.scala 54:13:@2491.4]
  assign io_outAck_4 = _T_433_4; // @[Switch.scala 54:13:@2492.4]
  assign io_outAck_5 = _T_433_5; // @[Switch.scala 54:13:@2493.4]
  assign io_outAck_6 = _T_433_6; // @[Switch.scala 54:13:@2494.4]
  assign io_outAck_7 = _T_433_7; // @[Switch.scala 54:13:@2495.4]
  assign io_outAck_8 = _T_433_8; // @[Switch.scala 54:13:@2496.4]
  assign io_outAck_9 = _T_433_9; // @[Switch.scala 54:13:@2497.4]
  assign io_outAck_10 = _T_433_10; // @[Switch.scala 54:13:@2498.4]
  assign io_outAck_11 = _T_433_11; // @[Switch.scala 54:13:@2499.4]
  assign io_outAck_12 = _T_433_12; // @[Switch.scala 54:13:@2500.4]
  assign io_outAck_13 = _T_433_13; // @[Switch.scala 54:13:@2501.4]
  assign io_outAck_14 = _T_433_14; // @[Switch.scala 54:13:@2502.4]
  assign io_outAck_15 = _T_433_15; // @[Switch.scala 54:13:@2503.4]
  assign io_outData_0 = _T_522_0; // @[Switch.scala 55:14:@2521.4]
  assign io_outData_1 = _T_522_1; // @[Switch.scala 55:14:@2522.4]
  assign io_outData_2 = _T_522_2; // @[Switch.scala 55:14:@2523.4]
  assign io_outData_3 = _T_522_3; // @[Switch.scala 55:14:@2524.4]
  assign io_outData_4 = _T_522_4; // @[Switch.scala 55:14:@2525.4]
  assign io_outData_5 = _T_522_5; // @[Switch.scala 55:14:@2526.4]
  assign io_outData_6 = _T_522_6; // @[Switch.scala 55:14:@2527.4]
  assign io_outData_7 = _T_522_7; // @[Switch.scala 55:14:@2528.4]
  assign io_outData_8 = _T_522_8; // @[Switch.scala 55:14:@2529.4]
  assign io_outData_9 = _T_522_9; // @[Switch.scala 55:14:@2530.4]
  assign io_outData_10 = _T_522_10; // @[Switch.scala 55:14:@2531.4]
  assign io_outData_11 = _T_522_11; // @[Switch.scala 55:14:@2532.4]
  assign io_outData_12 = _T_522_12; // @[Switch.scala 55:14:@2533.4]
  assign io_outData_13 = _T_522_13; // @[Switch.scala 55:14:@2534.4]
  assign io_outData_14 = _T_522_14; // @[Switch.scala 55:14:@2535.4]
  assign io_outData_15 = _T_522_15; // @[Switch.scala 55:14:@2536.4]
  assign io_outValid_0 = _T_611_0; // @[Switch.scala 56:15:@2554.4]
  assign io_outValid_1 = _T_611_1; // @[Switch.scala 56:15:@2555.4]
  assign io_outValid_2 = _T_611_2; // @[Switch.scala 56:15:@2556.4]
  assign io_outValid_3 = _T_611_3; // @[Switch.scala 56:15:@2557.4]
  assign io_outValid_4 = _T_611_4; // @[Switch.scala 56:15:@2558.4]
  assign io_outValid_5 = _T_611_5; // @[Switch.scala 56:15:@2559.4]
  assign io_outValid_6 = _T_611_6; // @[Switch.scala 56:15:@2560.4]
  assign io_outValid_7 = _T_611_7; // @[Switch.scala 56:15:@2561.4]
  assign io_outValid_8 = _T_611_8; // @[Switch.scala 56:15:@2562.4]
  assign io_outValid_9 = _T_611_9; // @[Switch.scala 56:15:@2563.4]
  assign io_outValid_10 = _T_611_10; // @[Switch.scala 56:15:@2564.4]
  assign io_outValid_11 = _T_611_11; // @[Switch.scala 56:15:@2565.4]
  assign io_outValid_12 = _T_611_12; // @[Switch.scala 56:15:@2566.4]
  assign io_outValid_13 = _T_611_13; // @[Switch.scala 56:15:@2567.4]
  assign io_outValid_14 = _T_611_14; // @[Switch.scala 56:15:@2568.4]
  assign io_outValid_15 = _T_611_15; // @[Switch.scala 56:15:@2569.4]
  assign switch_io_inAddr_0 = _T_166_0; // @[Switch.scala 51:20:@2389.4]
  assign switch_io_inAddr_1 = _T_166_1; // @[Switch.scala 51:20:@2390.4]
  assign switch_io_inAddr_2 = _T_166_2; // @[Switch.scala 51:20:@2391.4]
  assign switch_io_inAddr_3 = _T_166_3; // @[Switch.scala 51:20:@2392.4]
  assign switch_io_inAddr_4 = _T_166_4; // @[Switch.scala 51:20:@2393.4]
  assign switch_io_inAddr_5 = _T_166_5; // @[Switch.scala 51:20:@2394.4]
  assign switch_io_inAddr_6 = _T_166_6; // @[Switch.scala 51:20:@2395.4]
  assign switch_io_inAddr_7 = _T_166_7; // @[Switch.scala 51:20:@2396.4]
  assign switch_io_inAddr_8 = _T_166_8; // @[Switch.scala 51:20:@2397.4]
  assign switch_io_inAddr_9 = _T_166_9; // @[Switch.scala 51:20:@2398.4]
  assign switch_io_inAddr_10 = _T_166_10; // @[Switch.scala 51:20:@2399.4]
  assign switch_io_inAddr_11 = _T_166_11; // @[Switch.scala 51:20:@2400.4]
  assign switch_io_inAddr_12 = _T_166_12; // @[Switch.scala 51:20:@2401.4]
  assign switch_io_inAddr_13 = _T_166_13; // @[Switch.scala 51:20:@2402.4]
  assign switch_io_inAddr_14 = _T_166_14; // @[Switch.scala 51:20:@2403.4]
  assign switch_io_inAddr_15 = _T_166_15; // @[Switch.scala 51:20:@2404.4]
  assign switch_io_inData_0 = _T_255_0; // @[Switch.scala 52:20:@2422.4]
  assign switch_io_inData_1 = _T_255_1; // @[Switch.scala 52:20:@2423.4]
  assign switch_io_inData_2 = _T_255_2; // @[Switch.scala 52:20:@2424.4]
  assign switch_io_inData_3 = _T_255_3; // @[Switch.scala 52:20:@2425.4]
  assign switch_io_inData_4 = _T_255_4; // @[Switch.scala 52:20:@2426.4]
  assign switch_io_inData_5 = _T_255_5; // @[Switch.scala 52:20:@2427.4]
  assign switch_io_inData_6 = _T_255_6; // @[Switch.scala 52:20:@2428.4]
  assign switch_io_inData_7 = _T_255_7; // @[Switch.scala 52:20:@2429.4]
  assign switch_io_inData_8 = _T_255_8; // @[Switch.scala 52:20:@2430.4]
  assign switch_io_inData_9 = _T_255_9; // @[Switch.scala 52:20:@2431.4]
  assign switch_io_inData_10 = _T_255_10; // @[Switch.scala 52:20:@2432.4]
  assign switch_io_inData_11 = _T_255_11; // @[Switch.scala 52:20:@2433.4]
  assign switch_io_inData_12 = _T_255_12; // @[Switch.scala 52:20:@2434.4]
  assign switch_io_inData_13 = _T_255_13; // @[Switch.scala 52:20:@2435.4]
  assign switch_io_inData_14 = _T_255_14; // @[Switch.scala 52:20:@2436.4]
  assign switch_io_inData_15 = _T_255_15; // @[Switch.scala 52:20:@2437.4]
  assign switch_io_inValid_0 = _T_344_0; // @[Switch.scala 53:21:@2455.4]
  assign switch_io_inValid_1 = _T_344_1; // @[Switch.scala 53:21:@2456.4]
  assign switch_io_inValid_2 = _T_344_2; // @[Switch.scala 53:21:@2457.4]
  assign switch_io_inValid_3 = _T_344_3; // @[Switch.scala 53:21:@2458.4]
  assign switch_io_inValid_4 = _T_344_4; // @[Switch.scala 53:21:@2459.4]
  assign switch_io_inValid_5 = _T_344_5; // @[Switch.scala 53:21:@2460.4]
  assign switch_io_inValid_6 = _T_344_6; // @[Switch.scala 53:21:@2461.4]
  assign switch_io_inValid_7 = _T_344_7; // @[Switch.scala 53:21:@2462.4]
  assign switch_io_inValid_8 = _T_344_8; // @[Switch.scala 53:21:@2463.4]
  assign switch_io_inValid_9 = _T_344_9; // @[Switch.scala 53:21:@2464.4]
  assign switch_io_inValid_10 = _T_344_10; // @[Switch.scala 53:21:@2465.4]
  assign switch_io_inValid_11 = _T_344_11; // @[Switch.scala 53:21:@2466.4]
  assign switch_io_inValid_12 = _T_344_12; // @[Switch.scala 53:21:@2467.4]
  assign switch_io_inValid_13 = _T_344_13; // @[Switch.scala 53:21:@2468.4]
  assign switch_io_inValid_14 = _T_344_14; // @[Switch.scala 53:21:@2469.4]
  assign switch_io_inValid_15 = _T_344_15; // @[Switch.scala 53:21:@2470.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_166_0 = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_166_1 = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_166_2 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_166_3 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_166_4 = _RAND_4[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_166_5 = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_166_6 = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_166_7 = _RAND_7[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_166_8 = _RAND_8[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_166_9 = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_166_10 = _RAND_10[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_166_11 = _RAND_11[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_166_12 = _RAND_12[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_166_13 = _RAND_13[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_166_14 = _RAND_14[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_166_15 = _RAND_15[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {2{`RANDOM}};
  _T_255_0 = _RAND_16[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {2{`RANDOM}};
  _T_255_1 = _RAND_17[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {2{`RANDOM}};
  _T_255_2 = _RAND_18[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {2{`RANDOM}};
  _T_255_3 = _RAND_19[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {2{`RANDOM}};
  _T_255_4 = _RAND_20[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {2{`RANDOM}};
  _T_255_5 = _RAND_21[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {2{`RANDOM}};
  _T_255_6 = _RAND_22[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {2{`RANDOM}};
  _T_255_7 = _RAND_23[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {2{`RANDOM}};
  _T_255_8 = _RAND_24[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {2{`RANDOM}};
  _T_255_9 = _RAND_25[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {2{`RANDOM}};
  _T_255_10 = _RAND_26[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {2{`RANDOM}};
  _T_255_11 = _RAND_27[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {2{`RANDOM}};
  _T_255_12 = _RAND_28[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {2{`RANDOM}};
  _T_255_13 = _RAND_29[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {2{`RANDOM}};
  _T_255_14 = _RAND_30[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {2{`RANDOM}};
  _T_255_15 = _RAND_31[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_344_0 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_344_1 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_344_2 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_344_3 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_344_4 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_344_5 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_344_6 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_344_7 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_344_8 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_344_9 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_344_10 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_344_11 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_344_12 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_344_13 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_344_14 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_344_15 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_433_0 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_433_1 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_433_2 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_433_3 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_433_4 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_433_5 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_433_6 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_433_7 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_433_8 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_433_9 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_433_10 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_433_11 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_433_12 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_433_13 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_433_14 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_433_15 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {2{`RANDOM}};
  _T_522_0 = _RAND_64[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {2{`RANDOM}};
  _T_522_1 = _RAND_65[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {2{`RANDOM}};
  _T_522_2 = _RAND_66[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {2{`RANDOM}};
  _T_522_3 = _RAND_67[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {2{`RANDOM}};
  _T_522_4 = _RAND_68[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {2{`RANDOM}};
  _T_522_5 = _RAND_69[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {2{`RANDOM}};
  _T_522_6 = _RAND_70[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {2{`RANDOM}};
  _T_522_7 = _RAND_71[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {2{`RANDOM}};
  _T_522_8 = _RAND_72[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {2{`RANDOM}};
  _T_522_9 = _RAND_73[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {2{`RANDOM}};
  _T_522_10 = _RAND_74[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {2{`RANDOM}};
  _T_522_11 = _RAND_75[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {2{`RANDOM}};
  _T_522_12 = _RAND_76[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {2{`RANDOM}};
  _T_522_13 = _RAND_77[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {2{`RANDOM}};
  _T_522_14 = _RAND_78[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {2{`RANDOM}};
  _T_522_15 = _RAND_79[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_611_0 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_611_1 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_611_2 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_611_3 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_611_4 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_611_5 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_611_6 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_611_7 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_611_8 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_611_9 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_611_10 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_611_11 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_611_12 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_611_13 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_611_14 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_611_15 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    _T_166_0 <= io_inAddr_0;
    _T_166_1 <= io_inAddr_1;
    _T_166_2 <= io_inAddr_2;
    _T_166_3 <= io_inAddr_3;
    _T_166_4 <= io_inAddr_4;
    _T_166_5 <= io_inAddr_5;
    _T_166_6 <= io_inAddr_6;
    _T_166_7 <= io_inAddr_7;
    _T_166_8 <= io_inAddr_8;
    _T_166_9 <= io_inAddr_9;
    _T_166_10 <= io_inAddr_10;
    _T_166_11 <= io_inAddr_11;
    _T_166_12 <= io_inAddr_12;
    _T_166_13 <= io_inAddr_13;
    _T_166_14 <= io_inAddr_14;
    _T_166_15 <= io_inAddr_15;
    _T_255_0 <= io_inData_0;
    _T_255_1 <= io_inData_1;
    _T_255_2 <= io_inData_2;
    _T_255_3 <= io_inData_3;
    _T_255_4 <= io_inData_4;
    _T_255_5 <= io_inData_5;
    _T_255_6 <= io_inData_6;
    _T_255_7 <= io_inData_7;
    _T_255_8 <= io_inData_8;
    _T_255_9 <= io_inData_9;
    _T_255_10 <= io_inData_10;
    _T_255_11 <= io_inData_11;
    _T_255_12 <= io_inData_12;
    _T_255_13 <= io_inData_13;
    _T_255_14 <= io_inData_14;
    _T_255_15 <= io_inData_15;
    _T_344_0 <= io_inValid_0;
    _T_344_1 <= io_inValid_1;
    _T_344_2 <= io_inValid_2;
    _T_344_3 <= io_inValid_3;
    _T_344_4 <= io_inValid_4;
    _T_344_5 <= io_inValid_5;
    _T_344_6 <= io_inValid_6;
    _T_344_7 <= io_inValid_7;
    _T_344_8 <= io_inValid_8;
    _T_344_9 <= io_inValid_9;
    _T_344_10 <= io_inValid_10;
    _T_344_11 <= io_inValid_11;
    _T_344_12 <= io_inValid_12;
    _T_344_13 <= io_inValid_13;
    _T_344_14 <= io_inValid_14;
    _T_344_15 <= io_inValid_15;
    _T_433_0 <= switch_io_outAck_0;
    _T_433_1 <= switch_io_outAck_1;
    _T_433_2 <= switch_io_outAck_2;
    _T_433_3 <= switch_io_outAck_3;
    _T_433_4 <= switch_io_outAck_4;
    _T_433_5 <= switch_io_outAck_5;
    _T_433_6 <= switch_io_outAck_6;
    _T_433_7 <= switch_io_outAck_7;
    _T_433_8 <= switch_io_outAck_8;
    _T_433_9 <= switch_io_outAck_9;
    _T_433_10 <= switch_io_outAck_10;
    _T_433_11 <= switch_io_outAck_11;
    _T_433_12 <= switch_io_outAck_12;
    _T_433_13 <= switch_io_outAck_13;
    _T_433_14 <= switch_io_outAck_14;
    _T_433_15 <= switch_io_outAck_15;
    _T_522_0 <= switch_io_outData_0;
    _T_522_1 <= switch_io_outData_1;
    _T_522_2 <= switch_io_outData_2;
    _T_522_3 <= switch_io_outData_3;
    _T_522_4 <= switch_io_outData_4;
    _T_522_5 <= switch_io_outData_5;
    _T_522_6 <= switch_io_outData_6;
    _T_522_7 <= switch_io_outData_7;
    _T_522_8 <= switch_io_outData_8;
    _T_522_9 <= switch_io_outData_9;
    _T_522_10 <= switch_io_outData_10;
    _T_522_11 <= switch_io_outData_11;
    _T_522_12 <= switch_io_outData_12;
    _T_522_13 <= switch_io_outData_13;
    _T_522_14 <= switch_io_outData_14;
    _T_522_15 <= switch_io_outData_15;
    _T_611_0 <= switch_io_outValid_0;
    _T_611_1 <= switch_io_outValid_1;
    _T_611_2 <= switch_io_outValid_2;
    _T_611_3 <= switch_io_outValid_3;
    _T_611_4 <= switch_io_outValid_4;
    _T_611_5 <= switch_io_outValid_5;
    _T_611_6 <= switch_io_outValid_6;
    _T_611_7 <= switch_io_outValid_7;
    _T_611_8 <= switch_io_outValid_8;
    _T_611_9 <= switch_io_outValid_9;
    _T_611_10 <= switch_io_outValid_10;
    _T_611_11 <= switch_io_outValid_11;
    _T_611_12 <= switch_io_outValid_12;
    _T_611_13 <= switch_io_outValid_13;
    _T_611_14 <= switch_io_outValid_14;
    _T_611_15 <= switch_io_outValid_15;
  end
endmodule
