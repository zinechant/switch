module Switch( // @[:@3.2]
  input  [5:0]  io_inAddr_0, // @[:@6.4]
  input  [5:0]  io_inAddr_1, // @[:@6.4]
  input  [5:0]  io_inAddr_2, // @[:@6.4]
  input  [5:0]  io_inAddr_3, // @[:@6.4]
  input  [5:0]  io_inAddr_4, // @[:@6.4]
  input  [5:0]  io_inAddr_5, // @[:@6.4]
  input  [5:0]  io_inAddr_6, // @[:@6.4]
  input  [5:0]  io_inAddr_7, // @[:@6.4]
  input  [5:0]  io_inAddr_8, // @[:@6.4]
  input  [5:0]  io_inAddr_9, // @[:@6.4]
  input  [5:0]  io_inAddr_10, // @[:@6.4]
  input  [5:0]  io_inAddr_11, // @[:@6.4]
  input  [5:0]  io_inAddr_12, // @[:@6.4]
  input  [5:0]  io_inAddr_13, // @[:@6.4]
  input  [5:0]  io_inAddr_14, // @[:@6.4]
  input  [5:0]  io_inAddr_15, // @[:@6.4]
  input  [5:0]  io_inAddr_16, // @[:@6.4]
  input  [5:0]  io_inAddr_17, // @[:@6.4]
  input  [5:0]  io_inAddr_18, // @[:@6.4]
  input  [5:0]  io_inAddr_19, // @[:@6.4]
  input  [5:0]  io_inAddr_20, // @[:@6.4]
  input  [5:0]  io_inAddr_21, // @[:@6.4]
  input  [5:0]  io_inAddr_22, // @[:@6.4]
  input  [5:0]  io_inAddr_23, // @[:@6.4]
  input  [5:0]  io_inAddr_24, // @[:@6.4]
  input  [5:0]  io_inAddr_25, // @[:@6.4]
  input  [5:0]  io_inAddr_26, // @[:@6.4]
  input  [5:0]  io_inAddr_27, // @[:@6.4]
  input  [5:0]  io_inAddr_28, // @[:@6.4]
  input  [5:0]  io_inAddr_29, // @[:@6.4]
  input  [5:0]  io_inAddr_30, // @[:@6.4]
  input  [5:0]  io_inAddr_31, // @[:@6.4]
  input  [5:0]  io_inAddr_32, // @[:@6.4]
  input  [5:0]  io_inAddr_33, // @[:@6.4]
  input  [5:0]  io_inAddr_34, // @[:@6.4]
  input  [5:0]  io_inAddr_35, // @[:@6.4]
  input  [5:0]  io_inAddr_36, // @[:@6.4]
  input  [5:0]  io_inAddr_37, // @[:@6.4]
  input  [5:0]  io_inAddr_38, // @[:@6.4]
  input  [5:0]  io_inAddr_39, // @[:@6.4]
  input  [5:0]  io_inAddr_40, // @[:@6.4]
  input  [5:0]  io_inAddr_41, // @[:@6.4]
  input  [5:0]  io_inAddr_42, // @[:@6.4]
  input  [5:0]  io_inAddr_43, // @[:@6.4]
  input  [5:0]  io_inAddr_44, // @[:@6.4]
  input  [5:0]  io_inAddr_45, // @[:@6.4]
  input  [5:0]  io_inAddr_46, // @[:@6.4]
  input  [5:0]  io_inAddr_47, // @[:@6.4]
  input  [5:0]  io_inAddr_48, // @[:@6.4]
  input  [5:0]  io_inAddr_49, // @[:@6.4]
  input  [5:0]  io_inAddr_50, // @[:@6.4]
  input  [5:0]  io_inAddr_51, // @[:@6.4]
  input  [5:0]  io_inAddr_52, // @[:@6.4]
  input  [5:0]  io_inAddr_53, // @[:@6.4]
  input  [5:0]  io_inAddr_54, // @[:@6.4]
  input  [5:0]  io_inAddr_55, // @[:@6.4]
  input  [5:0]  io_inAddr_56, // @[:@6.4]
  input  [5:0]  io_inAddr_57, // @[:@6.4]
  input  [5:0]  io_inAddr_58, // @[:@6.4]
  input  [5:0]  io_inAddr_59, // @[:@6.4]
  input  [5:0]  io_inAddr_60, // @[:@6.4]
  input  [5:0]  io_inAddr_61, // @[:@6.4]
  input  [5:0]  io_inAddr_62, // @[:@6.4]
  input  [5:0]  io_inAddr_63, // @[:@6.4]
  input  [47:0] io_inData_0, // @[:@6.4]
  input  [47:0] io_inData_1, // @[:@6.4]
  input  [47:0] io_inData_2, // @[:@6.4]
  input  [47:0] io_inData_3, // @[:@6.4]
  input  [47:0] io_inData_4, // @[:@6.4]
  input  [47:0] io_inData_5, // @[:@6.4]
  input  [47:0] io_inData_6, // @[:@6.4]
  input  [47:0] io_inData_7, // @[:@6.4]
  input  [47:0] io_inData_8, // @[:@6.4]
  input  [47:0] io_inData_9, // @[:@6.4]
  input  [47:0] io_inData_10, // @[:@6.4]
  input  [47:0] io_inData_11, // @[:@6.4]
  input  [47:0] io_inData_12, // @[:@6.4]
  input  [47:0] io_inData_13, // @[:@6.4]
  input  [47:0] io_inData_14, // @[:@6.4]
  input  [47:0] io_inData_15, // @[:@6.4]
  input  [47:0] io_inData_16, // @[:@6.4]
  input  [47:0] io_inData_17, // @[:@6.4]
  input  [47:0] io_inData_18, // @[:@6.4]
  input  [47:0] io_inData_19, // @[:@6.4]
  input  [47:0] io_inData_20, // @[:@6.4]
  input  [47:0] io_inData_21, // @[:@6.4]
  input  [47:0] io_inData_22, // @[:@6.4]
  input  [47:0] io_inData_23, // @[:@6.4]
  input  [47:0] io_inData_24, // @[:@6.4]
  input  [47:0] io_inData_25, // @[:@6.4]
  input  [47:0] io_inData_26, // @[:@6.4]
  input  [47:0] io_inData_27, // @[:@6.4]
  input  [47:0] io_inData_28, // @[:@6.4]
  input  [47:0] io_inData_29, // @[:@6.4]
  input  [47:0] io_inData_30, // @[:@6.4]
  input  [47:0] io_inData_31, // @[:@6.4]
  input  [47:0] io_inData_32, // @[:@6.4]
  input  [47:0] io_inData_33, // @[:@6.4]
  input  [47:0] io_inData_34, // @[:@6.4]
  input  [47:0] io_inData_35, // @[:@6.4]
  input  [47:0] io_inData_36, // @[:@6.4]
  input  [47:0] io_inData_37, // @[:@6.4]
  input  [47:0] io_inData_38, // @[:@6.4]
  input  [47:0] io_inData_39, // @[:@6.4]
  input  [47:0] io_inData_40, // @[:@6.4]
  input  [47:0] io_inData_41, // @[:@6.4]
  input  [47:0] io_inData_42, // @[:@6.4]
  input  [47:0] io_inData_43, // @[:@6.4]
  input  [47:0] io_inData_44, // @[:@6.4]
  input  [47:0] io_inData_45, // @[:@6.4]
  input  [47:0] io_inData_46, // @[:@6.4]
  input  [47:0] io_inData_47, // @[:@6.4]
  input  [47:0] io_inData_48, // @[:@6.4]
  input  [47:0] io_inData_49, // @[:@6.4]
  input  [47:0] io_inData_50, // @[:@6.4]
  input  [47:0] io_inData_51, // @[:@6.4]
  input  [47:0] io_inData_52, // @[:@6.4]
  input  [47:0] io_inData_53, // @[:@6.4]
  input  [47:0] io_inData_54, // @[:@6.4]
  input  [47:0] io_inData_55, // @[:@6.4]
  input  [47:0] io_inData_56, // @[:@6.4]
  input  [47:0] io_inData_57, // @[:@6.4]
  input  [47:0] io_inData_58, // @[:@6.4]
  input  [47:0] io_inData_59, // @[:@6.4]
  input  [47:0] io_inData_60, // @[:@6.4]
  input  [47:0] io_inData_61, // @[:@6.4]
  input  [47:0] io_inData_62, // @[:@6.4]
  input  [47:0] io_inData_63, // @[:@6.4]
  input         io_inValid_0, // @[:@6.4]
  input         io_inValid_1, // @[:@6.4]
  input         io_inValid_2, // @[:@6.4]
  input         io_inValid_3, // @[:@6.4]
  input         io_inValid_4, // @[:@6.4]
  input         io_inValid_5, // @[:@6.4]
  input         io_inValid_6, // @[:@6.4]
  input         io_inValid_7, // @[:@6.4]
  input         io_inValid_8, // @[:@6.4]
  input         io_inValid_9, // @[:@6.4]
  input         io_inValid_10, // @[:@6.4]
  input         io_inValid_11, // @[:@6.4]
  input         io_inValid_12, // @[:@6.4]
  input         io_inValid_13, // @[:@6.4]
  input         io_inValid_14, // @[:@6.4]
  input         io_inValid_15, // @[:@6.4]
  input         io_inValid_16, // @[:@6.4]
  input         io_inValid_17, // @[:@6.4]
  input         io_inValid_18, // @[:@6.4]
  input         io_inValid_19, // @[:@6.4]
  input         io_inValid_20, // @[:@6.4]
  input         io_inValid_21, // @[:@6.4]
  input         io_inValid_22, // @[:@6.4]
  input         io_inValid_23, // @[:@6.4]
  input         io_inValid_24, // @[:@6.4]
  input         io_inValid_25, // @[:@6.4]
  input         io_inValid_26, // @[:@6.4]
  input         io_inValid_27, // @[:@6.4]
  input         io_inValid_28, // @[:@6.4]
  input         io_inValid_29, // @[:@6.4]
  input         io_inValid_30, // @[:@6.4]
  input         io_inValid_31, // @[:@6.4]
  input         io_inValid_32, // @[:@6.4]
  input         io_inValid_33, // @[:@6.4]
  input         io_inValid_34, // @[:@6.4]
  input         io_inValid_35, // @[:@6.4]
  input         io_inValid_36, // @[:@6.4]
  input         io_inValid_37, // @[:@6.4]
  input         io_inValid_38, // @[:@6.4]
  input         io_inValid_39, // @[:@6.4]
  input         io_inValid_40, // @[:@6.4]
  input         io_inValid_41, // @[:@6.4]
  input         io_inValid_42, // @[:@6.4]
  input         io_inValid_43, // @[:@6.4]
  input         io_inValid_44, // @[:@6.4]
  input         io_inValid_45, // @[:@6.4]
  input         io_inValid_46, // @[:@6.4]
  input         io_inValid_47, // @[:@6.4]
  input         io_inValid_48, // @[:@6.4]
  input         io_inValid_49, // @[:@6.4]
  input         io_inValid_50, // @[:@6.4]
  input         io_inValid_51, // @[:@6.4]
  input         io_inValid_52, // @[:@6.4]
  input         io_inValid_53, // @[:@6.4]
  input         io_inValid_54, // @[:@6.4]
  input         io_inValid_55, // @[:@6.4]
  input         io_inValid_56, // @[:@6.4]
  input         io_inValid_57, // @[:@6.4]
  input         io_inValid_58, // @[:@6.4]
  input         io_inValid_59, // @[:@6.4]
  input         io_inValid_60, // @[:@6.4]
  input         io_inValid_61, // @[:@6.4]
  input         io_inValid_62, // @[:@6.4]
  input         io_inValid_63, // @[:@6.4]
  output        io_outAck_0, // @[:@6.4]
  output        io_outAck_1, // @[:@6.4]
  output        io_outAck_2, // @[:@6.4]
  output        io_outAck_3, // @[:@6.4]
  output        io_outAck_4, // @[:@6.4]
  output        io_outAck_5, // @[:@6.4]
  output        io_outAck_6, // @[:@6.4]
  output        io_outAck_7, // @[:@6.4]
  output        io_outAck_8, // @[:@6.4]
  output        io_outAck_9, // @[:@6.4]
  output        io_outAck_10, // @[:@6.4]
  output        io_outAck_11, // @[:@6.4]
  output        io_outAck_12, // @[:@6.4]
  output        io_outAck_13, // @[:@6.4]
  output        io_outAck_14, // @[:@6.4]
  output        io_outAck_15, // @[:@6.4]
  output        io_outAck_16, // @[:@6.4]
  output        io_outAck_17, // @[:@6.4]
  output        io_outAck_18, // @[:@6.4]
  output        io_outAck_19, // @[:@6.4]
  output        io_outAck_20, // @[:@6.4]
  output        io_outAck_21, // @[:@6.4]
  output        io_outAck_22, // @[:@6.4]
  output        io_outAck_23, // @[:@6.4]
  output        io_outAck_24, // @[:@6.4]
  output        io_outAck_25, // @[:@6.4]
  output        io_outAck_26, // @[:@6.4]
  output        io_outAck_27, // @[:@6.4]
  output        io_outAck_28, // @[:@6.4]
  output        io_outAck_29, // @[:@6.4]
  output        io_outAck_30, // @[:@6.4]
  output        io_outAck_31, // @[:@6.4]
  output        io_outAck_32, // @[:@6.4]
  output        io_outAck_33, // @[:@6.4]
  output        io_outAck_34, // @[:@6.4]
  output        io_outAck_35, // @[:@6.4]
  output        io_outAck_36, // @[:@6.4]
  output        io_outAck_37, // @[:@6.4]
  output        io_outAck_38, // @[:@6.4]
  output        io_outAck_39, // @[:@6.4]
  output        io_outAck_40, // @[:@6.4]
  output        io_outAck_41, // @[:@6.4]
  output        io_outAck_42, // @[:@6.4]
  output        io_outAck_43, // @[:@6.4]
  output        io_outAck_44, // @[:@6.4]
  output        io_outAck_45, // @[:@6.4]
  output        io_outAck_46, // @[:@6.4]
  output        io_outAck_47, // @[:@6.4]
  output        io_outAck_48, // @[:@6.4]
  output        io_outAck_49, // @[:@6.4]
  output        io_outAck_50, // @[:@6.4]
  output        io_outAck_51, // @[:@6.4]
  output        io_outAck_52, // @[:@6.4]
  output        io_outAck_53, // @[:@6.4]
  output        io_outAck_54, // @[:@6.4]
  output        io_outAck_55, // @[:@6.4]
  output        io_outAck_56, // @[:@6.4]
  output        io_outAck_57, // @[:@6.4]
  output        io_outAck_58, // @[:@6.4]
  output        io_outAck_59, // @[:@6.4]
  output        io_outAck_60, // @[:@6.4]
  output        io_outAck_61, // @[:@6.4]
  output        io_outAck_62, // @[:@6.4]
  output        io_outAck_63, // @[:@6.4]
  output [47:0] io_outData_0, // @[:@6.4]
  output [47:0] io_outData_1, // @[:@6.4]
  output [47:0] io_outData_2, // @[:@6.4]
  output [47:0] io_outData_3, // @[:@6.4]
  output [47:0] io_outData_4, // @[:@6.4]
  output [47:0] io_outData_5, // @[:@6.4]
  output [47:0] io_outData_6, // @[:@6.4]
  output [47:0] io_outData_7, // @[:@6.4]
  output [47:0] io_outData_8, // @[:@6.4]
  output [47:0] io_outData_9, // @[:@6.4]
  output [47:0] io_outData_10, // @[:@6.4]
  output [47:0] io_outData_11, // @[:@6.4]
  output [47:0] io_outData_12, // @[:@6.4]
  output [47:0] io_outData_13, // @[:@6.4]
  output [47:0] io_outData_14, // @[:@6.4]
  output [47:0] io_outData_15, // @[:@6.4]
  output [47:0] io_outData_16, // @[:@6.4]
  output [47:0] io_outData_17, // @[:@6.4]
  output [47:0] io_outData_18, // @[:@6.4]
  output [47:0] io_outData_19, // @[:@6.4]
  output [47:0] io_outData_20, // @[:@6.4]
  output [47:0] io_outData_21, // @[:@6.4]
  output [47:0] io_outData_22, // @[:@6.4]
  output [47:0] io_outData_23, // @[:@6.4]
  output [47:0] io_outData_24, // @[:@6.4]
  output [47:0] io_outData_25, // @[:@6.4]
  output [47:0] io_outData_26, // @[:@6.4]
  output [47:0] io_outData_27, // @[:@6.4]
  output [47:0] io_outData_28, // @[:@6.4]
  output [47:0] io_outData_29, // @[:@6.4]
  output [47:0] io_outData_30, // @[:@6.4]
  output [47:0] io_outData_31, // @[:@6.4]
  output [47:0] io_outData_32, // @[:@6.4]
  output [47:0] io_outData_33, // @[:@6.4]
  output [47:0] io_outData_34, // @[:@6.4]
  output [47:0] io_outData_35, // @[:@6.4]
  output [47:0] io_outData_36, // @[:@6.4]
  output [47:0] io_outData_37, // @[:@6.4]
  output [47:0] io_outData_38, // @[:@6.4]
  output [47:0] io_outData_39, // @[:@6.4]
  output [47:0] io_outData_40, // @[:@6.4]
  output [47:0] io_outData_41, // @[:@6.4]
  output [47:0] io_outData_42, // @[:@6.4]
  output [47:0] io_outData_43, // @[:@6.4]
  output [47:0] io_outData_44, // @[:@6.4]
  output [47:0] io_outData_45, // @[:@6.4]
  output [47:0] io_outData_46, // @[:@6.4]
  output [47:0] io_outData_47, // @[:@6.4]
  output [47:0] io_outData_48, // @[:@6.4]
  output [47:0] io_outData_49, // @[:@6.4]
  output [47:0] io_outData_50, // @[:@6.4]
  output [47:0] io_outData_51, // @[:@6.4]
  output [47:0] io_outData_52, // @[:@6.4]
  output [47:0] io_outData_53, // @[:@6.4]
  output [47:0] io_outData_54, // @[:@6.4]
  output [47:0] io_outData_55, // @[:@6.4]
  output [47:0] io_outData_56, // @[:@6.4]
  output [47:0] io_outData_57, // @[:@6.4]
  output [47:0] io_outData_58, // @[:@6.4]
  output [47:0] io_outData_59, // @[:@6.4]
  output [47:0] io_outData_60, // @[:@6.4]
  output [47:0] io_outData_61, // @[:@6.4]
  output [47:0] io_outData_62, // @[:@6.4]
  output [47:0] io_outData_63, // @[:@6.4]
  output        io_outValid_0, // @[:@6.4]
  output        io_outValid_1, // @[:@6.4]
  output        io_outValid_2, // @[:@6.4]
  output        io_outValid_3, // @[:@6.4]
  output        io_outValid_4, // @[:@6.4]
  output        io_outValid_5, // @[:@6.4]
  output        io_outValid_6, // @[:@6.4]
  output        io_outValid_7, // @[:@6.4]
  output        io_outValid_8, // @[:@6.4]
  output        io_outValid_9, // @[:@6.4]
  output        io_outValid_10, // @[:@6.4]
  output        io_outValid_11, // @[:@6.4]
  output        io_outValid_12, // @[:@6.4]
  output        io_outValid_13, // @[:@6.4]
  output        io_outValid_14, // @[:@6.4]
  output        io_outValid_15, // @[:@6.4]
  output        io_outValid_16, // @[:@6.4]
  output        io_outValid_17, // @[:@6.4]
  output        io_outValid_18, // @[:@6.4]
  output        io_outValid_19, // @[:@6.4]
  output        io_outValid_20, // @[:@6.4]
  output        io_outValid_21, // @[:@6.4]
  output        io_outValid_22, // @[:@6.4]
  output        io_outValid_23, // @[:@6.4]
  output        io_outValid_24, // @[:@6.4]
  output        io_outValid_25, // @[:@6.4]
  output        io_outValid_26, // @[:@6.4]
  output        io_outValid_27, // @[:@6.4]
  output        io_outValid_28, // @[:@6.4]
  output        io_outValid_29, // @[:@6.4]
  output        io_outValid_30, // @[:@6.4]
  output        io_outValid_31, // @[:@6.4]
  output        io_outValid_32, // @[:@6.4]
  output        io_outValid_33, // @[:@6.4]
  output        io_outValid_34, // @[:@6.4]
  output        io_outValid_35, // @[:@6.4]
  output        io_outValid_36, // @[:@6.4]
  output        io_outValid_37, // @[:@6.4]
  output        io_outValid_38, // @[:@6.4]
  output        io_outValid_39, // @[:@6.4]
  output        io_outValid_40, // @[:@6.4]
  output        io_outValid_41, // @[:@6.4]
  output        io_outValid_42, // @[:@6.4]
  output        io_outValid_43, // @[:@6.4]
  output        io_outValid_44, // @[:@6.4]
  output        io_outValid_45, // @[:@6.4]
  output        io_outValid_46, // @[:@6.4]
  output        io_outValid_47, // @[:@6.4]
  output        io_outValid_48, // @[:@6.4]
  output        io_outValid_49, // @[:@6.4]
  output        io_outValid_50, // @[:@6.4]
  output        io_outValid_51, // @[:@6.4]
  output        io_outValid_52, // @[:@6.4]
  output        io_outValid_53, // @[:@6.4]
  output        io_outValid_54, // @[:@6.4]
  output        io_outValid_55, // @[:@6.4]
  output        io_outValid_56, // @[:@6.4]
  output        io_outValid_57, // @[:@6.4]
  output        io_outValid_58, // @[:@6.4]
  output        io_outValid_59, // @[:@6.4]
  output        io_outValid_60, // @[:@6.4]
  output        io_outValid_61, // @[:@6.4]
  output        io_outValid_62, // @[:@6.4]
  output        io_outValid_63 // @[:@6.4]
);
  wire  _T_17654; // @[Switch.scala 30:53:@10.4]
  wire  valid_0_0; // @[Switch.scala 30:36:@11.4]
  wire  _T_17657; // @[Switch.scala 30:53:@13.4]
  wire  valid_0_1; // @[Switch.scala 30:36:@14.4]
  wire  _T_17660; // @[Switch.scala 30:53:@16.4]
  wire  valid_0_2; // @[Switch.scala 30:36:@17.4]
  wire  _T_17663; // @[Switch.scala 30:53:@19.4]
  wire  valid_0_3; // @[Switch.scala 30:36:@20.4]
  wire  _T_17666; // @[Switch.scala 30:53:@22.4]
  wire  valid_0_4; // @[Switch.scala 30:36:@23.4]
  wire  _T_17669; // @[Switch.scala 30:53:@25.4]
  wire  valid_0_5; // @[Switch.scala 30:36:@26.4]
  wire  _T_17672; // @[Switch.scala 30:53:@28.4]
  wire  valid_0_6; // @[Switch.scala 30:36:@29.4]
  wire  _T_17675; // @[Switch.scala 30:53:@31.4]
  wire  valid_0_7; // @[Switch.scala 30:36:@32.4]
  wire  _T_17678; // @[Switch.scala 30:53:@34.4]
  wire  valid_0_8; // @[Switch.scala 30:36:@35.4]
  wire  _T_17681; // @[Switch.scala 30:53:@37.4]
  wire  valid_0_9; // @[Switch.scala 30:36:@38.4]
  wire  _T_17684; // @[Switch.scala 30:53:@40.4]
  wire  valid_0_10; // @[Switch.scala 30:36:@41.4]
  wire  _T_17687; // @[Switch.scala 30:53:@43.4]
  wire  valid_0_11; // @[Switch.scala 30:36:@44.4]
  wire  _T_17690; // @[Switch.scala 30:53:@46.4]
  wire  valid_0_12; // @[Switch.scala 30:36:@47.4]
  wire  _T_17693; // @[Switch.scala 30:53:@49.4]
  wire  valid_0_13; // @[Switch.scala 30:36:@50.4]
  wire  _T_17696; // @[Switch.scala 30:53:@52.4]
  wire  valid_0_14; // @[Switch.scala 30:36:@53.4]
  wire  _T_17699; // @[Switch.scala 30:53:@55.4]
  wire  valid_0_15; // @[Switch.scala 30:36:@56.4]
  wire  _T_17702; // @[Switch.scala 30:53:@58.4]
  wire  valid_0_16; // @[Switch.scala 30:36:@59.4]
  wire  _T_17705; // @[Switch.scala 30:53:@61.4]
  wire  valid_0_17; // @[Switch.scala 30:36:@62.4]
  wire  _T_17708; // @[Switch.scala 30:53:@64.4]
  wire  valid_0_18; // @[Switch.scala 30:36:@65.4]
  wire  _T_17711; // @[Switch.scala 30:53:@67.4]
  wire  valid_0_19; // @[Switch.scala 30:36:@68.4]
  wire  _T_17714; // @[Switch.scala 30:53:@70.4]
  wire  valid_0_20; // @[Switch.scala 30:36:@71.4]
  wire  _T_17717; // @[Switch.scala 30:53:@73.4]
  wire  valid_0_21; // @[Switch.scala 30:36:@74.4]
  wire  _T_17720; // @[Switch.scala 30:53:@76.4]
  wire  valid_0_22; // @[Switch.scala 30:36:@77.4]
  wire  _T_17723; // @[Switch.scala 30:53:@79.4]
  wire  valid_0_23; // @[Switch.scala 30:36:@80.4]
  wire  _T_17726; // @[Switch.scala 30:53:@82.4]
  wire  valid_0_24; // @[Switch.scala 30:36:@83.4]
  wire  _T_17729; // @[Switch.scala 30:53:@85.4]
  wire  valid_0_25; // @[Switch.scala 30:36:@86.4]
  wire  _T_17732; // @[Switch.scala 30:53:@88.4]
  wire  valid_0_26; // @[Switch.scala 30:36:@89.4]
  wire  _T_17735; // @[Switch.scala 30:53:@91.4]
  wire  valid_0_27; // @[Switch.scala 30:36:@92.4]
  wire  _T_17738; // @[Switch.scala 30:53:@94.4]
  wire  valid_0_28; // @[Switch.scala 30:36:@95.4]
  wire  _T_17741; // @[Switch.scala 30:53:@97.4]
  wire  valid_0_29; // @[Switch.scala 30:36:@98.4]
  wire  _T_17744; // @[Switch.scala 30:53:@100.4]
  wire  valid_0_30; // @[Switch.scala 30:36:@101.4]
  wire  _T_17747; // @[Switch.scala 30:53:@103.4]
  wire  valid_0_31; // @[Switch.scala 30:36:@104.4]
  wire  _T_17750; // @[Switch.scala 30:53:@106.4]
  wire  valid_0_32; // @[Switch.scala 30:36:@107.4]
  wire  _T_17753; // @[Switch.scala 30:53:@109.4]
  wire  valid_0_33; // @[Switch.scala 30:36:@110.4]
  wire  _T_17756; // @[Switch.scala 30:53:@112.4]
  wire  valid_0_34; // @[Switch.scala 30:36:@113.4]
  wire  _T_17759; // @[Switch.scala 30:53:@115.4]
  wire  valid_0_35; // @[Switch.scala 30:36:@116.4]
  wire  _T_17762; // @[Switch.scala 30:53:@118.4]
  wire  valid_0_36; // @[Switch.scala 30:36:@119.4]
  wire  _T_17765; // @[Switch.scala 30:53:@121.4]
  wire  valid_0_37; // @[Switch.scala 30:36:@122.4]
  wire  _T_17768; // @[Switch.scala 30:53:@124.4]
  wire  valid_0_38; // @[Switch.scala 30:36:@125.4]
  wire  _T_17771; // @[Switch.scala 30:53:@127.4]
  wire  valid_0_39; // @[Switch.scala 30:36:@128.4]
  wire  _T_17774; // @[Switch.scala 30:53:@130.4]
  wire  valid_0_40; // @[Switch.scala 30:36:@131.4]
  wire  _T_17777; // @[Switch.scala 30:53:@133.4]
  wire  valid_0_41; // @[Switch.scala 30:36:@134.4]
  wire  _T_17780; // @[Switch.scala 30:53:@136.4]
  wire  valid_0_42; // @[Switch.scala 30:36:@137.4]
  wire  _T_17783; // @[Switch.scala 30:53:@139.4]
  wire  valid_0_43; // @[Switch.scala 30:36:@140.4]
  wire  _T_17786; // @[Switch.scala 30:53:@142.4]
  wire  valid_0_44; // @[Switch.scala 30:36:@143.4]
  wire  _T_17789; // @[Switch.scala 30:53:@145.4]
  wire  valid_0_45; // @[Switch.scala 30:36:@146.4]
  wire  _T_17792; // @[Switch.scala 30:53:@148.4]
  wire  valid_0_46; // @[Switch.scala 30:36:@149.4]
  wire  _T_17795; // @[Switch.scala 30:53:@151.4]
  wire  valid_0_47; // @[Switch.scala 30:36:@152.4]
  wire  _T_17798; // @[Switch.scala 30:53:@154.4]
  wire  valid_0_48; // @[Switch.scala 30:36:@155.4]
  wire  _T_17801; // @[Switch.scala 30:53:@157.4]
  wire  valid_0_49; // @[Switch.scala 30:36:@158.4]
  wire  _T_17804; // @[Switch.scala 30:53:@160.4]
  wire  valid_0_50; // @[Switch.scala 30:36:@161.4]
  wire  _T_17807; // @[Switch.scala 30:53:@163.4]
  wire  valid_0_51; // @[Switch.scala 30:36:@164.4]
  wire  _T_17810; // @[Switch.scala 30:53:@166.4]
  wire  valid_0_52; // @[Switch.scala 30:36:@167.4]
  wire  _T_17813; // @[Switch.scala 30:53:@169.4]
  wire  valid_0_53; // @[Switch.scala 30:36:@170.4]
  wire  _T_17816; // @[Switch.scala 30:53:@172.4]
  wire  valid_0_54; // @[Switch.scala 30:36:@173.4]
  wire  _T_17819; // @[Switch.scala 30:53:@175.4]
  wire  valid_0_55; // @[Switch.scala 30:36:@176.4]
  wire  _T_17822; // @[Switch.scala 30:53:@178.4]
  wire  valid_0_56; // @[Switch.scala 30:36:@179.4]
  wire  _T_17825; // @[Switch.scala 30:53:@181.4]
  wire  valid_0_57; // @[Switch.scala 30:36:@182.4]
  wire  _T_17828; // @[Switch.scala 30:53:@184.4]
  wire  valid_0_58; // @[Switch.scala 30:36:@185.4]
  wire  _T_17831; // @[Switch.scala 30:53:@187.4]
  wire  valid_0_59; // @[Switch.scala 30:36:@188.4]
  wire  _T_17834; // @[Switch.scala 30:53:@190.4]
  wire  valid_0_60; // @[Switch.scala 30:36:@191.4]
  wire  _T_17837; // @[Switch.scala 30:53:@193.4]
  wire  valid_0_61; // @[Switch.scala 30:36:@194.4]
  wire  _T_17840; // @[Switch.scala 30:53:@196.4]
  wire  valid_0_62; // @[Switch.scala 30:36:@197.4]
  wire  _T_17843; // @[Switch.scala 30:53:@199.4]
  wire  valid_0_63; // @[Switch.scala 30:36:@200.4]
  wire [5:0] _T_17909; // @[Mux.scala 31:69:@202.4]
  wire [5:0] _T_17910; // @[Mux.scala 31:69:@203.4]
  wire [5:0] _T_17911; // @[Mux.scala 31:69:@204.4]
  wire [5:0] _T_17912; // @[Mux.scala 31:69:@205.4]
  wire [5:0] _T_17913; // @[Mux.scala 31:69:@206.4]
  wire [5:0] _T_17914; // @[Mux.scala 31:69:@207.4]
  wire [5:0] _T_17915; // @[Mux.scala 31:69:@208.4]
  wire [5:0] _T_17916; // @[Mux.scala 31:69:@209.4]
  wire [5:0] _T_17917; // @[Mux.scala 31:69:@210.4]
  wire [5:0] _T_17918; // @[Mux.scala 31:69:@211.4]
  wire [5:0] _T_17919; // @[Mux.scala 31:69:@212.4]
  wire [5:0] _T_17920; // @[Mux.scala 31:69:@213.4]
  wire [5:0] _T_17921; // @[Mux.scala 31:69:@214.4]
  wire [5:0] _T_17922; // @[Mux.scala 31:69:@215.4]
  wire [5:0] _T_17923; // @[Mux.scala 31:69:@216.4]
  wire [5:0] _T_17924; // @[Mux.scala 31:69:@217.4]
  wire [5:0] _T_17925; // @[Mux.scala 31:69:@218.4]
  wire [5:0] _T_17926; // @[Mux.scala 31:69:@219.4]
  wire [5:0] _T_17927; // @[Mux.scala 31:69:@220.4]
  wire [5:0] _T_17928; // @[Mux.scala 31:69:@221.4]
  wire [5:0] _T_17929; // @[Mux.scala 31:69:@222.4]
  wire [5:0] _T_17930; // @[Mux.scala 31:69:@223.4]
  wire [5:0] _T_17931; // @[Mux.scala 31:69:@224.4]
  wire [5:0] _T_17932; // @[Mux.scala 31:69:@225.4]
  wire [5:0] _T_17933; // @[Mux.scala 31:69:@226.4]
  wire [5:0] _T_17934; // @[Mux.scala 31:69:@227.4]
  wire [5:0] _T_17935; // @[Mux.scala 31:69:@228.4]
  wire [5:0] _T_17936; // @[Mux.scala 31:69:@229.4]
  wire [5:0] _T_17937; // @[Mux.scala 31:69:@230.4]
  wire [5:0] _T_17938; // @[Mux.scala 31:69:@231.4]
  wire [5:0] _T_17939; // @[Mux.scala 31:69:@232.4]
  wire [5:0] _T_17940; // @[Mux.scala 31:69:@233.4]
  wire [5:0] _T_17941; // @[Mux.scala 31:69:@234.4]
  wire [5:0] _T_17942; // @[Mux.scala 31:69:@235.4]
  wire [5:0] _T_17943; // @[Mux.scala 31:69:@236.4]
  wire [5:0] _T_17944; // @[Mux.scala 31:69:@237.4]
  wire [5:0] _T_17945; // @[Mux.scala 31:69:@238.4]
  wire [5:0] _T_17946; // @[Mux.scala 31:69:@239.4]
  wire [5:0] _T_17947; // @[Mux.scala 31:69:@240.4]
  wire [5:0] _T_17948; // @[Mux.scala 31:69:@241.4]
  wire [5:0] _T_17949; // @[Mux.scala 31:69:@242.4]
  wire [5:0] _T_17950; // @[Mux.scala 31:69:@243.4]
  wire [5:0] _T_17951; // @[Mux.scala 31:69:@244.4]
  wire [5:0] _T_17952; // @[Mux.scala 31:69:@245.4]
  wire [5:0] _T_17953; // @[Mux.scala 31:69:@246.4]
  wire [5:0] _T_17954; // @[Mux.scala 31:69:@247.4]
  wire [5:0] _T_17955; // @[Mux.scala 31:69:@248.4]
  wire [5:0] _T_17956; // @[Mux.scala 31:69:@249.4]
  wire [5:0] _T_17957; // @[Mux.scala 31:69:@250.4]
  wire [5:0] _T_17958; // @[Mux.scala 31:69:@251.4]
  wire [5:0] _T_17959; // @[Mux.scala 31:69:@252.4]
  wire [5:0] _T_17960; // @[Mux.scala 31:69:@253.4]
  wire [5:0] _T_17961; // @[Mux.scala 31:69:@254.4]
  wire [5:0] _T_17962; // @[Mux.scala 31:69:@255.4]
  wire [5:0] _T_17963; // @[Mux.scala 31:69:@256.4]
  wire [5:0] _T_17964; // @[Mux.scala 31:69:@257.4]
  wire [5:0] _T_17965; // @[Mux.scala 31:69:@258.4]
  wire [5:0] _T_17966; // @[Mux.scala 31:69:@259.4]
  wire [5:0] _T_17967; // @[Mux.scala 31:69:@260.4]
  wire [5:0] _T_17968; // @[Mux.scala 31:69:@261.4]
  wire [5:0] _T_17969; // @[Mux.scala 31:69:@262.4]
  wire [5:0] _T_17970; // @[Mux.scala 31:69:@263.4]
  wire [5:0] select_0; // @[Mux.scala 31:69:@264.4]
  wire [47:0] _GEN_1; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_2; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_3; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_4; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_5; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_6; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_7; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_8; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_9; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_10; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_11; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_12; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_13; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_14; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_15; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_16; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_17; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_18; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_19; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_20; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_21; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_22; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_23; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_24; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_25; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_26; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_27; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_28; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_29; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_30; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_31; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_32; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_33; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_34; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_35; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_36; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_37; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_38; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_39; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_40; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_41; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_42; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_43; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_44; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_45; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_46; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_47; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_48; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_49; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_50; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_51; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_52; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_53; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_54; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_55; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_56; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_57; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_58; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_59; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_60; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_61; // @[Switch.scala 33:19:@266.4]
  wire [47:0] _GEN_62; // @[Switch.scala 33:19:@266.4]
  wire [7:0] _T_17979; // @[Switch.scala 34:32:@273.4]
  wire [15:0] _T_17987; // @[Switch.scala 34:32:@281.4]
  wire [7:0] _T_17994; // @[Switch.scala 34:32:@288.4]
  wire [31:0] _T_18003; // @[Switch.scala 34:32:@297.4]
  wire [7:0] _T_18010; // @[Switch.scala 34:32:@304.4]
  wire [15:0] _T_18018; // @[Switch.scala 34:32:@312.4]
  wire [7:0] _T_18025; // @[Switch.scala 34:32:@319.4]
  wire [31:0] _T_18034; // @[Switch.scala 34:32:@328.4]
  wire [63:0] _T_18035; // @[Switch.scala 34:32:@329.4]
  wire  _T_18039; // @[Switch.scala 30:53:@332.4]
  wire  valid_1_0; // @[Switch.scala 30:36:@333.4]
  wire  _T_18042; // @[Switch.scala 30:53:@335.4]
  wire  valid_1_1; // @[Switch.scala 30:36:@336.4]
  wire  _T_18045; // @[Switch.scala 30:53:@338.4]
  wire  valid_1_2; // @[Switch.scala 30:36:@339.4]
  wire  _T_18048; // @[Switch.scala 30:53:@341.4]
  wire  valid_1_3; // @[Switch.scala 30:36:@342.4]
  wire  _T_18051; // @[Switch.scala 30:53:@344.4]
  wire  valid_1_4; // @[Switch.scala 30:36:@345.4]
  wire  _T_18054; // @[Switch.scala 30:53:@347.4]
  wire  valid_1_5; // @[Switch.scala 30:36:@348.4]
  wire  _T_18057; // @[Switch.scala 30:53:@350.4]
  wire  valid_1_6; // @[Switch.scala 30:36:@351.4]
  wire  _T_18060; // @[Switch.scala 30:53:@353.4]
  wire  valid_1_7; // @[Switch.scala 30:36:@354.4]
  wire  _T_18063; // @[Switch.scala 30:53:@356.4]
  wire  valid_1_8; // @[Switch.scala 30:36:@357.4]
  wire  _T_18066; // @[Switch.scala 30:53:@359.4]
  wire  valid_1_9; // @[Switch.scala 30:36:@360.4]
  wire  _T_18069; // @[Switch.scala 30:53:@362.4]
  wire  valid_1_10; // @[Switch.scala 30:36:@363.4]
  wire  _T_18072; // @[Switch.scala 30:53:@365.4]
  wire  valid_1_11; // @[Switch.scala 30:36:@366.4]
  wire  _T_18075; // @[Switch.scala 30:53:@368.4]
  wire  valid_1_12; // @[Switch.scala 30:36:@369.4]
  wire  _T_18078; // @[Switch.scala 30:53:@371.4]
  wire  valid_1_13; // @[Switch.scala 30:36:@372.4]
  wire  _T_18081; // @[Switch.scala 30:53:@374.4]
  wire  valid_1_14; // @[Switch.scala 30:36:@375.4]
  wire  _T_18084; // @[Switch.scala 30:53:@377.4]
  wire  valid_1_15; // @[Switch.scala 30:36:@378.4]
  wire  _T_18087; // @[Switch.scala 30:53:@380.4]
  wire  valid_1_16; // @[Switch.scala 30:36:@381.4]
  wire  _T_18090; // @[Switch.scala 30:53:@383.4]
  wire  valid_1_17; // @[Switch.scala 30:36:@384.4]
  wire  _T_18093; // @[Switch.scala 30:53:@386.4]
  wire  valid_1_18; // @[Switch.scala 30:36:@387.4]
  wire  _T_18096; // @[Switch.scala 30:53:@389.4]
  wire  valid_1_19; // @[Switch.scala 30:36:@390.4]
  wire  _T_18099; // @[Switch.scala 30:53:@392.4]
  wire  valid_1_20; // @[Switch.scala 30:36:@393.4]
  wire  _T_18102; // @[Switch.scala 30:53:@395.4]
  wire  valid_1_21; // @[Switch.scala 30:36:@396.4]
  wire  _T_18105; // @[Switch.scala 30:53:@398.4]
  wire  valid_1_22; // @[Switch.scala 30:36:@399.4]
  wire  _T_18108; // @[Switch.scala 30:53:@401.4]
  wire  valid_1_23; // @[Switch.scala 30:36:@402.4]
  wire  _T_18111; // @[Switch.scala 30:53:@404.4]
  wire  valid_1_24; // @[Switch.scala 30:36:@405.4]
  wire  _T_18114; // @[Switch.scala 30:53:@407.4]
  wire  valid_1_25; // @[Switch.scala 30:36:@408.4]
  wire  _T_18117; // @[Switch.scala 30:53:@410.4]
  wire  valid_1_26; // @[Switch.scala 30:36:@411.4]
  wire  _T_18120; // @[Switch.scala 30:53:@413.4]
  wire  valid_1_27; // @[Switch.scala 30:36:@414.4]
  wire  _T_18123; // @[Switch.scala 30:53:@416.4]
  wire  valid_1_28; // @[Switch.scala 30:36:@417.4]
  wire  _T_18126; // @[Switch.scala 30:53:@419.4]
  wire  valid_1_29; // @[Switch.scala 30:36:@420.4]
  wire  _T_18129; // @[Switch.scala 30:53:@422.4]
  wire  valid_1_30; // @[Switch.scala 30:36:@423.4]
  wire  _T_18132; // @[Switch.scala 30:53:@425.4]
  wire  valid_1_31; // @[Switch.scala 30:36:@426.4]
  wire  _T_18135; // @[Switch.scala 30:53:@428.4]
  wire  valid_1_32; // @[Switch.scala 30:36:@429.4]
  wire  _T_18138; // @[Switch.scala 30:53:@431.4]
  wire  valid_1_33; // @[Switch.scala 30:36:@432.4]
  wire  _T_18141; // @[Switch.scala 30:53:@434.4]
  wire  valid_1_34; // @[Switch.scala 30:36:@435.4]
  wire  _T_18144; // @[Switch.scala 30:53:@437.4]
  wire  valid_1_35; // @[Switch.scala 30:36:@438.4]
  wire  _T_18147; // @[Switch.scala 30:53:@440.4]
  wire  valid_1_36; // @[Switch.scala 30:36:@441.4]
  wire  _T_18150; // @[Switch.scala 30:53:@443.4]
  wire  valid_1_37; // @[Switch.scala 30:36:@444.4]
  wire  _T_18153; // @[Switch.scala 30:53:@446.4]
  wire  valid_1_38; // @[Switch.scala 30:36:@447.4]
  wire  _T_18156; // @[Switch.scala 30:53:@449.4]
  wire  valid_1_39; // @[Switch.scala 30:36:@450.4]
  wire  _T_18159; // @[Switch.scala 30:53:@452.4]
  wire  valid_1_40; // @[Switch.scala 30:36:@453.4]
  wire  _T_18162; // @[Switch.scala 30:53:@455.4]
  wire  valid_1_41; // @[Switch.scala 30:36:@456.4]
  wire  _T_18165; // @[Switch.scala 30:53:@458.4]
  wire  valid_1_42; // @[Switch.scala 30:36:@459.4]
  wire  _T_18168; // @[Switch.scala 30:53:@461.4]
  wire  valid_1_43; // @[Switch.scala 30:36:@462.4]
  wire  _T_18171; // @[Switch.scala 30:53:@464.4]
  wire  valid_1_44; // @[Switch.scala 30:36:@465.4]
  wire  _T_18174; // @[Switch.scala 30:53:@467.4]
  wire  valid_1_45; // @[Switch.scala 30:36:@468.4]
  wire  _T_18177; // @[Switch.scala 30:53:@470.4]
  wire  valid_1_46; // @[Switch.scala 30:36:@471.4]
  wire  _T_18180; // @[Switch.scala 30:53:@473.4]
  wire  valid_1_47; // @[Switch.scala 30:36:@474.4]
  wire  _T_18183; // @[Switch.scala 30:53:@476.4]
  wire  valid_1_48; // @[Switch.scala 30:36:@477.4]
  wire  _T_18186; // @[Switch.scala 30:53:@479.4]
  wire  valid_1_49; // @[Switch.scala 30:36:@480.4]
  wire  _T_18189; // @[Switch.scala 30:53:@482.4]
  wire  valid_1_50; // @[Switch.scala 30:36:@483.4]
  wire  _T_18192; // @[Switch.scala 30:53:@485.4]
  wire  valid_1_51; // @[Switch.scala 30:36:@486.4]
  wire  _T_18195; // @[Switch.scala 30:53:@488.4]
  wire  valid_1_52; // @[Switch.scala 30:36:@489.4]
  wire  _T_18198; // @[Switch.scala 30:53:@491.4]
  wire  valid_1_53; // @[Switch.scala 30:36:@492.4]
  wire  _T_18201; // @[Switch.scala 30:53:@494.4]
  wire  valid_1_54; // @[Switch.scala 30:36:@495.4]
  wire  _T_18204; // @[Switch.scala 30:53:@497.4]
  wire  valid_1_55; // @[Switch.scala 30:36:@498.4]
  wire  _T_18207; // @[Switch.scala 30:53:@500.4]
  wire  valid_1_56; // @[Switch.scala 30:36:@501.4]
  wire  _T_18210; // @[Switch.scala 30:53:@503.4]
  wire  valid_1_57; // @[Switch.scala 30:36:@504.4]
  wire  _T_18213; // @[Switch.scala 30:53:@506.4]
  wire  valid_1_58; // @[Switch.scala 30:36:@507.4]
  wire  _T_18216; // @[Switch.scala 30:53:@509.4]
  wire  valid_1_59; // @[Switch.scala 30:36:@510.4]
  wire  _T_18219; // @[Switch.scala 30:53:@512.4]
  wire  valid_1_60; // @[Switch.scala 30:36:@513.4]
  wire  _T_18222; // @[Switch.scala 30:53:@515.4]
  wire  valid_1_61; // @[Switch.scala 30:36:@516.4]
  wire  _T_18225; // @[Switch.scala 30:53:@518.4]
  wire  valid_1_62; // @[Switch.scala 30:36:@519.4]
  wire  _T_18228; // @[Switch.scala 30:53:@521.4]
  wire  valid_1_63; // @[Switch.scala 30:36:@522.4]
  wire [5:0] _T_18294; // @[Mux.scala 31:69:@524.4]
  wire [5:0] _T_18295; // @[Mux.scala 31:69:@525.4]
  wire [5:0] _T_18296; // @[Mux.scala 31:69:@526.4]
  wire [5:0] _T_18297; // @[Mux.scala 31:69:@527.4]
  wire [5:0] _T_18298; // @[Mux.scala 31:69:@528.4]
  wire [5:0] _T_18299; // @[Mux.scala 31:69:@529.4]
  wire [5:0] _T_18300; // @[Mux.scala 31:69:@530.4]
  wire [5:0] _T_18301; // @[Mux.scala 31:69:@531.4]
  wire [5:0] _T_18302; // @[Mux.scala 31:69:@532.4]
  wire [5:0] _T_18303; // @[Mux.scala 31:69:@533.4]
  wire [5:0] _T_18304; // @[Mux.scala 31:69:@534.4]
  wire [5:0] _T_18305; // @[Mux.scala 31:69:@535.4]
  wire [5:0] _T_18306; // @[Mux.scala 31:69:@536.4]
  wire [5:0] _T_18307; // @[Mux.scala 31:69:@537.4]
  wire [5:0] _T_18308; // @[Mux.scala 31:69:@538.4]
  wire [5:0] _T_18309; // @[Mux.scala 31:69:@539.4]
  wire [5:0] _T_18310; // @[Mux.scala 31:69:@540.4]
  wire [5:0] _T_18311; // @[Mux.scala 31:69:@541.4]
  wire [5:0] _T_18312; // @[Mux.scala 31:69:@542.4]
  wire [5:0] _T_18313; // @[Mux.scala 31:69:@543.4]
  wire [5:0] _T_18314; // @[Mux.scala 31:69:@544.4]
  wire [5:0] _T_18315; // @[Mux.scala 31:69:@545.4]
  wire [5:0] _T_18316; // @[Mux.scala 31:69:@546.4]
  wire [5:0] _T_18317; // @[Mux.scala 31:69:@547.4]
  wire [5:0] _T_18318; // @[Mux.scala 31:69:@548.4]
  wire [5:0] _T_18319; // @[Mux.scala 31:69:@549.4]
  wire [5:0] _T_18320; // @[Mux.scala 31:69:@550.4]
  wire [5:0] _T_18321; // @[Mux.scala 31:69:@551.4]
  wire [5:0] _T_18322; // @[Mux.scala 31:69:@552.4]
  wire [5:0] _T_18323; // @[Mux.scala 31:69:@553.4]
  wire [5:0] _T_18324; // @[Mux.scala 31:69:@554.4]
  wire [5:0] _T_18325; // @[Mux.scala 31:69:@555.4]
  wire [5:0] _T_18326; // @[Mux.scala 31:69:@556.4]
  wire [5:0] _T_18327; // @[Mux.scala 31:69:@557.4]
  wire [5:0] _T_18328; // @[Mux.scala 31:69:@558.4]
  wire [5:0] _T_18329; // @[Mux.scala 31:69:@559.4]
  wire [5:0] _T_18330; // @[Mux.scala 31:69:@560.4]
  wire [5:0] _T_18331; // @[Mux.scala 31:69:@561.4]
  wire [5:0] _T_18332; // @[Mux.scala 31:69:@562.4]
  wire [5:0] _T_18333; // @[Mux.scala 31:69:@563.4]
  wire [5:0] _T_18334; // @[Mux.scala 31:69:@564.4]
  wire [5:0] _T_18335; // @[Mux.scala 31:69:@565.4]
  wire [5:0] _T_18336; // @[Mux.scala 31:69:@566.4]
  wire [5:0] _T_18337; // @[Mux.scala 31:69:@567.4]
  wire [5:0] _T_18338; // @[Mux.scala 31:69:@568.4]
  wire [5:0] _T_18339; // @[Mux.scala 31:69:@569.4]
  wire [5:0] _T_18340; // @[Mux.scala 31:69:@570.4]
  wire [5:0] _T_18341; // @[Mux.scala 31:69:@571.4]
  wire [5:0] _T_18342; // @[Mux.scala 31:69:@572.4]
  wire [5:0] _T_18343; // @[Mux.scala 31:69:@573.4]
  wire [5:0] _T_18344; // @[Mux.scala 31:69:@574.4]
  wire [5:0] _T_18345; // @[Mux.scala 31:69:@575.4]
  wire [5:0] _T_18346; // @[Mux.scala 31:69:@576.4]
  wire [5:0] _T_18347; // @[Mux.scala 31:69:@577.4]
  wire [5:0] _T_18348; // @[Mux.scala 31:69:@578.4]
  wire [5:0] _T_18349; // @[Mux.scala 31:69:@579.4]
  wire [5:0] _T_18350; // @[Mux.scala 31:69:@580.4]
  wire [5:0] _T_18351; // @[Mux.scala 31:69:@581.4]
  wire [5:0] _T_18352; // @[Mux.scala 31:69:@582.4]
  wire [5:0] _T_18353; // @[Mux.scala 31:69:@583.4]
  wire [5:0] _T_18354; // @[Mux.scala 31:69:@584.4]
  wire [5:0] _T_18355; // @[Mux.scala 31:69:@585.4]
  wire [5:0] select_1; // @[Mux.scala 31:69:@586.4]
  wire [47:0] _GEN_65; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_66; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_67; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_68; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_69; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_70; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_71; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_72; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_73; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_74; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_75; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_76; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_77; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_78; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_79; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_80; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_81; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_82; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_83; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_84; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_85; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_86; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_87; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_88; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_89; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_90; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_91; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_92; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_93; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_94; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_95; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_96; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_97; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_98; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_99; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_100; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_101; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_102; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_103; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_104; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_105; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_106; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_107; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_108; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_109; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_110; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_111; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_112; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_113; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_114; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_115; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_116; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_117; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_118; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_119; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_120; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_121; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_122; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_123; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_124; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_125; // @[Switch.scala 33:19:@588.4]
  wire [47:0] _GEN_126; // @[Switch.scala 33:19:@588.4]
  wire [7:0] _T_18364; // @[Switch.scala 34:32:@595.4]
  wire [15:0] _T_18372; // @[Switch.scala 34:32:@603.4]
  wire [7:0] _T_18379; // @[Switch.scala 34:32:@610.4]
  wire [31:0] _T_18388; // @[Switch.scala 34:32:@619.4]
  wire [7:0] _T_18395; // @[Switch.scala 34:32:@626.4]
  wire [15:0] _T_18403; // @[Switch.scala 34:32:@634.4]
  wire [7:0] _T_18410; // @[Switch.scala 34:32:@641.4]
  wire [31:0] _T_18419; // @[Switch.scala 34:32:@650.4]
  wire [63:0] _T_18420; // @[Switch.scala 34:32:@651.4]
  wire  _T_18424; // @[Switch.scala 30:53:@654.4]
  wire  valid_2_0; // @[Switch.scala 30:36:@655.4]
  wire  _T_18427; // @[Switch.scala 30:53:@657.4]
  wire  valid_2_1; // @[Switch.scala 30:36:@658.4]
  wire  _T_18430; // @[Switch.scala 30:53:@660.4]
  wire  valid_2_2; // @[Switch.scala 30:36:@661.4]
  wire  _T_18433; // @[Switch.scala 30:53:@663.4]
  wire  valid_2_3; // @[Switch.scala 30:36:@664.4]
  wire  _T_18436; // @[Switch.scala 30:53:@666.4]
  wire  valid_2_4; // @[Switch.scala 30:36:@667.4]
  wire  _T_18439; // @[Switch.scala 30:53:@669.4]
  wire  valid_2_5; // @[Switch.scala 30:36:@670.4]
  wire  _T_18442; // @[Switch.scala 30:53:@672.4]
  wire  valid_2_6; // @[Switch.scala 30:36:@673.4]
  wire  _T_18445; // @[Switch.scala 30:53:@675.4]
  wire  valid_2_7; // @[Switch.scala 30:36:@676.4]
  wire  _T_18448; // @[Switch.scala 30:53:@678.4]
  wire  valid_2_8; // @[Switch.scala 30:36:@679.4]
  wire  _T_18451; // @[Switch.scala 30:53:@681.4]
  wire  valid_2_9; // @[Switch.scala 30:36:@682.4]
  wire  _T_18454; // @[Switch.scala 30:53:@684.4]
  wire  valid_2_10; // @[Switch.scala 30:36:@685.4]
  wire  _T_18457; // @[Switch.scala 30:53:@687.4]
  wire  valid_2_11; // @[Switch.scala 30:36:@688.4]
  wire  _T_18460; // @[Switch.scala 30:53:@690.4]
  wire  valid_2_12; // @[Switch.scala 30:36:@691.4]
  wire  _T_18463; // @[Switch.scala 30:53:@693.4]
  wire  valid_2_13; // @[Switch.scala 30:36:@694.4]
  wire  _T_18466; // @[Switch.scala 30:53:@696.4]
  wire  valid_2_14; // @[Switch.scala 30:36:@697.4]
  wire  _T_18469; // @[Switch.scala 30:53:@699.4]
  wire  valid_2_15; // @[Switch.scala 30:36:@700.4]
  wire  _T_18472; // @[Switch.scala 30:53:@702.4]
  wire  valid_2_16; // @[Switch.scala 30:36:@703.4]
  wire  _T_18475; // @[Switch.scala 30:53:@705.4]
  wire  valid_2_17; // @[Switch.scala 30:36:@706.4]
  wire  _T_18478; // @[Switch.scala 30:53:@708.4]
  wire  valid_2_18; // @[Switch.scala 30:36:@709.4]
  wire  _T_18481; // @[Switch.scala 30:53:@711.4]
  wire  valid_2_19; // @[Switch.scala 30:36:@712.4]
  wire  _T_18484; // @[Switch.scala 30:53:@714.4]
  wire  valid_2_20; // @[Switch.scala 30:36:@715.4]
  wire  _T_18487; // @[Switch.scala 30:53:@717.4]
  wire  valid_2_21; // @[Switch.scala 30:36:@718.4]
  wire  _T_18490; // @[Switch.scala 30:53:@720.4]
  wire  valid_2_22; // @[Switch.scala 30:36:@721.4]
  wire  _T_18493; // @[Switch.scala 30:53:@723.4]
  wire  valid_2_23; // @[Switch.scala 30:36:@724.4]
  wire  _T_18496; // @[Switch.scala 30:53:@726.4]
  wire  valid_2_24; // @[Switch.scala 30:36:@727.4]
  wire  _T_18499; // @[Switch.scala 30:53:@729.4]
  wire  valid_2_25; // @[Switch.scala 30:36:@730.4]
  wire  _T_18502; // @[Switch.scala 30:53:@732.4]
  wire  valid_2_26; // @[Switch.scala 30:36:@733.4]
  wire  _T_18505; // @[Switch.scala 30:53:@735.4]
  wire  valid_2_27; // @[Switch.scala 30:36:@736.4]
  wire  _T_18508; // @[Switch.scala 30:53:@738.4]
  wire  valid_2_28; // @[Switch.scala 30:36:@739.4]
  wire  _T_18511; // @[Switch.scala 30:53:@741.4]
  wire  valid_2_29; // @[Switch.scala 30:36:@742.4]
  wire  _T_18514; // @[Switch.scala 30:53:@744.4]
  wire  valid_2_30; // @[Switch.scala 30:36:@745.4]
  wire  _T_18517; // @[Switch.scala 30:53:@747.4]
  wire  valid_2_31; // @[Switch.scala 30:36:@748.4]
  wire  _T_18520; // @[Switch.scala 30:53:@750.4]
  wire  valid_2_32; // @[Switch.scala 30:36:@751.4]
  wire  _T_18523; // @[Switch.scala 30:53:@753.4]
  wire  valid_2_33; // @[Switch.scala 30:36:@754.4]
  wire  _T_18526; // @[Switch.scala 30:53:@756.4]
  wire  valid_2_34; // @[Switch.scala 30:36:@757.4]
  wire  _T_18529; // @[Switch.scala 30:53:@759.4]
  wire  valid_2_35; // @[Switch.scala 30:36:@760.4]
  wire  _T_18532; // @[Switch.scala 30:53:@762.4]
  wire  valid_2_36; // @[Switch.scala 30:36:@763.4]
  wire  _T_18535; // @[Switch.scala 30:53:@765.4]
  wire  valid_2_37; // @[Switch.scala 30:36:@766.4]
  wire  _T_18538; // @[Switch.scala 30:53:@768.4]
  wire  valid_2_38; // @[Switch.scala 30:36:@769.4]
  wire  _T_18541; // @[Switch.scala 30:53:@771.4]
  wire  valid_2_39; // @[Switch.scala 30:36:@772.4]
  wire  _T_18544; // @[Switch.scala 30:53:@774.4]
  wire  valid_2_40; // @[Switch.scala 30:36:@775.4]
  wire  _T_18547; // @[Switch.scala 30:53:@777.4]
  wire  valid_2_41; // @[Switch.scala 30:36:@778.4]
  wire  _T_18550; // @[Switch.scala 30:53:@780.4]
  wire  valid_2_42; // @[Switch.scala 30:36:@781.4]
  wire  _T_18553; // @[Switch.scala 30:53:@783.4]
  wire  valid_2_43; // @[Switch.scala 30:36:@784.4]
  wire  _T_18556; // @[Switch.scala 30:53:@786.4]
  wire  valid_2_44; // @[Switch.scala 30:36:@787.4]
  wire  _T_18559; // @[Switch.scala 30:53:@789.4]
  wire  valid_2_45; // @[Switch.scala 30:36:@790.4]
  wire  _T_18562; // @[Switch.scala 30:53:@792.4]
  wire  valid_2_46; // @[Switch.scala 30:36:@793.4]
  wire  _T_18565; // @[Switch.scala 30:53:@795.4]
  wire  valid_2_47; // @[Switch.scala 30:36:@796.4]
  wire  _T_18568; // @[Switch.scala 30:53:@798.4]
  wire  valid_2_48; // @[Switch.scala 30:36:@799.4]
  wire  _T_18571; // @[Switch.scala 30:53:@801.4]
  wire  valid_2_49; // @[Switch.scala 30:36:@802.4]
  wire  _T_18574; // @[Switch.scala 30:53:@804.4]
  wire  valid_2_50; // @[Switch.scala 30:36:@805.4]
  wire  _T_18577; // @[Switch.scala 30:53:@807.4]
  wire  valid_2_51; // @[Switch.scala 30:36:@808.4]
  wire  _T_18580; // @[Switch.scala 30:53:@810.4]
  wire  valid_2_52; // @[Switch.scala 30:36:@811.4]
  wire  _T_18583; // @[Switch.scala 30:53:@813.4]
  wire  valid_2_53; // @[Switch.scala 30:36:@814.4]
  wire  _T_18586; // @[Switch.scala 30:53:@816.4]
  wire  valid_2_54; // @[Switch.scala 30:36:@817.4]
  wire  _T_18589; // @[Switch.scala 30:53:@819.4]
  wire  valid_2_55; // @[Switch.scala 30:36:@820.4]
  wire  _T_18592; // @[Switch.scala 30:53:@822.4]
  wire  valid_2_56; // @[Switch.scala 30:36:@823.4]
  wire  _T_18595; // @[Switch.scala 30:53:@825.4]
  wire  valid_2_57; // @[Switch.scala 30:36:@826.4]
  wire  _T_18598; // @[Switch.scala 30:53:@828.4]
  wire  valid_2_58; // @[Switch.scala 30:36:@829.4]
  wire  _T_18601; // @[Switch.scala 30:53:@831.4]
  wire  valid_2_59; // @[Switch.scala 30:36:@832.4]
  wire  _T_18604; // @[Switch.scala 30:53:@834.4]
  wire  valid_2_60; // @[Switch.scala 30:36:@835.4]
  wire  _T_18607; // @[Switch.scala 30:53:@837.4]
  wire  valid_2_61; // @[Switch.scala 30:36:@838.4]
  wire  _T_18610; // @[Switch.scala 30:53:@840.4]
  wire  valid_2_62; // @[Switch.scala 30:36:@841.4]
  wire  _T_18613; // @[Switch.scala 30:53:@843.4]
  wire  valid_2_63; // @[Switch.scala 30:36:@844.4]
  wire [5:0] _T_18679; // @[Mux.scala 31:69:@846.4]
  wire [5:0] _T_18680; // @[Mux.scala 31:69:@847.4]
  wire [5:0] _T_18681; // @[Mux.scala 31:69:@848.4]
  wire [5:0] _T_18682; // @[Mux.scala 31:69:@849.4]
  wire [5:0] _T_18683; // @[Mux.scala 31:69:@850.4]
  wire [5:0] _T_18684; // @[Mux.scala 31:69:@851.4]
  wire [5:0] _T_18685; // @[Mux.scala 31:69:@852.4]
  wire [5:0] _T_18686; // @[Mux.scala 31:69:@853.4]
  wire [5:0] _T_18687; // @[Mux.scala 31:69:@854.4]
  wire [5:0] _T_18688; // @[Mux.scala 31:69:@855.4]
  wire [5:0] _T_18689; // @[Mux.scala 31:69:@856.4]
  wire [5:0] _T_18690; // @[Mux.scala 31:69:@857.4]
  wire [5:0] _T_18691; // @[Mux.scala 31:69:@858.4]
  wire [5:0] _T_18692; // @[Mux.scala 31:69:@859.4]
  wire [5:0] _T_18693; // @[Mux.scala 31:69:@860.4]
  wire [5:0] _T_18694; // @[Mux.scala 31:69:@861.4]
  wire [5:0] _T_18695; // @[Mux.scala 31:69:@862.4]
  wire [5:0] _T_18696; // @[Mux.scala 31:69:@863.4]
  wire [5:0] _T_18697; // @[Mux.scala 31:69:@864.4]
  wire [5:0] _T_18698; // @[Mux.scala 31:69:@865.4]
  wire [5:0] _T_18699; // @[Mux.scala 31:69:@866.4]
  wire [5:0] _T_18700; // @[Mux.scala 31:69:@867.4]
  wire [5:0] _T_18701; // @[Mux.scala 31:69:@868.4]
  wire [5:0] _T_18702; // @[Mux.scala 31:69:@869.4]
  wire [5:0] _T_18703; // @[Mux.scala 31:69:@870.4]
  wire [5:0] _T_18704; // @[Mux.scala 31:69:@871.4]
  wire [5:0] _T_18705; // @[Mux.scala 31:69:@872.4]
  wire [5:0] _T_18706; // @[Mux.scala 31:69:@873.4]
  wire [5:0] _T_18707; // @[Mux.scala 31:69:@874.4]
  wire [5:0] _T_18708; // @[Mux.scala 31:69:@875.4]
  wire [5:0] _T_18709; // @[Mux.scala 31:69:@876.4]
  wire [5:0] _T_18710; // @[Mux.scala 31:69:@877.4]
  wire [5:0] _T_18711; // @[Mux.scala 31:69:@878.4]
  wire [5:0] _T_18712; // @[Mux.scala 31:69:@879.4]
  wire [5:0] _T_18713; // @[Mux.scala 31:69:@880.4]
  wire [5:0] _T_18714; // @[Mux.scala 31:69:@881.4]
  wire [5:0] _T_18715; // @[Mux.scala 31:69:@882.4]
  wire [5:0] _T_18716; // @[Mux.scala 31:69:@883.4]
  wire [5:0] _T_18717; // @[Mux.scala 31:69:@884.4]
  wire [5:0] _T_18718; // @[Mux.scala 31:69:@885.4]
  wire [5:0] _T_18719; // @[Mux.scala 31:69:@886.4]
  wire [5:0] _T_18720; // @[Mux.scala 31:69:@887.4]
  wire [5:0] _T_18721; // @[Mux.scala 31:69:@888.4]
  wire [5:0] _T_18722; // @[Mux.scala 31:69:@889.4]
  wire [5:0] _T_18723; // @[Mux.scala 31:69:@890.4]
  wire [5:0] _T_18724; // @[Mux.scala 31:69:@891.4]
  wire [5:0] _T_18725; // @[Mux.scala 31:69:@892.4]
  wire [5:0] _T_18726; // @[Mux.scala 31:69:@893.4]
  wire [5:0] _T_18727; // @[Mux.scala 31:69:@894.4]
  wire [5:0] _T_18728; // @[Mux.scala 31:69:@895.4]
  wire [5:0] _T_18729; // @[Mux.scala 31:69:@896.4]
  wire [5:0] _T_18730; // @[Mux.scala 31:69:@897.4]
  wire [5:0] _T_18731; // @[Mux.scala 31:69:@898.4]
  wire [5:0] _T_18732; // @[Mux.scala 31:69:@899.4]
  wire [5:0] _T_18733; // @[Mux.scala 31:69:@900.4]
  wire [5:0] _T_18734; // @[Mux.scala 31:69:@901.4]
  wire [5:0] _T_18735; // @[Mux.scala 31:69:@902.4]
  wire [5:0] _T_18736; // @[Mux.scala 31:69:@903.4]
  wire [5:0] _T_18737; // @[Mux.scala 31:69:@904.4]
  wire [5:0] _T_18738; // @[Mux.scala 31:69:@905.4]
  wire [5:0] _T_18739; // @[Mux.scala 31:69:@906.4]
  wire [5:0] _T_18740; // @[Mux.scala 31:69:@907.4]
  wire [5:0] select_2; // @[Mux.scala 31:69:@908.4]
  wire [47:0] _GEN_129; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_130; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_131; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_132; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_133; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_134; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_135; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_136; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_137; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_138; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_139; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_140; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_141; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_142; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_143; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_144; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_145; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_146; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_147; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_148; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_149; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_150; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_151; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_152; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_153; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_154; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_155; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_156; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_157; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_158; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_159; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_160; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_161; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_162; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_163; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_164; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_165; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_166; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_167; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_168; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_169; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_170; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_171; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_172; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_173; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_174; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_175; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_176; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_177; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_178; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_179; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_180; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_181; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_182; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_183; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_184; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_185; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_186; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_187; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_188; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_189; // @[Switch.scala 33:19:@910.4]
  wire [47:0] _GEN_190; // @[Switch.scala 33:19:@910.4]
  wire [7:0] _T_18749; // @[Switch.scala 34:32:@917.4]
  wire [15:0] _T_18757; // @[Switch.scala 34:32:@925.4]
  wire [7:0] _T_18764; // @[Switch.scala 34:32:@932.4]
  wire [31:0] _T_18773; // @[Switch.scala 34:32:@941.4]
  wire [7:0] _T_18780; // @[Switch.scala 34:32:@948.4]
  wire [15:0] _T_18788; // @[Switch.scala 34:32:@956.4]
  wire [7:0] _T_18795; // @[Switch.scala 34:32:@963.4]
  wire [31:0] _T_18804; // @[Switch.scala 34:32:@972.4]
  wire [63:0] _T_18805; // @[Switch.scala 34:32:@973.4]
  wire  _T_18809; // @[Switch.scala 30:53:@976.4]
  wire  valid_3_0; // @[Switch.scala 30:36:@977.4]
  wire  _T_18812; // @[Switch.scala 30:53:@979.4]
  wire  valid_3_1; // @[Switch.scala 30:36:@980.4]
  wire  _T_18815; // @[Switch.scala 30:53:@982.4]
  wire  valid_3_2; // @[Switch.scala 30:36:@983.4]
  wire  _T_18818; // @[Switch.scala 30:53:@985.4]
  wire  valid_3_3; // @[Switch.scala 30:36:@986.4]
  wire  _T_18821; // @[Switch.scala 30:53:@988.4]
  wire  valid_3_4; // @[Switch.scala 30:36:@989.4]
  wire  _T_18824; // @[Switch.scala 30:53:@991.4]
  wire  valid_3_5; // @[Switch.scala 30:36:@992.4]
  wire  _T_18827; // @[Switch.scala 30:53:@994.4]
  wire  valid_3_6; // @[Switch.scala 30:36:@995.4]
  wire  _T_18830; // @[Switch.scala 30:53:@997.4]
  wire  valid_3_7; // @[Switch.scala 30:36:@998.4]
  wire  _T_18833; // @[Switch.scala 30:53:@1000.4]
  wire  valid_3_8; // @[Switch.scala 30:36:@1001.4]
  wire  _T_18836; // @[Switch.scala 30:53:@1003.4]
  wire  valid_3_9; // @[Switch.scala 30:36:@1004.4]
  wire  _T_18839; // @[Switch.scala 30:53:@1006.4]
  wire  valid_3_10; // @[Switch.scala 30:36:@1007.4]
  wire  _T_18842; // @[Switch.scala 30:53:@1009.4]
  wire  valid_3_11; // @[Switch.scala 30:36:@1010.4]
  wire  _T_18845; // @[Switch.scala 30:53:@1012.4]
  wire  valid_3_12; // @[Switch.scala 30:36:@1013.4]
  wire  _T_18848; // @[Switch.scala 30:53:@1015.4]
  wire  valid_3_13; // @[Switch.scala 30:36:@1016.4]
  wire  _T_18851; // @[Switch.scala 30:53:@1018.4]
  wire  valid_3_14; // @[Switch.scala 30:36:@1019.4]
  wire  _T_18854; // @[Switch.scala 30:53:@1021.4]
  wire  valid_3_15; // @[Switch.scala 30:36:@1022.4]
  wire  _T_18857; // @[Switch.scala 30:53:@1024.4]
  wire  valid_3_16; // @[Switch.scala 30:36:@1025.4]
  wire  _T_18860; // @[Switch.scala 30:53:@1027.4]
  wire  valid_3_17; // @[Switch.scala 30:36:@1028.4]
  wire  _T_18863; // @[Switch.scala 30:53:@1030.4]
  wire  valid_3_18; // @[Switch.scala 30:36:@1031.4]
  wire  _T_18866; // @[Switch.scala 30:53:@1033.4]
  wire  valid_3_19; // @[Switch.scala 30:36:@1034.4]
  wire  _T_18869; // @[Switch.scala 30:53:@1036.4]
  wire  valid_3_20; // @[Switch.scala 30:36:@1037.4]
  wire  _T_18872; // @[Switch.scala 30:53:@1039.4]
  wire  valid_3_21; // @[Switch.scala 30:36:@1040.4]
  wire  _T_18875; // @[Switch.scala 30:53:@1042.4]
  wire  valid_3_22; // @[Switch.scala 30:36:@1043.4]
  wire  _T_18878; // @[Switch.scala 30:53:@1045.4]
  wire  valid_3_23; // @[Switch.scala 30:36:@1046.4]
  wire  _T_18881; // @[Switch.scala 30:53:@1048.4]
  wire  valid_3_24; // @[Switch.scala 30:36:@1049.4]
  wire  _T_18884; // @[Switch.scala 30:53:@1051.4]
  wire  valid_3_25; // @[Switch.scala 30:36:@1052.4]
  wire  _T_18887; // @[Switch.scala 30:53:@1054.4]
  wire  valid_3_26; // @[Switch.scala 30:36:@1055.4]
  wire  _T_18890; // @[Switch.scala 30:53:@1057.4]
  wire  valid_3_27; // @[Switch.scala 30:36:@1058.4]
  wire  _T_18893; // @[Switch.scala 30:53:@1060.4]
  wire  valid_3_28; // @[Switch.scala 30:36:@1061.4]
  wire  _T_18896; // @[Switch.scala 30:53:@1063.4]
  wire  valid_3_29; // @[Switch.scala 30:36:@1064.4]
  wire  _T_18899; // @[Switch.scala 30:53:@1066.4]
  wire  valid_3_30; // @[Switch.scala 30:36:@1067.4]
  wire  _T_18902; // @[Switch.scala 30:53:@1069.4]
  wire  valid_3_31; // @[Switch.scala 30:36:@1070.4]
  wire  _T_18905; // @[Switch.scala 30:53:@1072.4]
  wire  valid_3_32; // @[Switch.scala 30:36:@1073.4]
  wire  _T_18908; // @[Switch.scala 30:53:@1075.4]
  wire  valid_3_33; // @[Switch.scala 30:36:@1076.4]
  wire  _T_18911; // @[Switch.scala 30:53:@1078.4]
  wire  valid_3_34; // @[Switch.scala 30:36:@1079.4]
  wire  _T_18914; // @[Switch.scala 30:53:@1081.4]
  wire  valid_3_35; // @[Switch.scala 30:36:@1082.4]
  wire  _T_18917; // @[Switch.scala 30:53:@1084.4]
  wire  valid_3_36; // @[Switch.scala 30:36:@1085.4]
  wire  _T_18920; // @[Switch.scala 30:53:@1087.4]
  wire  valid_3_37; // @[Switch.scala 30:36:@1088.4]
  wire  _T_18923; // @[Switch.scala 30:53:@1090.4]
  wire  valid_3_38; // @[Switch.scala 30:36:@1091.4]
  wire  _T_18926; // @[Switch.scala 30:53:@1093.4]
  wire  valid_3_39; // @[Switch.scala 30:36:@1094.4]
  wire  _T_18929; // @[Switch.scala 30:53:@1096.4]
  wire  valid_3_40; // @[Switch.scala 30:36:@1097.4]
  wire  _T_18932; // @[Switch.scala 30:53:@1099.4]
  wire  valid_3_41; // @[Switch.scala 30:36:@1100.4]
  wire  _T_18935; // @[Switch.scala 30:53:@1102.4]
  wire  valid_3_42; // @[Switch.scala 30:36:@1103.4]
  wire  _T_18938; // @[Switch.scala 30:53:@1105.4]
  wire  valid_3_43; // @[Switch.scala 30:36:@1106.4]
  wire  _T_18941; // @[Switch.scala 30:53:@1108.4]
  wire  valid_3_44; // @[Switch.scala 30:36:@1109.4]
  wire  _T_18944; // @[Switch.scala 30:53:@1111.4]
  wire  valid_3_45; // @[Switch.scala 30:36:@1112.4]
  wire  _T_18947; // @[Switch.scala 30:53:@1114.4]
  wire  valid_3_46; // @[Switch.scala 30:36:@1115.4]
  wire  _T_18950; // @[Switch.scala 30:53:@1117.4]
  wire  valid_3_47; // @[Switch.scala 30:36:@1118.4]
  wire  _T_18953; // @[Switch.scala 30:53:@1120.4]
  wire  valid_3_48; // @[Switch.scala 30:36:@1121.4]
  wire  _T_18956; // @[Switch.scala 30:53:@1123.4]
  wire  valid_3_49; // @[Switch.scala 30:36:@1124.4]
  wire  _T_18959; // @[Switch.scala 30:53:@1126.4]
  wire  valid_3_50; // @[Switch.scala 30:36:@1127.4]
  wire  _T_18962; // @[Switch.scala 30:53:@1129.4]
  wire  valid_3_51; // @[Switch.scala 30:36:@1130.4]
  wire  _T_18965; // @[Switch.scala 30:53:@1132.4]
  wire  valid_3_52; // @[Switch.scala 30:36:@1133.4]
  wire  _T_18968; // @[Switch.scala 30:53:@1135.4]
  wire  valid_3_53; // @[Switch.scala 30:36:@1136.4]
  wire  _T_18971; // @[Switch.scala 30:53:@1138.4]
  wire  valid_3_54; // @[Switch.scala 30:36:@1139.4]
  wire  _T_18974; // @[Switch.scala 30:53:@1141.4]
  wire  valid_3_55; // @[Switch.scala 30:36:@1142.4]
  wire  _T_18977; // @[Switch.scala 30:53:@1144.4]
  wire  valid_3_56; // @[Switch.scala 30:36:@1145.4]
  wire  _T_18980; // @[Switch.scala 30:53:@1147.4]
  wire  valid_3_57; // @[Switch.scala 30:36:@1148.4]
  wire  _T_18983; // @[Switch.scala 30:53:@1150.4]
  wire  valid_3_58; // @[Switch.scala 30:36:@1151.4]
  wire  _T_18986; // @[Switch.scala 30:53:@1153.4]
  wire  valid_3_59; // @[Switch.scala 30:36:@1154.4]
  wire  _T_18989; // @[Switch.scala 30:53:@1156.4]
  wire  valid_3_60; // @[Switch.scala 30:36:@1157.4]
  wire  _T_18992; // @[Switch.scala 30:53:@1159.4]
  wire  valid_3_61; // @[Switch.scala 30:36:@1160.4]
  wire  _T_18995; // @[Switch.scala 30:53:@1162.4]
  wire  valid_3_62; // @[Switch.scala 30:36:@1163.4]
  wire  _T_18998; // @[Switch.scala 30:53:@1165.4]
  wire  valid_3_63; // @[Switch.scala 30:36:@1166.4]
  wire [5:0] _T_19064; // @[Mux.scala 31:69:@1168.4]
  wire [5:0] _T_19065; // @[Mux.scala 31:69:@1169.4]
  wire [5:0] _T_19066; // @[Mux.scala 31:69:@1170.4]
  wire [5:0] _T_19067; // @[Mux.scala 31:69:@1171.4]
  wire [5:0] _T_19068; // @[Mux.scala 31:69:@1172.4]
  wire [5:0] _T_19069; // @[Mux.scala 31:69:@1173.4]
  wire [5:0] _T_19070; // @[Mux.scala 31:69:@1174.4]
  wire [5:0] _T_19071; // @[Mux.scala 31:69:@1175.4]
  wire [5:0] _T_19072; // @[Mux.scala 31:69:@1176.4]
  wire [5:0] _T_19073; // @[Mux.scala 31:69:@1177.4]
  wire [5:0] _T_19074; // @[Mux.scala 31:69:@1178.4]
  wire [5:0] _T_19075; // @[Mux.scala 31:69:@1179.4]
  wire [5:0] _T_19076; // @[Mux.scala 31:69:@1180.4]
  wire [5:0] _T_19077; // @[Mux.scala 31:69:@1181.4]
  wire [5:0] _T_19078; // @[Mux.scala 31:69:@1182.4]
  wire [5:0] _T_19079; // @[Mux.scala 31:69:@1183.4]
  wire [5:0] _T_19080; // @[Mux.scala 31:69:@1184.4]
  wire [5:0] _T_19081; // @[Mux.scala 31:69:@1185.4]
  wire [5:0] _T_19082; // @[Mux.scala 31:69:@1186.4]
  wire [5:0] _T_19083; // @[Mux.scala 31:69:@1187.4]
  wire [5:0] _T_19084; // @[Mux.scala 31:69:@1188.4]
  wire [5:0] _T_19085; // @[Mux.scala 31:69:@1189.4]
  wire [5:0] _T_19086; // @[Mux.scala 31:69:@1190.4]
  wire [5:0] _T_19087; // @[Mux.scala 31:69:@1191.4]
  wire [5:0] _T_19088; // @[Mux.scala 31:69:@1192.4]
  wire [5:0] _T_19089; // @[Mux.scala 31:69:@1193.4]
  wire [5:0] _T_19090; // @[Mux.scala 31:69:@1194.4]
  wire [5:0] _T_19091; // @[Mux.scala 31:69:@1195.4]
  wire [5:0] _T_19092; // @[Mux.scala 31:69:@1196.4]
  wire [5:0] _T_19093; // @[Mux.scala 31:69:@1197.4]
  wire [5:0] _T_19094; // @[Mux.scala 31:69:@1198.4]
  wire [5:0] _T_19095; // @[Mux.scala 31:69:@1199.4]
  wire [5:0] _T_19096; // @[Mux.scala 31:69:@1200.4]
  wire [5:0] _T_19097; // @[Mux.scala 31:69:@1201.4]
  wire [5:0] _T_19098; // @[Mux.scala 31:69:@1202.4]
  wire [5:0] _T_19099; // @[Mux.scala 31:69:@1203.4]
  wire [5:0] _T_19100; // @[Mux.scala 31:69:@1204.4]
  wire [5:0] _T_19101; // @[Mux.scala 31:69:@1205.4]
  wire [5:0] _T_19102; // @[Mux.scala 31:69:@1206.4]
  wire [5:0] _T_19103; // @[Mux.scala 31:69:@1207.4]
  wire [5:0] _T_19104; // @[Mux.scala 31:69:@1208.4]
  wire [5:0] _T_19105; // @[Mux.scala 31:69:@1209.4]
  wire [5:0] _T_19106; // @[Mux.scala 31:69:@1210.4]
  wire [5:0] _T_19107; // @[Mux.scala 31:69:@1211.4]
  wire [5:0] _T_19108; // @[Mux.scala 31:69:@1212.4]
  wire [5:0] _T_19109; // @[Mux.scala 31:69:@1213.4]
  wire [5:0] _T_19110; // @[Mux.scala 31:69:@1214.4]
  wire [5:0] _T_19111; // @[Mux.scala 31:69:@1215.4]
  wire [5:0] _T_19112; // @[Mux.scala 31:69:@1216.4]
  wire [5:0] _T_19113; // @[Mux.scala 31:69:@1217.4]
  wire [5:0] _T_19114; // @[Mux.scala 31:69:@1218.4]
  wire [5:0] _T_19115; // @[Mux.scala 31:69:@1219.4]
  wire [5:0] _T_19116; // @[Mux.scala 31:69:@1220.4]
  wire [5:0] _T_19117; // @[Mux.scala 31:69:@1221.4]
  wire [5:0] _T_19118; // @[Mux.scala 31:69:@1222.4]
  wire [5:0] _T_19119; // @[Mux.scala 31:69:@1223.4]
  wire [5:0] _T_19120; // @[Mux.scala 31:69:@1224.4]
  wire [5:0] _T_19121; // @[Mux.scala 31:69:@1225.4]
  wire [5:0] _T_19122; // @[Mux.scala 31:69:@1226.4]
  wire [5:0] _T_19123; // @[Mux.scala 31:69:@1227.4]
  wire [5:0] _T_19124; // @[Mux.scala 31:69:@1228.4]
  wire [5:0] _T_19125; // @[Mux.scala 31:69:@1229.4]
  wire [5:0] select_3; // @[Mux.scala 31:69:@1230.4]
  wire [47:0] _GEN_193; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_194; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_195; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_196; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_197; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_198; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_199; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_200; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_201; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_202; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_203; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_204; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_205; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_206; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_207; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_208; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_209; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_210; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_211; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_212; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_213; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_214; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_215; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_216; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_217; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_218; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_219; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_220; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_221; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_222; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_223; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_224; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_225; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_226; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_227; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_228; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_229; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_230; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_231; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_232; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_233; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_234; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_235; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_236; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_237; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_238; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_239; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_240; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_241; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_242; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_243; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_244; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_245; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_246; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_247; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_248; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_249; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_250; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_251; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_252; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_253; // @[Switch.scala 33:19:@1232.4]
  wire [47:0] _GEN_254; // @[Switch.scala 33:19:@1232.4]
  wire [7:0] _T_19134; // @[Switch.scala 34:32:@1239.4]
  wire [15:0] _T_19142; // @[Switch.scala 34:32:@1247.4]
  wire [7:0] _T_19149; // @[Switch.scala 34:32:@1254.4]
  wire [31:0] _T_19158; // @[Switch.scala 34:32:@1263.4]
  wire [7:0] _T_19165; // @[Switch.scala 34:32:@1270.4]
  wire [15:0] _T_19173; // @[Switch.scala 34:32:@1278.4]
  wire [7:0] _T_19180; // @[Switch.scala 34:32:@1285.4]
  wire [31:0] _T_19189; // @[Switch.scala 34:32:@1294.4]
  wire [63:0] _T_19190; // @[Switch.scala 34:32:@1295.4]
  wire  _T_19194; // @[Switch.scala 30:53:@1298.4]
  wire  valid_4_0; // @[Switch.scala 30:36:@1299.4]
  wire  _T_19197; // @[Switch.scala 30:53:@1301.4]
  wire  valid_4_1; // @[Switch.scala 30:36:@1302.4]
  wire  _T_19200; // @[Switch.scala 30:53:@1304.4]
  wire  valid_4_2; // @[Switch.scala 30:36:@1305.4]
  wire  _T_19203; // @[Switch.scala 30:53:@1307.4]
  wire  valid_4_3; // @[Switch.scala 30:36:@1308.4]
  wire  _T_19206; // @[Switch.scala 30:53:@1310.4]
  wire  valid_4_4; // @[Switch.scala 30:36:@1311.4]
  wire  _T_19209; // @[Switch.scala 30:53:@1313.4]
  wire  valid_4_5; // @[Switch.scala 30:36:@1314.4]
  wire  _T_19212; // @[Switch.scala 30:53:@1316.4]
  wire  valid_4_6; // @[Switch.scala 30:36:@1317.4]
  wire  _T_19215; // @[Switch.scala 30:53:@1319.4]
  wire  valid_4_7; // @[Switch.scala 30:36:@1320.4]
  wire  _T_19218; // @[Switch.scala 30:53:@1322.4]
  wire  valid_4_8; // @[Switch.scala 30:36:@1323.4]
  wire  _T_19221; // @[Switch.scala 30:53:@1325.4]
  wire  valid_4_9; // @[Switch.scala 30:36:@1326.4]
  wire  _T_19224; // @[Switch.scala 30:53:@1328.4]
  wire  valid_4_10; // @[Switch.scala 30:36:@1329.4]
  wire  _T_19227; // @[Switch.scala 30:53:@1331.4]
  wire  valid_4_11; // @[Switch.scala 30:36:@1332.4]
  wire  _T_19230; // @[Switch.scala 30:53:@1334.4]
  wire  valid_4_12; // @[Switch.scala 30:36:@1335.4]
  wire  _T_19233; // @[Switch.scala 30:53:@1337.4]
  wire  valid_4_13; // @[Switch.scala 30:36:@1338.4]
  wire  _T_19236; // @[Switch.scala 30:53:@1340.4]
  wire  valid_4_14; // @[Switch.scala 30:36:@1341.4]
  wire  _T_19239; // @[Switch.scala 30:53:@1343.4]
  wire  valid_4_15; // @[Switch.scala 30:36:@1344.4]
  wire  _T_19242; // @[Switch.scala 30:53:@1346.4]
  wire  valid_4_16; // @[Switch.scala 30:36:@1347.4]
  wire  _T_19245; // @[Switch.scala 30:53:@1349.4]
  wire  valid_4_17; // @[Switch.scala 30:36:@1350.4]
  wire  _T_19248; // @[Switch.scala 30:53:@1352.4]
  wire  valid_4_18; // @[Switch.scala 30:36:@1353.4]
  wire  _T_19251; // @[Switch.scala 30:53:@1355.4]
  wire  valid_4_19; // @[Switch.scala 30:36:@1356.4]
  wire  _T_19254; // @[Switch.scala 30:53:@1358.4]
  wire  valid_4_20; // @[Switch.scala 30:36:@1359.4]
  wire  _T_19257; // @[Switch.scala 30:53:@1361.4]
  wire  valid_4_21; // @[Switch.scala 30:36:@1362.4]
  wire  _T_19260; // @[Switch.scala 30:53:@1364.4]
  wire  valid_4_22; // @[Switch.scala 30:36:@1365.4]
  wire  _T_19263; // @[Switch.scala 30:53:@1367.4]
  wire  valid_4_23; // @[Switch.scala 30:36:@1368.4]
  wire  _T_19266; // @[Switch.scala 30:53:@1370.4]
  wire  valid_4_24; // @[Switch.scala 30:36:@1371.4]
  wire  _T_19269; // @[Switch.scala 30:53:@1373.4]
  wire  valid_4_25; // @[Switch.scala 30:36:@1374.4]
  wire  _T_19272; // @[Switch.scala 30:53:@1376.4]
  wire  valid_4_26; // @[Switch.scala 30:36:@1377.4]
  wire  _T_19275; // @[Switch.scala 30:53:@1379.4]
  wire  valid_4_27; // @[Switch.scala 30:36:@1380.4]
  wire  _T_19278; // @[Switch.scala 30:53:@1382.4]
  wire  valid_4_28; // @[Switch.scala 30:36:@1383.4]
  wire  _T_19281; // @[Switch.scala 30:53:@1385.4]
  wire  valid_4_29; // @[Switch.scala 30:36:@1386.4]
  wire  _T_19284; // @[Switch.scala 30:53:@1388.4]
  wire  valid_4_30; // @[Switch.scala 30:36:@1389.4]
  wire  _T_19287; // @[Switch.scala 30:53:@1391.4]
  wire  valid_4_31; // @[Switch.scala 30:36:@1392.4]
  wire  _T_19290; // @[Switch.scala 30:53:@1394.4]
  wire  valid_4_32; // @[Switch.scala 30:36:@1395.4]
  wire  _T_19293; // @[Switch.scala 30:53:@1397.4]
  wire  valid_4_33; // @[Switch.scala 30:36:@1398.4]
  wire  _T_19296; // @[Switch.scala 30:53:@1400.4]
  wire  valid_4_34; // @[Switch.scala 30:36:@1401.4]
  wire  _T_19299; // @[Switch.scala 30:53:@1403.4]
  wire  valid_4_35; // @[Switch.scala 30:36:@1404.4]
  wire  _T_19302; // @[Switch.scala 30:53:@1406.4]
  wire  valid_4_36; // @[Switch.scala 30:36:@1407.4]
  wire  _T_19305; // @[Switch.scala 30:53:@1409.4]
  wire  valid_4_37; // @[Switch.scala 30:36:@1410.4]
  wire  _T_19308; // @[Switch.scala 30:53:@1412.4]
  wire  valid_4_38; // @[Switch.scala 30:36:@1413.4]
  wire  _T_19311; // @[Switch.scala 30:53:@1415.4]
  wire  valid_4_39; // @[Switch.scala 30:36:@1416.4]
  wire  _T_19314; // @[Switch.scala 30:53:@1418.4]
  wire  valid_4_40; // @[Switch.scala 30:36:@1419.4]
  wire  _T_19317; // @[Switch.scala 30:53:@1421.4]
  wire  valid_4_41; // @[Switch.scala 30:36:@1422.4]
  wire  _T_19320; // @[Switch.scala 30:53:@1424.4]
  wire  valid_4_42; // @[Switch.scala 30:36:@1425.4]
  wire  _T_19323; // @[Switch.scala 30:53:@1427.4]
  wire  valid_4_43; // @[Switch.scala 30:36:@1428.4]
  wire  _T_19326; // @[Switch.scala 30:53:@1430.4]
  wire  valid_4_44; // @[Switch.scala 30:36:@1431.4]
  wire  _T_19329; // @[Switch.scala 30:53:@1433.4]
  wire  valid_4_45; // @[Switch.scala 30:36:@1434.4]
  wire  _T_19332; // @[Switch.scala 30:53:@1436.4]
  wire  valid_4_46; // @[Switch.scala 30:36:@1437.4]
  wire  _T_19335; // @[Switch.scala 30:53:@1439.4]
  wire  valid_4_47; // @[Switch.scala 30:36:@1440.4]
  wire  _T_19338; // @[Switch.scala 30:53:@1442.4]
  wire  valid_4_48; // @[Switch.scala 30:36:@1443.4]
  wire  _T_19341; // @[Switch.scala 30:53:@1445.4]
  wire  valid_4_49; // @[Switch.scala 30:36:@1446.4]
  wire  _T_19344; // @[Switch.scala 30:53:@1448.4]
  wire  valid_4_50; // @[Switch.scala 30:36:@1449.4]
  wire  _T_19347; // @[Switch.scala 30:53:@1451.4]
  wire  valid_4_51; // @[Switch.scala 30:36:@1452.4]
  wire  _T_19350; // @[Switch.scala 30:53:@1454.4]
  wire  valid_4_52; // @[Switch.scala 30:36:@1455.4]
  wire  _T_19353; // @[Switch.scala 30:53:@1457.4]
  wire  valid_4_53; // @[Switch.scala 30:36:@1458.4]
  wire  _T_19356; // @[Switch.scala 30:53:@1460.4]
  wire  valid_4_54; // @[Switch.scala 30:36:@1461.4]
  wire  _T_19359; // @[Switch.scala 30:53:@1463.4]
  wire  valid_4_55; // @[Switch.scala 30:36:@1464.4]
  wire  _T_19362; // @[Switch.scala 30:53:@1466.4]
  wire  valid_4_56; // @[Switch.scala 30:36:@1467.4]
  wire  _T_19365; // @[Switch.scala 30:53:@1469.4]
  wire  valid_4_57; // @[Switch.scala 30:36:@1470.4]
  wire  _T_19368; // @[Switch.scala 30:53:@1472.4]
  wire  valid_4_58; // @[Switch.scala 30:36:@1473.4]
  wire  _T_19371; // @[Switch.scala 30:53:@1475.4]
  wire  valid_4_59; // @[Switch.scala 30:36:@1476.4]
  wire  _T_19374; // @[Switch.scala 30:53:@1478.4]
  wire  valid_4_60; // @[Switch.scala 30:36:@1479.4]
  wire  _T_19377; // @[Switch.scala 30:53:@1481.4]
  wire  valid_4_61; // @[Switch.scala 30:36:@1482.4]
  wire  _T_19380; // @[Switch.scala 30:53:@1484.4]
  wire  valid_4_62; // @[Switch.scala 30:36:@1485.4]
  wire  _T_19383; // @[Switch.scala 30:53:@1487.4]
  wire  valid_4_63; // @[Switch.scala 30:36:@1488.4]
  wire [5:0] _T_19449; // @[Mux.scala 31:69:@1490.4]
  wire [5:0] _T_19450; // @[Mux.scala 31:69:@1491.4]
  wire [5:0] _T_19451; // @[Mux.scala 31:69:@1492.4]
  wire [5:0] _T_19452; // @[Mux.scala 31:69:@1493.4]
  wire [5:0] _T_19453; // @[Mux.scala 31:69:@1494.4]
  wire [5:0] _T_19454; // @[Mux.scala 31:69:@1495.4]
  wire [5:0] _T_19455; // @[Mux.scala 31:69:@1496.4]
  wire [5:0] _T_19456; // @[Mux.scala 31:69:@1497.4]
  wire [5:0] _T_19457; // @[Mux.scala 31:69:@1498.4]
  wire [5:0] _T_19458; // @[Mux.scala 31:69:@1499.4]
  wire [5:0] _T_19459; // @[Mux.scala 31:69:@1500.4]
  wire [5:0] _T_19460; // @[Mux.scala 31:69:@1501.4]
  wire [5:0] _T_19461; // @[Mux.scala 31:69:@1502.4]
  wire [5:0] _T_19462; // @[Mux.scala 31:69:@1503.4]
  wire [5:0] _T_19463; // @[Mux.scala 31:69:@1504.4]
  wire [5:0] _T_19464; // @[Mux.scala 31:69:@1505.4]
  wire [5:0] _T_19465; // @[Mux.scala 31:69:@1506.4]
  wire [5:0] _T_19466; // @[Mux.scala 31:69:@1507.4]
  wire [5:0] _T_19467; // @[Mux.scala 31:69:@1508.4]
  wire [5:0] _T_19468; // @[Mux.scala 31:69:@1509.4]
  wire [5:0] _T_19469; // @[Mux.scala 31:69:@1510.4]
  wire [5:0] _T_19470; // @[Mux.scala 31:69:@1511.4]
  wire [5:0] _T_19471; // @[Mux.scala 31:69:@1512.4]
  wire [5:0] _T_19472; // @[Mux.scala 31:69:@1513.4]
  wire [5:0] _T_19473; // @[Mux.scala 31:69:@1514.4]
  wire [5:0] _T_19474; // @[Mux.scala 31:69:@1515.4]
  wire [5:0] _T_19475; // @[Mux.scala 31:69:@1516.4]
  wire [5:0] _T_19476; // @[Mux.scala 31:69:@1517.4]
  wire [5:0] _T_19477; // @[Mux.scala 31:69:@1518.4]
  wire [5:0] _T_19478; // @[Mux.scala 31:69:@1519.4]
  wire [5:0] _T_19479; // @[Mux.scala 31:69:@1520.4]
  wire [5:0] _T_19480; // @[Mux.scala 31:69:@1521.4]
  wire [5:0] _T_19481; // @[Mux.scala 31:69:@1522.4]
  wire [5:0] _T_19482; // @[Mux.scala 31:69:@1523.4]
  wire [5:0] _T_19483; // @[Mux.scala 31:69:@1524.4]
  wire [5:0] _T_19484; // @[Mux.scala 31:69:@1525.4]
  wire [5:0] _T_19485; // @[Mux.scala 31:69:@1526.4]
  wire [5:0] _T_19486; // @[Mux.scala 31:69:@1527.4]
  wire [5:0] _T_19487; // @[Mux.scala 31:69:@1528.4]
  wire [5:0] _T_19488; // @[Mux.scala 31:69:@1529.4]
  wire [5:0] _T_19489; // @[Mux.scala 31:69:@1530.4]
  wire [5:0] _T_19490; // @[Mux.scala 31:69:@1531.4]
  wire [5:0] _T_19491; // @[Mux.scala 31:69:@1532.4]
  wire [5:0] _T_19492; // @[Mux.scala 31:69:@1533.4]
  wire [5:0] _T_19493; // @[Mux.scala 31:69:@1534.4]
  wire [5:0] _T_19494; // @[Mux.scala 31:69:@1535.4]
  wire [5:0] _T_19495; // @[Mux.scala 31:69:@1536.4]
  wire [5:0] _T_19496; // @[Mux.scala 31:69:@1537.4]
  wire [5:0] _T_19497; // @[Mux.scala 31:69:@1538.4]
  wire [5:0] _T_19498; // @[Mux.scala 31:69:@1539.4]
  wire [5:0] _T_19499; // @[Mux.scala 31:69:@1540.4]
  wire [5:0] _T_19500; // @[Mux.scala 31:69:@1541.4]
  wire [5:0] _T_19501; // @[Mux.scala 31:69:@1542.4]
  wire [5:0] _T_19502; // @[Mux.scala 31:69:@1543.4]
  wire [5:0] _T_19503; // @[Mux.scala 31:69:@1544.4]
  wire [5:0] _T_19504; // @[Mux.scala 31:69:@1545.4]
  wire [5:0] _T_19505; // @[Mux.scala 31:69:@1546.4]
  wire [5:0] _T_19506; // @[Mux.scala 31:69:@1547.4]
  wire [5:0] _T_19507; // @[Mux.scala 31:69:@1548.4]
  wire [5:0] _T_19508; // @[Mux.scala 31:69:@1549.4]
  wire [5:0] _T_19509; // @[Mux.scala 31:69:@1550.4]
  wire [5:0] _T_19510; // @[Mux.scala 31:69:@1551.4]
  wire [5:0] select_4; // @[Mux.scala 31:69:@1552.4]
  wire [47:0] _GEN_257; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_258; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_259; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_260; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_261; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_262; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_263; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_264; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_265; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_266; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_267; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_268; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_269; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_270; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_271; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_272; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_273; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_274; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_275; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_276; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_277; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_278; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_279; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_280; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_281; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_282; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_283; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_284; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_285; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_286; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_287; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_288; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_289; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_290; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_291; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_292; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_293; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_294; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_295; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_296; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_297; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_298; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_299; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_300; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_301; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_302; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_303; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_304; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_305; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_306; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_307; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_308; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_309; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_310; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_311; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_312; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_313; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_314; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_315; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_316; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_317; // @[Switch.scala 33:19:@1554.4]
  wire [47:0] _GEN_318; // @[Switch.scala 33:19:@1554.4]
  wire [7:0] _T_19519; // @[Switch.scala 34:32:@1561.4]
  wire [15:0] _T_19527; // @[Switch.scala 34:32:@1569.4]
  wire [7:0] _T_19534; // @[Switch.scala 34:32:@1576.4]
  wire [31:0] _T_19543; // @[Switch.scala 34:32:@1585.4]
  wire [7:0] _T_19550; // @[Switch.scala 34:32:@1592.4]
  wire [15:0] _T_19558; // @[Switch.scala 34:32:@1600.4]
  wire [7:0] _T_19565; // @[Switch.scala 34:32:@1607.4]
  wire [31:0] _T_19574; // @[Switch.scala 34:32:@1616.4]
  wire [63:0] _T_19575; // @[Switch.scala 34:32:@1617.4]
  wire  _T_19579; // @[Switch.scala 30:53:@1620.4]
  wire  valid_5_0; // @[Switch.scala 30:36:@1621.4]
  wire  _T_19582; // @[Switch.scala 30:53:@1623.4]
  wire  valid_5_1; // @[Switch.scala 30:36:@1624.4]
  wire  _T_19585; // @[Switch.scala 30:53:@1626.4]
  wire  valid_5_2; // @[Switch.scala 30:36:@1627.4]
  wire  _T_19588; // @[Switch.scala 30:53:@1629.4]
  wire  valid_5_3; // @[Switch.scala 30:36:@1630.4]
  wire  _T_19591; // @[Switch.scala 30:53:@1632.4]
  wire  valid_5_4; // @[Switch.scala 30:36:@1633.4]
  wire  _T_19594; // @[Switch.scala 30:53:@1635.4]
  wire  valid_5_5; // @[Switch.scala 30:36:@1636.4]
  wire  _T_19597; // @[Switch.scala 30:53:@1638.4]
  wire  valid_5_6; // @[Switch.scala 30:36:@1639.4]
  wire  _T_19600; // @[Switch.scala 30:53:@1641.4]
  wire  valid_5_7; // @[Switch.scala 30:36:@1642.4]
  wire  _T_19603; // @[Switch.scala 30:53:@1644.4]
  wire  valid_5_8; // @[Switch.scala 30:36:@1645.4]
  wire  _T_19606; // @[Switch.scala 30:53:@1647.4]
  wire  valid_5_9; // @[Switch.scala 30:36:@1648.4]
  wire  _T_19609; // @[Switch.scala 30:53:@1650.4]
  wire  valid_5_10; // @[Switch.scala 30:36:@1651.4]
  wire  _T_19612; // @[Switch.scala 30:53:@1653.4]
  wire  valid_5_11; // @[Switch.scala 30:36:@1654.4]
  wire  _T_19615; // @[Switch.scala 30:53:@1656.4]
  wire  valid_5_12; // @[Switch.scala 30:36:@1657.4]
  wire  _T_19618; // @[Switch.scala 30:53:@1659.4]
  wire  valid_5_13; // @[Switch.scala 30:36:@1660.4]
  wire  _T_19621; // @[Switch.scala 30:53:@1662.4]
  wire  valid_5_14; // @[Switch.scala 30:36:@1663.4]
  wire  _T_19624; // @[Switch.scala 30:53:@1665.4]
  wire  valid_5_15; // @[Switch.scala 30:36:@1666.4]
  wire  _T_19627; // @[Switch.scala 30:53:@1668.4]
  wire  valid_5_16; // @[Switch.scala 30:36:@1669.4]
  wire  _T_19630; // @[Switch.scala 30:53:@1671.4]
  wire  valid_5_17; // @[Switch.scala 30:36:@1672.4]
  wire  _T_19633; // @[Switch.scala 30:53:@1674.4]
  wire  valid_5_18; // @[Switch.scala 30:36:@1675.4]
  wire  _T_19636; // @[Switch.scala 30:53:@1677.4]
  wire  valid_5_19; // @[Switch.scala 30:36:@1678.4]
  wire  _T_19639; // @[Switch.scala 30:53:@1680.4]
  wire  valid_5_20; // @[Switch.scala 30:36:@1681.4]
  wire  _T_19642; // @[Switch.scala 30:53:@1683.4]
  wire  valid_5_21; // @[Switch.scala 30:36:@1684.4]
  wire  _T_19645; // @[Switch.scala 30:53:@1686.4]
  wire  valid_5_22; // @[Switch.scala 30:36:@1687.4]
  wire  _T_19648; // @[Switch.scala 30:53:@1689.4]
  wire  valid_5_23; // @[Switch.scala 30:36:@1690.4]
  wire  _T_19651; // @[Switch.scala 30:53:@1692.4]
  wire  valid_5_24; // @[Switch.scala 30:36:@1693.4]
  wire  _T_19654; // @[Switch.scala 30:53:@1695.4]
  wire  valid_5_25; // @[Switch.scala 30:36:@1696.4]
  wire  _T_19657; // @[Switch.scala 30:53:@1698.4]
  wire  valid_5_26; // @[Switch.scala 30:36:@1699.4]
  wire  _T_19660; // @[Switch.scala 30:53:@1701.4]
  wire  valid_5_27; // @[Switch.scala 30:36:@1702.4]
  wire  _T_19663; // @[Switch.scala 30:53:@1704.4]
  wire  valid_5_28; // @[Switch.scala 30:36:@1705.4]
  wire  _T_19666; // @[Switch.scala 30:53:@1707.4]
  wire  valid_5_29; // @[Switch.scala 30:36:@1708.4]
  wire  _T_19669; // @[Switch.scala 30:53:@1710.4]
  wire  valid_5_30; // @[Switch.scala 30:36:@1711.4]
  wire  _T_19672; // @[Switch.scala 30:53:@1713.4]
  wire  valid_5_31; // @[Switch.scala 30:36:@1714.4]
  wire  _T_19675; // @[Switch.scala 30:53:@1716.4]
  wire  valid_5_32; // @[Switch.scala 30:36:@1717.4]
  wire  _T_19678; // @[Switch.scala 30:53:@1719.4]
  wire  valid_5_33; // @[Switch.scala 30:36:@1720.4]
  wire  _T_19681; // @[Switch.scala 30:53:@1722.4]
  wire  valid_5_34; // @[Switch.scala 30:36:@1723.4]
  wire  _T_19684; // @[Switch.scala 30:53:@1725.4]
  wire  valid_5_35; // @[Switch.scala 30:36:@1726.4]
  wire  _T_19687; // @[Switch.scala 30:53:@1728.4]
  wire  valid_5_36; // @[Switch.scala 30:36:@1729.4]
  wire  _T_19690; // @[Switch.scala 30:53:@1731.4]
  wire  valid_5_37; // @[Switch.scala 30:36:@1732.4]
  wire  _T_19693; // @[Switch.scala 30:53:@1734.4]
  wire  valid_5_38; // @[Switch.scala 30:36:@1735.4]
  wire  _T_19696; // @[Switch.scala 30:53:@1737.4]
  wire  valid_5_39; // @[Switch.scala 30:36:@1738.4]
  wire  _T_19699; // @[Switch.scala 30:53:@1740.4]
  wire  valid_5_40; // @[Switch.scala 30:36:@1741.4]
  wire  _T_19702; // @[Switch.scala 30:53:@1743.4]
  wire  valid_5_41; // @[Switch.scala 30:36:@1744.4]
  wire  _T_19705; // @[Switch.scala 30:53:@1746.4]
  wire  valid_5_42; // @[Switch.scala 30:36:@1747.4]
  wire  _T_19708; // @[Switch.scala 30:53:@1749.4]
  wire  valid_5_43; // @[Switch.scala 30:36:@1750.4]
  wire  _T_19711; // @[Switch.scala 30:53:@1752.4]
  wire  valid_5_44; // @[Switch.scala 30:36:@1753.4]
  wire  _T_19714; // @[Switch.scala 30:53:@1755.4]
  wire  valid_5_45; // @[Switch.scala 30:36:@1756.4]
  wire  _T_19717; // @[Switch.scala 30:53:@1758.4]
  wire  valid_5_46; // @[Switch.scala 30:36:@1759.4]
  wire  _T_19720; // @[Switch.scala 30:53:@1761.4]
  wire  valid_5_47; // @[Switch.scala 30:36:@1762.4]
  wire  _T_19723; // @[Switch.scala 30:53:@1764.4]
  wire  valid_5_48; // @[Switch.scala 30:36:@1765.4]
  wire  _T_19726; // @[Switch.scala 30:53:@1767.4]
  wire  valid_5_49; // @[Switch.scala 30:36:@1768.4]
  wire  _T_19729; // @[Switch.scala 30:53:@1770.4]
  wire  valid_5_50; // @[Switch.scala 30:36:@1771.4]
  wire  _T_19732; // @[Switch.scala 30:53:@1773.4]
  wire  valid_5_51; // @[Switch.scala 30:36:@1774.4]
  wire  _T_19735; // @[Switch.scala 30:53:@1776.4]
  wire  valid_5_52; // @[Switch.scala 30:36:@1777.4]
  wire  _T_19738; // @[Switch.scala 30:53:@1779.4]
  wire  valid_5_53; // @[Switch.scala 30:36:@1780.4]
  wire  _T_19741; // @[Switch.scala 30:53:@1782.4]
  wire  valid_5_54; // @[Switch.scala 30:36:@1783.4]
  wire  _T_19744; // @[Switch.scala 30:53:@1785.4]
  wire  valid_5_55; // @[Switch.scala 30:36:@1786.4]
  wire  _T_19747; // @[Switch.scala 30:53:@1788.4]
  wire  valid_5_56; // @[Switch.scala 30:36:@1789.4]
  wire  _T_19750; // @[Switch.scala 30:53:@1791.4]
  wire  valid_5_57; // @[Switch.scala 30:36:@1792.4]
  wire  _T_19753; // @[Switch.scala 30:53:@1794.4]
  wire  valid_5_58; // @[Switch.scala 30:36:@1795.4]
  wire  _T_19756; // @[Switch.scala 30:53:@1797.4]
  wire  valid_5_59; // @[Switch.scala 30:36:@1798.4]
  wire  _T_19759; // @[Switch.scala 30:53:@1800.4]
  wire  valid_5_60; // @[Switch.scala 30:36:@1801.4]
  wire  _T_19762; // @[Switch.scala 30:53:@1803.4]
  wire  valid_5_61; // @[Switch.scala 30:36:@1804.4]
  wire  _T_19765; // @[Switch.scala 30:53:@1806.4]
  wire  valid_5_62; // @[Switch.scala 30:36:@1807.4]
  wire  _T_19768; // @[Switch.scala 30:53:@1809.4]
  wire  valid_5_63; // @[Switch.scala 30:36:@1810.4]
  wire [5:0] _T_19834; // @[Mux.scala 31:69:@1812.4]
  wire [5:0] _T_19835; // @[Mux.scala 31:69:@1813.4]
  wire [5:0] _T_19836; // @[Mux.scala 31:69:@1814.4]
  wire [5:0] _T_19837; // @[Mux.scala 31:69:@1815.4]
  wire [5:0] _T_19838; // @[Mux.scala 31:69:@1816.4]
  wire [5:0] _T_19839; // @[Mux.scala 31:69:@1817.4]
  wire [5:0] _T_19840; // @[Mux.scala 31:69:@1818.4]
  wire [5:0] _T_19841; // @[Mux.scala 31:69:@1819.4]
  wire [5:0] _T_19842; // @[Mux.scala 31:69:@1820.4]
  wire [5:0] _T_19843; // @[Mux.scala 31:69:@1821.4]
  wire [5:0] _T_19844; // @[Mux.scala 31:69:@1822.4]
  wire [5:0] _T_19845; // @[Mux.scala 31:69:@1823.4]
  wire [5:0] _T_19846; // @[Mux.scala 31:69:@1824.4]
  wire [5:0] _T_19847; // @[Mux.scala 31:69:@1825.4]
  wire [5:0] _T_19848; // @[Mux.scala 31:69:@1826.4]
  wire [5:0] _T_19849; // @[Mux.scala 31:69:@1827.4]
  wire [5:0] _T_19850; // @[Mux.scala 31:69:@1828.4]
  wire [5:0] _T_19851; // @[Mux.scala 31:69:@1829.4]
  wire [5:0] _T_19852; // @[Mux.scala 31:69:@1830.4]
  wire [5:0] _T_19853; // @[Mux.scala 31:69:@1831.4]
  wire [5:0] _T_19854; // @[Mux.scala 31:69:@1832.4]
  wire [5:0] _T_19855; // @[Mux.scala 31:69:@1833.4]
  wire [5:0] _T_19856; // @[Mux.scala 31:69:@1834.4]
  wire [5:0] _T_19857; // @[Mux.scala 31:69:@1835.4]
  wire [5:0] _T_19858; // @[Mux.scala 31:69:@1836.4]
  wire [5:0] _T_19859; // @[Mux.scala 31:69:@1837.4]
  wire [5:0] _T_19860; // @[Mux.scala 31:69:@1838.4]
  wire [5:0] _T_19861; // @[Mux.scala 31:69:@1839.4]
  wire [5:0] _T_19862; // @[Mux.scala 31:69:@1840.4]
  wire [5:0] _T_19863; // @[Mux.scala 31:69:@1841.4]
  wire [5:0] _T_19864; // @[Mux.scala 31:69:@1842.4]
  wire [5:0] _T_19865; // @[Mux.scala 31:69:@1843.4]
  wire [5:0] _T_19866; // @[Mux.scala 31:69:@1844.4]
  wire [5:0] _T_19867; // @[Mux.scala 31:69:@1845.4]
  wire [5:0] _T_19868; // @[Mux.scala 31:69:@1846.4]
  wire [5:0] _T_19869; // @[Mux.scala 31:69:@1847.4]
  wire [5:0] _T_19870; // @[Mux.scala 31:69:@1848.4]
  wire [5:0] _T_19871; // @[Mux.scala 31:69:@1849.4]
  wire [5:0] _T_19872; // @[Mux.scala 31:69:@1850.4]
  wire [5:0] _T_19873; // @[Mux.scala 31:69:@1851.4]
  wire [5:0] _T_19874; // @[Mux.scala 31:69:@1852.4]
  wire [5:0] _T_19875; // @[Mux.scala 31:69:@1853.4]
  wire [5:0] _T_19876; // @[Mux.scala 31:69:@1854.4]
  wire [5:0] _T_19877; // @[Mux.scala 31:69:@1855.4]
  wire [5:0] _T_19878; // @[Mux.scala 31:69:@1856.4]
  wire [5:0] _T_19879; // @[Mux.scala 31:69:@1857.4]
  wire [5:0] _T_19880; // @[Mux.scala 31:69:@1858.4]
  wire [5:0] _T_19881; // @[Mux.scala 31:69:@1859.4]
  wire [5:0] _T_19882; // @[Mux.scala 31:69:@1860.4]
  wire [5:0] _T_19883; // @[Mux.scala 31:69:@1861.4]
  wire [5:0] _T_19884; // @[Mux.scala 31:69:@1862.4]
  wire [5:0] _T_19885; // @[Mux.scala 31:69:@1863.4]
  wire [5:0] _T_19886; // @[Mux.scala 31:69:@1864.4]
  wire [5:0] _T_19887; // @[Mux.scala 31:69:@1865.4]
  wire [5:0] _T_19888; // @[Mux.scala 31:69:@1866.4]
  wire [5:0] _T_19889; // @[Mux.scala 31:69:@1867.4]
  wire [5:0] _T_19890; // @[Mux.scala 31:69:@1868.4]
  wire [5:0] _T_19891; // @[Mux.scala 31:69:@1869.4]
  wire [5:0] _T_19892; // @[Mux.scala 31:69:@1870.4]
  wire [5:0] _T_19893; // @[Mux.scala 31:69:@1871.4]
  wire [5:0] _T_19894; // @[Mux.scala 31:69:@1872.4]
  wire [5:0] _T_19895; // @[Mux.scala 31:69:@1873.4]
  wire [5:0] select_5; // @[Mux.scala 31:69:@1874.4]
  wire [47:0] _GEN_321; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_322; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_323; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_324; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_325; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_326; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_327; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_328; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_329; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_330; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_331; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_332; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_333; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_334; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_335; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_336; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_337; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_338; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_339; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_340; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_341; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_342; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_343; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_344; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_345; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_346; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_347; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_348; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_349; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_350; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_351; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_352; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_353; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_354; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_355; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_356; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_357; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_358; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_359; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_360; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_361; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_362; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_363; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_364; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_365; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_366; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_367; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_368; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_369; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_370; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_371; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_372; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_373; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_374; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_375; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_376; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_377; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_378; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_379; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_380; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_381; // @[Switch.scala 33:19:@1876.4]
  wire [47:0] _GEN_382; // @[Switch.scala 33:19:@1876.4]
  wire [7:0] _T_19904; // @[Switch.scala 34:32:@1883.4]
  wire [15:0] _T_19912; // @[Switch.scala 34:32:@1891.4]
  wire [7:0] _T_19919; // @[Switch.scala 34:32:@1898.4]
  wire [31:0] _T_19928; // @[Switch.scala 34:32:@1907.4]
  wire [7:0] _T_19935; // @[Switch.scala 34:32:@1914.4]
  wire [15:0] _T_19943; // @[Switch.scala 34:32:@1922.4]
  wire [7:0] _T_19950; // @[Switch.scala 34:32:@1929.4]
  wire [31:0] _T_19959; // @[Switch.scala 34:32:@1938.4]
  wire [63:0] _T_19960; // @[Switch.scala 34:32:@1939.4]
  wire  _T_19964; // @[Switch.scala 30:53:@1942.4]
  wire  valid_6_0; // @[Switch.scala 30:36:@1943.4]
  wire  _T_19967; // @[Switch.scala 30:53:@1945.4]
  wire  valid_6_1; // @[Switch.scala 30:36:@1946.4]
  wire  _T_19970; // @[Switch.scala 30:53:@1948.4]
  wire  valid_6_2; // @[Switch.scala 30:36:@1949.4]
  wire  _T_19973; // @[Switch.scala 30:53:@1951.4]
  wire  valid_6_3; // @[Switch.scala 30:36:@1952.4]
  wire  _T_19976; // @[Switch.scala 30:53:@1954.4]
  wire  valid_6_4; // @[Switch.scala 30:36:@1955.4]
  wire  _T_19979; // @[Switch.scala 30:53:@1957.4]
  wire  valid_6_5; // @[Switch.scala 30:36:@1958.4]
  wire  _T_19982; // @[Switch.scala 30:53:@1960.4]
  wire  valid_6_6; // @[Switch.scala 30:36:@1961.4]
  wire  _T_19985; // @[Switch.scala 30:53:@1963.4]
  wire  valid_6_7; // @[Switch.scala 30:36:@1964.4]
  wire  _T_19988; // @[Switch.scala 30:53:@1966.4]
  wire  valid_6_8; // @[Switch.scala 30:36:@1967.4]
  wire  _T_19991; // @[Switch.scala 30:53:@1969.4]
  wire  valid_6_9; // @[Switch.scala 30:36:@1970.4]
  wire  _T_19994; // @[Switch.scala 30:53:@1972.4]
  wire  valid_6_10; // @[Switch.scala 30:36:@1973.4]
  wire  _T_19997; // @[Switch.scala 30:53:@1975.4]
  wire  valid_6_11; // @[Switch.scala 30:36:@1976.4]
  wire  _T_20000; // @[Switch.scala 30:53:@1978.4]
  wire  valid_6_12; // @[Switch.scala 30:36:@1979.4]
  wire  _T_20003; // @[Switch.scala 30:53:@1981.4]
  wire  valid_6_13; // @[Switch.scala 30:36:@1982.4]
  wire  _T_20006; // @[Switch.scala 30:53:@1984.4]
  wire  valid_6_14; // @[Switch.scala 30:36:@1985.4]
  wire  _T_20009; // @[Switch.scala 30:53:@1987.4]
  wire  valid_6_15; // @[Switch.scala 30:36:@1988.4]
  wire  _T_20012; // @[Switch.scala 30:53:@1990.4]
  wire  valid_6_16; // @[Switch.scala 30:36:@1991.4]
  wire  _T_20015; // @[Switch.scala 30:53:@1993.4]
  wire  valid_6_17; // @[Switch.scala 30:36:@1994.4]
  wire  _T_20018; // @[Switch.scala 30:53:@1996.4]
  wire  valid_6_18; // @[Switch.scala 30:36:@1997.4]
  wire  _T_20021; // @[Switch.scala 30:53:@1999.4]
  wire  valid_6_19; // @[Switch.scala 30:36:@2000.4]
  wire  _T_20024; // @[Switch.scala 30:53:@2002.4]
  wire  valid_6_20; // @[Switch.scala 30:36:@2003.4]
  wire  _T_20027; // @[Switch.scala 30:53:@2005.4]
  wire  valid_6_21; // @[Switch.scala 30:36:@2006.4]
  wire  _T_20030; // @[Switch.scala 30:53:@2008.4]
  wire  valid_6_22; // @[Switch.scala 30:36:@2009.4]
  wire  _T_20033; // @[Switch.scala 30:53:@2011.4]
  wire  valid_6_23; // @[Switch.scala 30:36:@2012.4]
  wire  _T_20036; // @[Switch.scala 30:53:@2014.4]
  wire  valid_6_24; // @[Switch.scala 30:36:@2015.4]
  wire  _T_20039; // @[Switch.scala 30:53:@2017.4]
  wire  valid_6_25; // @[Switch.scala 30:36:@2018.4]
  wire  _T_20042; // @[Switch.scala 30:53:@2020.4]
  wire  valid_6_26; // @[Switch.scala 30:36:@2021.4]
  wire  _T_20045; // @[Switch.scala 30:53:@2023.4]
  wire  valid_6_27; // @[Switch.scala 30:36:@2024.4]
  wire  _T_20048; // @[Switch.scala 30:53:@2026.4]
  wire  valid_6_28; // @[Switch.scala 30:36:@2027.4]
  wire  _T_20051; // @[Switch.scala 30:53:@2029.4]
  wire  valid_6_29; // @[Switch.scala 30:36:@2030.4]
  wire  _T_20054; // @[Switch.scala 30:53:@2032.4]
  wire  valid_6_30; // @[Switch.scala 30:36:@2033.4]
  wire  _T_20057; // @[Switch.scala 30:53:@2035.4]
  wire  valid_6_31; // @[Switch.scala 30:36:@2036.4]
  wire  _T_20060; // @[Switch.scala 30:53:@2038.4]
  wire  valid_6_32; // @[Switch.scala 30:36:@2039.4]
  wire  _T_20063; // @[Switch.scala 30:53:@2041.4]
  wire  valid_6_33; // @[Switch.scala 30:36:@2042.4]
  wire  _T_20066; // @[Switch.scala 30:53:@2044.4]
  wire  valid_6_34; // @[Switch.scala 30:36:@2045.4]
  wire  _T_20069; // @[Switch.scala 30:53:@2047.4]
  wire  valid_6_35; // @[Switch.scala 30:36:@2048.4]
  wire  _T_20072; // @[Switch.scala 30:53:@2050.4]
  wire  valid_6_36; // @[Switch.scala 30:36:@2051.4]
  wire  _T_20075; // @[Switch.scala 30:53:@2053.4]
  wire  valid_6_37; // @[Switch.scala 30:36:@2054.4]
  wire  _T_20078; // @[Switch.scala 30:53:@2056.4]
  wire  valid_6_38; // @[Switch.scala 30:36:@2057.4]
  wire  _T_20081; // @[Switch.scala 30:53:@2059.4]
  wire  valid_6_39; // @[Switch.scala 30:36:@2060.4]
  wire  _T_20084; // @[Switch.scala 30:53:@2062.4]
  wire  valid_6_40; // @[Switch.scala 30:36:@2063.4]
  wire  _T_20087; // @[Switch.scala 30:53:@2065.4]
  wire  valid_6_41; // @[Switch.scala 30:36:@2066.4]
  wire  _T_20090; // @[Switch.scala 30:53:@2068.4]
  wire  valid_6_42; // @[Switch.scala 30:36:@2069.4]
  wire  _T_20093; // @[Switch.scala 30:53:@2071.4]
  wire  valid_6_43; // @[Switch.scala 30:36:@2072.4]
  wire  _T_20096; // @[Switch.scala 30:53:@2074.4]
  wire  valid_6_44; // @[Switch.scala 30:36:@2075.4]
  wire  _T_20099; // @[Switch.scala 30:53:@2077.4]
  wire  valid_6_45; // @[Switch.scala 30:36:@2078.4]
  wire  _T_20102; // @[Switch.scala 30:53:@2080.4]
  wire  valid_6_46; // @[Switch.scala 30:36:@2081.4]
  wire  _T_20105; // @[Switch.scala 30:53:@2083.4]
  wire  valid_6_47; // @[Switch.scala 30:36:@2084.4]
  wire  _T_20108; // @[Switch.scala 30:53:@2086.4]
  wire  valid_6_48; // @[Switch.scala 30:36:@2087.4]
  wire  _T_20111; // @[Switch.scala 30:53:@2089.4]
  wire  valid_6_49; // @[Switch.scala 30:36:@2090.4]
  wire  _T_20114; // @[Switch.scala 30:53:@2092.4]
  wire  valid_6_50; // @[Switch.scala 30:36:@2093.4]
  wire  _T_20117; // @[Switch.scala 30:53:@2095.4]
  wire  valid_6_51; // @[Switch.scala 30:36:@2096.4]
  wire  _T_20120; // @[Switch.scala 30:53:@2098.4]
  wire  valid_6_52; // @[Switch.scala 30:36:@2099.4]
  wire  _T_20123; // @[Switch.scala 30:53:@2101.4]
  wire  valid_6_53; // @[Switch.scala 30:36:@2102.4]
  wire  _T_20126; // @[Switch.scala 30:53:@2104.4]
  wire  valid_6_54; // @[Switch.scala 30:36:@2105.4]
  wire  _T_20129; // @[Switch.scala 30:53:@2107.4]
  wire  valid_6_55; // @[Switch.scala 30:36:@2108.4]
  wire  _T_20132; // @[Switch.scala 30:53:@2110.4]
  wire  valid_6_56; // @[Switch.scala 30:36:@2111.4]
  wire  _T_20135; // @[Switch.scala 30:53:@2113.4]
  wire  valid_6_57; // @[Switch.scala 30:36:@2114.4]
  wire  _T_20138; // @[Switch.scala 30:53:@2116.4]
  wire  valid_6_58; // @[Switch.scala 30:36:@2117.4]
  wire  _T_20141; // @[Switch.scala 30:53:@2119.4]
  wire  valid_6_59; // @[Switch.scala 30:36:@2120.4]
  wire  _T_20144; // @[Switch.scala 30:53:@2122.4]
  wire  valid_6_60; // @[Switch.scala 30:36:@2123.4]
  wire  _T_20147; // @[Switch.scala 30:53:@2125.4]
  wire  valid_6_61; // @[Switch.scala 30:36:@2126.4]
  wire  _T_20150; // @[Switch.scala 30:53:@2128.4]
  wire  valid_6_62; // @[Switch.scala 30:36:@2129.4]
  wire  _T_20153; // @[Switch.scala 30:53:@2131.4]
  wire  valid_6_63; // @[Switch.scala 30:36:@2132.4]
  wire [5:0] _T_20219; // @[Mux.scala 31:69:@2134.4]
  wire [5:0] _T_20220; // @[Mux.scala 31:69:@2135.4]
  wire [5:0] _T_20221; // @[Mux.scala 31:69:@2136.4]
  wire [5:0] _T_20222; // @[Mux.scala 31:69:@2137.4]
  wire [5:0] _T_20223; // @[Mux.scala 31:69:@2138.4]
  wire [5:0] _T_20224; // @[Mux.scala 31:69:@2139.4]
  wire [5:0] _T_20225; // @[Mux.scala 31:69:@2140.4]
  wire [5:0] _T_20226; // @[Mux.scala 31:69:@2141.4]
  wire [5:0] _T_20227; // @[Mux.scala 31:69:@2142.4]
  wire [5:0] _T_20228; // @[Mux.scala 31:69:@2143.4]
  wire [5:0] _T_20229; // @[Mux.scala 31:69:@2144.4]
  wire [5:0] _T_20230; // @[Mux.scala 31:69:@2145.4]
  wire [5:0] _T_20231; // @[Mux.scala 31:69:@2146.4]
  wire [5:0] _T_20232; // @[Mux.scala 31:69:@2147.4]
  wire [5:0] _T_20233; // @[Mux.scala 31:69:@2148.4]
  wire [5:0] _T_20234; // @[Mux.scala 31:69:@2149.4]
  wire [5:0] _T_20235; // @[Mux.scala 31:69:@2150.4]
  wire [5:0] _T_20236; // @[Mux.scala 31:69:@2151.4]
  wire [5:0] _T_20237; // @[Mux.scala 31:69:@2152.4]
  wire [5:0] _T_20238; // @[Mux.scala 31:69:@2153.4]
  wire [5:0] _T_20239; // @[Mux.scala 31:69:@2154.4]
  wire [5:0] _T_20240; // @[Mux.scala 31:69:@2155.4]
  wire [5:0] _T_20241; // @[Mux.scala 31:69:@2156.4]
  wire [5:0] _T_20242; // @[Mux.scala 31:69:@2157.4]
  wire [5:0] _T_20243; // @[Mux.scala 31:69:@2158.4]
  wire [5:0] _T_20244; // @[Mux.scala 31:69:@2159.4]
  wire [5:0] _T_20245; // @[Mux.scala 31:69:@2160.4]
  wire [5:0] _T_20246; // @[Mux.scala 31:69:@2161.4]
  wire [5:0] _T_20247; // @[Mux.scala 31:69:@2162.4]
  wire [5:0] _T_20248; // @[Mux.scala 31:69:@2163.4]
  wire [5:0] _T_20249; // @[Mux.scala 31:69:@2164.4]
  wire [5:0] _T_20250; // @[Mux.scala 31:69:@2165.4]
  wire [5:0] _T_20251; // @[Mux.scala 31:69:@2166.4]
  wire [5:0] _T_20252; // @[Mux.scala 31:69:@2167.4]
  wire [5:0] _T_20253; // @[Mux.scala 31:69:@2168.4]
  wire [5:0] _T_20254; // @[Mux.scala 31:69:@2169.4]
  wire [5:0] _T_20255; // @[Mux.scala 31:69:@2170.4]
  wire [5:0] _T_20256; // @[Mux.scala 31:69:@2171.4]
  wire [5:0] _T_20257; // @[Mux.scala 31:69:@2172.4]
  wire [5:0] _T_20258; // @[Mux.scala 31:69:@2173.4]
  wire [5:0] _T_20259; // @[Mux.scala 31:69:@2174.4]
  wire [5:0] _T_20260; // @[Mux.scala 31:69:@2175.4]
  wire [5:0] _T_20261; // @[Mux.scala 31:69:@2176.4]
  wire [5:0] _T_20262; // @[Mux.scala 31:69:@2177.4]
  wire [5:0] _T_20263; // @[Mux.scala 31:69:@2178.4]
  wire [5:0] _T_20264; // @[Mux.scala 31:69:@2179.4]
  wire [5:0] _T_20265; // @[Mux.scala 31:69:@2180.4]
  wire [5:0] _T_20266; // @[Mux.scala 31:69:@2181.4]
  wire [5:0] _T_20267; // @[Mux.scala 31:69:@2182.4]
  wire [5:0] _T_20268; // @[Mux.scala 31:69:@2183.4]
  wire [5:0] _T_20269; // @[Mux.scala 31:69:@2184.4]
  wire [5:0] _T_20270; // @[Mux.scala 31:69:@2185.4]
  wire [5:0] _T_20271; // @[Mux.scala 31:69:@2186.4]
  wire [5:0] _T_20272; // @[Mux.scala 31:69:@2187.4]
  wire [5:0] _T_20273; // @[Mux.scala 31:69:@2188.4]
  wire [5:0] _T_20274; // @[Mux.scala 31:69:@2189.4]
  wire [5:0] _T_20275; // @[Mux.scala 31:69:@2190.4]
  wire [5:0] _T_20276; // @[Mux.scala 31:69:@2191.4]
  wire [5:0] _T_20277; // @[Mux.scala 31:69:@2192.4]
  wire [5:0] _T_20278; // @[Mux.scala 31:69:@2193.4]
  wire [5:0] _T_20279; // @[Mux.scala 31:69:@2194.4]
  wire [5:0] _T_20280; // @[Mux.scala 31:69:@2195.4]
  wire [5:0] select_6; // @[Mux.scala 31:69:@2196.4]
  wire [47:0] _GEN_385; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_386; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_387; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_388; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_389; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_390; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_391; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_392; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_393; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_394; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_395; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_396; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_397; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_398; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_399; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_400; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_401; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_402; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_403; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_404; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_405; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_406; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_407; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_408; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_409; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_410; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_411; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_412; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_413; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_414; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_415; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_416; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_417; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_418; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_419; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_420; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_421; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_422; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_423; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_424; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_425; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_426; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_427; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_428; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_429; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_430; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_431; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_432; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_433; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_434; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_435; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_436; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_437; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_438; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_439; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_440; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_441; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_442; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_443; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_444; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_445; // @[Switch.scala 33:19:@2198.4]
  wire [47:0] _GEN_446; // @[Switch.scala 33:19:@2198.4]
  wire [7:0] _T_20289; // @[Switch.scala 34:32:@2205.4]
  wire [15:0] _T_20297; // @[Switch.scala 34:32:@2213.4]
  wire [7:0] _T_20304; // @[Switch.scala 34:32:@2220.4]
  wire [31:0] _T_20313; // @[Switch.scala 34:32:@2229.4]
  wire [7:0] _T_20320; // @[Switch.scala 34:32:@2236.4]
  wire [15:0] _T_20328; // @[Switch.scala 34:32:@2244.4]
  wire [7:0] _T_20335; // @[Switch.scala 34:32:@2251.4]
  wire [31:0] _T_20344; // @[Switch.scala 34:32:@2260.4]
  wire [63:0] _T_20345; // @[Switch.scala 34:32:@2261.4]
  wire  _T_20349; // @[Switch.scala 30:53:@2264.4]
  wire  valid_7_0; // @[Switch.scala 30:36:@2265.4]
  wire  _T_20352; // @[Switch.scala 30:53:@2267.4]
  wire  valid_7_1; // @[Switch.scala 30:36:@2268.4]
  wire  _T_20355; // @[Switch.scala 30:53:@2270.4]
  wire  valid_7_2; // @[Switch.scala 30:36:@2271.4]
  wire  _T_20358; // @[Switch.scala 30:53:@2273.4]
  wire  valid_7_3; // @[Switch.scala 30:36:@2274.4]
  wire  _T_20361; // @[Switch.scala 30:53:@2276.4]
  wire  valid_7_4; // @[Switch.scala 30:36:@2277.4]
  wire  _T_20364; // @[Switch.scala 30:53:@2279.4]
  wire  valid_7_5; // @[Switch.scala 30:36:@2280.4]
  wire  _T_20367; // @[Switch.scala 30:53:@2282.4]
  wire  valid_7_6; // @[Switch.scala 30:36:@2283.4]
  wire  _T_20370; // @[Switch.scala 30:53:@2285.4]
  wire  valid_7_7; // @[Switch.scala 30:36:@2286.4]
  wire  _T_20373; // @[Switch.scala 30:53:@2288.4]
  wire  valid_7_8; // @[Switch.scala 30:36:@2289.4]
  wire  _T_20376; // @[Switch.scala 30:53:@2291.4]
  wire  valid_7_9; // @[Switch.scala 30:36:@2292.4]
  wire  _T_20379; // @[Switch.scala 30:53:@2294.4]
  wire  valid_7_10; // @[Switch.scala 30:36:@2295.4]
  wire  _T_20382; // @[Switch.scala 30:53:@2297.4]
  wire  valid_7_11; // @[Switch.scala 30:36:@2298.4]
  wire  _T_20385; // @[Switch.scala 30:53:@2300.4]
  wire  valid_7_12; // @[Switch.scala 30:36:@2301.4]
  wire  _T_20388; // @[Switch.scala 30:53:@2303.4]
  wire  valid_7_13; // @[Switch.scala 30:36:@2304.4]
  wire  _T_20391; // @[Switch.scala 30:53:@2306.4]
  wire  valid_7_14; // @[Switch.scala 30:36:@2307.4]
  wire  _T_20394; // @[Switch.scala 30:53:@2309.4]
  wire  valid_7_15; // @[Switch.scala 30:36:@2310.4]
  wire  _T_20397; // @[Switch.scala 30:53:@2312.4]
  wire  valid_7_16; // @[Switch.scala 30:36:@2313.4]
  wire  _T_20400; // @[Switch.scala 30:53:@2315.4]
  wire  valid_7_17; // @[Switch.scala 30:36:@2316.4]
  wire  _T_20403; // @[Switch.scala 30:53:@2318.4]
  wire  valid_7_18; // @[Switch.scala 30:36:@2319.4]
  wire  _T_20406; // @[Switch.scala 30:53:@2321.4]
  wire  valid_7_19; // @[Switch.scala 30:36:@2322.4]
  wire  _T_20409; // @[Switch.scala 30:53:@2324.4]
  wire  valid_7_20; // @[Switch.scala 30:36:@2325.4]
  wire  _T_20412; // @[Switch.scala 30:53:@2327.4]
  wire  valid_7_21; // @[Switch.scala 30:36:@2328.4]
  wire  _T_20415; // @[Switch.scala 30:53:@2330.4]
  wire  valid_7_22; // @[Switch.scala 30:36:@2331.4]
  wire  _T_20418; // @[Switch.scala 30:53:@2333.4]
  wire  valid_7_23; // @[Switch.scala 30:36:@2334.4]
  wire  _T_20421; // @[Switch.scala 30:53:@2336.4]
  wire  valid_7_24; // @[Switch.scala 30:36:@2337.4]
  wire  _T_20424; // @[Switch.scala 30:53:@2339.4]
  wire  valid_7_25; // @[Switch.scala 30:36:@2340.4]
  wire  _T_20427; // @[Switch.scala 30:53:@2342.4]
  wire  valid_7_26; // @[Switch.scala 30:36:@2343.4]
  wire  _T_20430; // @[Switch.scala 30:53:@2345.4]
  wire  valid_7_27; // @[Switch.scala 30:36:@2346.4]
  wire  _T_20433; // @[Switch.scala 30:53:@2348.4]
  wire  valid_7_28; // @[Switch.scala 30:36:@2349.4]
  wire  _T_20436; // @[Switch.scala 30:53:@2351.4]
  wire  valid_7_29; // @[Switch.scala 30:36:@2352.4]
  wire  _T_20439; // @[Switch.scala 30:53:@2354.4]
  wire  valid_7_30; // @[Switch.scala 30:36:@2355.4]
  wire  _T_20442; // @[Switch.scala 30:53:@2357.4]
  wire  valid_7_31; // @[Switch.scala 30:36:@2358.4]
  wire  _T_20445; // @[Switch.scala 30:53:@2360.4]
  wire  valid_7_32; // @[Switch.scala 30:36:@2361.4]
  wire  _T_20448; // @[Switch.scala 30:53:@2363.4]
  wire  valid_7_33; // @[Switch.scala 30:36:@2364.4]
  wire  _T_20451; // @[Switch.scala 30:53:@2366.4]
  wire  valid_7_34; // @[Switch.scala 30:36:@2367.4]
  wire  _T_20454; // @[Switch.scala 30:53:@2369.4]
  wire  valid_7_35; // @[Switch.scala 30:36:@2370.4]
  wire  _T_20457; // @[Switch.scala 30:53:@2372.4]
  wire  valid_7_36; // @[Switch.scala 30:36:@2373.4]
  wire  _T_20460; // @[Switch.scala 30:53:@2375.4]
  wire  valid_7_37; // @[Switch.scala 30:36:@2376.4]
  wire  _T_20463; // @[Switch.scala 30:53:@2378.4]
  wire  valid_7_38; // @[Switch.scala 30:36:@2379.4]
  wire  _T_20466; // @[Switch.scala 30:53:@2381.4]
  wire  valid_7_39; // @[Switch.scala 30:36:@2382.4]
  wire  _T_20469; // @[Switch.scala 30:53:@2384.4]
  wire  valid_7_40; // @[Switch.scala 30:36:@2385.4]
  wire  _T_20472; // @[Switch.scala 30:53:@2387.4]
  wire  valid_7_41; // @[Switch.scala 30:36:@2388.4]
  wire  _T_20475; // @[Switch.scala 30:53:@2390.4]
  wire  valid_7_42; // @[Switch.scala 30:36:@2391.4]
  wire  _T_20478; // @[Switch.scala 30:53:@2393.4]
  wire  valid_7_43; // @[Switch.scala 30:36:@2394.4]
  wire  _T_20481; // @[Switch.scala 30:53:@2396.4]
  wire  valid_7_44; // @[Switch.scala 30:36:@2397.4]
  wire  _T_20484; // @[Switch.scala 30:53:@2399.4]
  wire  valid_7_45; // @[Switch.scala 30:36:@2400.4]
  wire  _T_20487; // @[Switch.scala 30:53:@2402.4]
  wire  valid_7_46; // @[Switch.scala 30:36:@2403.4]
  wire  _T_20490; // @[Switch.scala 30:53:@2405.4]
  wire  valid_7_47; // @[Switch.scala 30:36:@2406.4]
  wire  _T_20493; // @[Switch.scala 30:53:@2408.4]
  wire  valid_7_48; // @[Switch.scala 30:36:@2409.4]
  wire  _T_20496; // @[Switch.scala 30:53:@2411.4]
  wire  valid_7_49; // @[Switch.scala 30:36:@2412.4]
  wire  _T_20499; // @[Switch.scala 30:53:@2414.4]
  wire  valid_7_50; // @[Switch.scala 30:36:@2415.4]
  wire  _T_20502; // @[Switch.scala 30:53:@2417.4]
  wire  valid_7_51; // @[Switch.scala 30:36:@2418.4]
  wire  _T_20505; // @[Switch.scala 30:53:@2420.4]
  wire  valid_7_52; // @[Switch.scala 30:36:@2421.4]
  wire  _T_20508; // @[Switch.scala 30:53:@2423.4]
  wire  valid_7_53; // @[Switch.scala 30:36:@2424.4]
  wire  _T_20511; // @[Switch.scala 30:53:@2426.4]
  wire  valid_7_54; // @[Switch.scala 30:36:@2427.4]
  wire  _T_20514; // @[Switch.scala 30:53:@2429.4]
  wire  valid_7_55; // @[Switch.scala 30:36:@2430.4]
  wire  _T_20517; // @[Switch.scala 30:53:@2432.4]
  wire  valid_7_56; // @[Switch.scala 30:36:@2433.4]
  wire  _T_20520; // @[Switch.scala 30:53:@2435.4]
  wire  valid_7_57; // @[Switch.scala 30:36:@2436.4]
  wire  _T_20523; // @[Switch.scala 30:53:@2438.4]
  wire  valid_7_58; // @[Switch.scala 30:36:@2439.4]
  wire  _T_20526; // @[Switch.scala 30:53:@2441.4]
  wire  valid_7_59; // @[Switch.scala 30:36:@2442.4]
  wire  _T_20529; // @[Switch.scala 30:53:@2444.4]
  wire  valid_7_60; // @[Switch.scala 30:36:@2445.4]
  wire  _T_20532; // @[Switch.scala 30:53:@2447.4]
  wire  valid_7_61; // @[Switch.scala 30:36:@2448.4]
  wire  _T_20535; // @[Switch.scala 30:53:@2450.4]
  wire  valid_7_62; // @[Switch.scala 30:36:@2451.4]
  wire  _T_20538; // @[Switch.scala 30:53:@2453.4]
  wire  valid_7_63; // @[Switch.scala 30:36:@2454.4]
  wire [5:0] _T_20604; // @[Mux.scala 31:69:@2456.4]
  wire [5:0] _T_20605; // @[Mux.scala 31:69:@2457.4]
  wire [5:0] _T_20606; // @[Mux.scala 31:69:@2458.4]
  wire [5:0] _T_20607; // @[Mux.scala 31:69:@2459.4]
  wire [5:0] _T_20608; // @[Mux.scala 31:69:@2460.4]
  wire [5:0] _T_20609; // @[Mux.scala 31:69:@2461.4]
  wire [5:0] _T_20610; // @[Mux.scala 31:69:@2462.4]
  wire [5:0] _T_20611; // @[Mux.scala 31:69:@2463.4]
  wire [5:0] _T_20612; // @[Mux.scala 31:69:@2464.4]
  wire [5:0] _T_20613; // @[Mux.scala 31:69:@2465.4]
  wire [5:0] _T_20614; // @[Mux.scala 31:69:@2466.4]
  wire [5:0] _T_20615; // @[Mux.scala 31:69:@2467.4]
  wire [5:0] _T_20616; // @[Mux.scala 31:69:@2468.4]
  wire [5:0] _T_20617; // @[Mux.scala 31:69:@2469.4]
  wire [5:0] _T_20618; // @[Mux.scala 31:69:@2470.4]
  wire [5:0] _T_20619; // @[Mux.scala 31:69:@2471.4]
  wire [5:0] _T_20620; // @[Mux.scala 31:69:@2472.4]
  wire [5:0] _T_20621; // @[Mux.scala 31:69:@2473.4]
  wire [5:0] _T_20622; // @[Mux.scala 31:69:@2474.4]
  wire [5:0] _T_20623; // @[Mux.scala 31:69:@2475.4]
  wire [5:0] _T_20624; // @[Mux.scala 31:69:@2476.4]
  wire [5:0] _T_20625; // @[Mux.scala 31:69:@2477.4]
  wire [5:0] _T_20626; // @[Mux.scala 31:69:@2478.4]
  wire [5:0] _T_20627; // @[Mux.scala 31:69:@2479.4]
  wire [5:0] _T_20628; // @[Mux.scala 31:69:@2480.4]
  wire [5:0] _T_20629; // @[Mux.scala 31:69:@2481.4]
  wire [5:0] _T_20630; // @[Mux.scala 31:69:@2482.4]
  wire [5:0] _T_20631; // @[Mux.scala 31:69:@2483.4]
  wire [5:0] _T_20632; // @[Mux.scala 31:69:@2484.4]
  wire [5:0] _T_20633; // @[Mux.scala 31:69:@2485.4]
  wire [5:0] _T_20634; // @[Mux.scala 31:69:@2486.4]
  wire [5:0] _T_20635; // @[Mux.scala 31:69:@2487.4]
  wire [5:0] _T_20636; // @[Mux.scala 31:69:@2488.4]
  wire [5:0] _T_20637; // @[Mux.scala 31:69:@2489.4]
  wire [5:0] _T_20638; // @[Mux.scala 31:69:@2490.4]
  wire [5:0] _T_20639; // @[Mux.scala 31:69:@2491.4]
  wire [5:0] _T_20640; // @[Mux.scala 31:69:@2492.4]
  wire [5:0] _T_20641; // @[Mux.scala 31:69:@2493.4]
  wire [5:0] _T_20642; // @[Mux.scala 31:69:@2494.4]
  wire [5:0] _T_20643; // @[Mux.scala 31:69:@2495.4]
  wire [5:0] _T_20644; // @[Mux.scala 31:69:@2496.4]
  wire [5:0] _T_20645; // @[Mux.scala 31:69:@2497.4]
  wire [5:0] _T_20646; // @[Mux.scala 31:69:@2498.4]
  wire [5:0] _T_20647; // @[Mux.scala 31:69:@2499.4]
  wire [5:0] _T_20648; // @[Mux.scala 31:69:@2500.4]
  wire [5:0] _T_20649; // @[Mux.scala 31:69:@2501.4]
  wire [5:0] _T_20650; // @[Mux.scala 31:69:@2502.4]
  wire [5:0] _T_20651; // @[Mux.scala 31:69:@2503.4]
  wire [5:0] _T_20652; // @[Mux.scala 31:69:@2504.4]
  wire [5:0] _T_20653; // @[Mux.scala 31:69:@2505.4]
  wire [5:0] _T_20654; // @[Mux.scala 31:69:@2506.4]
  wire [5:0] _T_20655; // @[Mux.scala 31:69:@2507.4]
  wire [5:0] _T_20656; // @[Mux.scala 31:69:@2508.4]
  wire [5:0] _T_20657; // @[Mux.scala 31:69:@2509.4]
  wire [5:0] _T_20658; // @[Mux.scala 31:69:@2510.4]
  wire [5:0] _T_20659; // @[Mux.scala 31:69:@2511.4]
  wire [5:0] _T_20660; // @[Mux.scala 31:69:@2512.4]
  wire [5:0] _T_20661; // @[Mux.scala 31:69:@2513.4]
  wire [5:0] _T_20662; // @[Mux.scala 31:69:@2514.4]
  wire [5:0] _T_20663; // @[Mux.scala 31:69:@2515.4]
  wire [5:0] _T_20664; // @[Mux.scala 31:69:@2516.4]
  wire [5:0] _T_20665; // @[Mux.scala 31:69:@2517.4]
  wire [5:0] select_7; // @[Mux.scala 31:69:@2518.4]
  wire [47:0] _GEN_449; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_450; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_451; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_452; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_453; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_454; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_455; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_456; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_457; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_458; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_459; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_460; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_461; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_462; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_463; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_464; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_465; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_466; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_467; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_468; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_469; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_470; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_471; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_472; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_473; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_474; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_475; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_476; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_477; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_478; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_479; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_480; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_481; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_482; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_483; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_484; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_485; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_486; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_487; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_488; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_489; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_490; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_491; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_492; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_493; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_494; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_495; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_496; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_497; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_498; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_499; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_500; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_501; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_502; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_503; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_504; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_505; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_506; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_507; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_508; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_509; // @[Switch.scala 33:19:@2520.4]
  wire [47:0] _GEN_510; // @[Switch.scala 33:19:@2520.4]
  wire [7:0] _T_20674; // @[Switch.scala 34:32:@2527.4]
  wire [15:0] _T_20682; // @[Switch.scala 34:32:@2535.4]
  wire [7:0] _T_20689; // @[Switch.scala 34:32:@2542.4]
  wire [31:0] _T_20698; // @[Switch.scala 34:32:@2551.4]
  wire [7:0] _T_20705; // @[Switch.scala 34:32:@2558.4]
  wire [15:0] _T_20713; // @[Switch.scala 34:32:@2566.4]
  wire [7:0] _T_20720; // @[Switch.scala 34:32:@2573.4]
  wire [31:0] _T_20729; // @[Switch.scala 34:32:@2582.4]
  wire [63:0] _T_20730; // @[Switch.scala 34:32:@2583.4]
  wire  _T_20734; // @[Switch.scala 30:53:@2586.4]
  wire  valid_8_0; // @[Switch.scala 30:36:@2587.4]
  wire  _T_20737; // @[Switch.scala 30:53:@2589.4]
  wire  valid_8_1; // @[Switch.scala 30:36:@2590.4]
  wire  _T_20740; // @[Switch.scala 30:53:@2592.4]
  wire  valid_8_2; // @[Switch.scala 30:36:@2593.4]
  wire  _T_20743; // @[Switch.scala 30:53:@2595.4]
  wire  valid_8_3; // @[Switch.scala 30:36:@2596.4]
  wire  _T_20746; // @[Switch.scala 30:53:@2598.4]
  wire  valid_8_4; // @[Switch.scala 30:36:@2599.4]
  wire  _T_20749; // @[Switch.scala 30:53:@2601.4]
  wire  valid_8_5; // @[Switch.scala 30:36:@2602.4]
  wire  _T_20752; // @[Switch.scala 30:53:@2604.4]
  wire  valid_8_6; // @[Switch.scala 30:36:@2605.4]
  wire  _T_20755; // @[Switch.scala 30:53:@2607.4]
  wire  valid_8_7; // @[Switch.scala 30:36:@2608.4]
  wire  _T_20758; // @[Switch.scala 30:53:@2610.4]
  wire  valid_8_8; // @[Switch.scala 30:36:@2611.4]
  wire  _T_20761; // @[Switch.scala 30:53:@2613.4]
  wire  valid_8_9; // @[Switch.scala 30:36:@2614.4]
  wire  _T_20764; // @[Switch.scala 30:53:@2616.4]
  wire  valid_8_10; // @[Switch.scala 30:36:@2617.4]
  wire  _T_20767; // @[Switch.scala 30:53:@2619.4]
  wire  valid_8_11; // @[Switch.scala 30:36:@2620.4]
  wire  _T_20770; // @[Switch.scala 30:53:@2622.4]
  wire  valid_8_12; // @[Switch.scala 30:36:@2623.4]
  wire  _T_20773; // @[Switch.scala 30:53:@2625.4]
  wire  valid_8_13; // @[Switch.scala 30:36:@2626.4]
  wire  _T_20776; // @[Switch.scala 30:53:@2628.4]
  wire  valid_8_14; // @[Switch.scala 30:36:@2629.4]
  wire  _T_20779; // @[Switch.scala 30:53:@2631.4]
  wire  valid_8_15; // @[Switch.scala 30:36:@2632.4]
  wire  _T_20782; // @[Switch.scala 30:53:@2634.4]
  wire  valid_8_16; // @[Switch.scala 30:36:@2635.4]
  wire  _T_20785; // @[Switch.scala 30:53:@2637.4]
  wire  valid_8_17; // @[Switch.scala 30:36:@2638.4]
  wire  _T_20788; // @[Switch.scala 30:53:@2640.4]
  wire  valid_8_18; // @[Switch.scala 30:36:@2641.4]
  wire  _T_20791; // @[Switch.scala 30:53:@2643.4]
  wire  valid_8_19; // @[Switch.scala 30:36:@2644.4]
  wire  _T_20794; // @[Switch.scala 30:53:@2646.4]
  wire  valid_8_20; // @[Switch.scala 30:36:@2647.4]
  wire  _T_20797; // @[Switch.scala 30:53:@2649.4]
  wire  valid_8_21; // @[Switch.scala 30:36:@2650.4]
  wire  _T_20800; // @[Switch.scala 30:53:@2652.4]
  wire  valid_8_22; // @[Switch.scala 30:36:@2653.4]
  wire  _T_20803; // @[Switch.scala 30:53:@2655.4]
  wire  valid_8_23; // @[Switch.scala 30:36:@2656.4]
  wire  _T_20806; // @[Switch.scala 30:53:@2658.4]
  wire  valid_8_24; // @[Switch.scala 30:36:@2659.4]
  wire  _T_20809; // @[Switch.scala 30:53:@2661.4]
  wire  valid_8_25; // @[Switch.scala 30:36:@2662.4]
  wire  _T_20812; // @[Switch.scala 30:53:@2664.4]
  wire  valid_8_26; // @[Switch.scala 30:36:@2665.4]
  wire  _T_20815; // @[Switch.scala 30:53:@2667.4]
  wire  valid_8_27; // @[Switch.scala 30:36:@2668.4]
  wire  _T_20818; // @[Switch.scala 30:53:@2670.4]
  wire  valid_8_28; // @[Switch.scala 30:36:@2671.4]
  wire  _T_20821; // @[Switch.scala 30:53:@2673.4]
  wire  valid_8_29; // @[Switch.scala 30:36:@2674.4]
  wire  _T_20824; // @[Switch.scala 30:53:@2676.4]
  wire  valid_8_30; // @[Switch.scala 30:36:@2677.4]
  wire  _T_20827; // @[Switch.scala 30:53:@2679.4]
  wire  valid_8_31; // @[Switch.scala 30:36:@2680.4]
  wire  _T_20830; // @[Switch.scala 30:53:@2682.4]
  wire  valid_8_32; // @[Switch.scala 30:36:@2683.4]
  wire  _T_20833; // @[Switch.scala 30:53:@2685.4]
  wire  valid_8_33; // @[Switch.scala 30:36:@2686.4]
  wire  _T_20836; // @[Switch.scala 30:53:@2688.4]
  wire  valid_8_34; // @[Switch.scala 30:36:@2689.4]
  wire  _T_20839; // @[Switch.scala 30:53:@2691.4]
  wire  valid_8_35; // @[Switch.scala 30:36:@2692.4]
  wire  _T_20842; // @[Switch.scala 30:53:@2694.4]
  wire  valid_8_36; // @[Switch.scala 30:36:@2695.4]
  wire  _T_20845; // @[Switch.scala 30:53:@2697.4]
  wire  valid_8_37; // @[Switch.scala 30:36:@2698.4]
  wire  _T_20848; // @[Switch.scala 30:53:@2700.4]
  wire  valid_8_38; // @[Switch.scala 30:36:@2701.4]
  wire  _T_20851; // @[Switch.scala 30:53:@2703.4]
  wire  valid_8_39; // @[Switch.scala 30:36:@2704.4]
  wire  _T_20854; // @[Switch.scala 30:53:@2706.4]
  wire  valid_8_40; // @[Switch.scala 30:36:@2707.4]
  wire  _T_20857; // @[Switch.scala 30:53:@2709.4]
  wire  valid_8_41; // @[Switch.scala 30:36:@2710.4]
  wire  _T_20860; // @[Switch.scala 30:53:@2712.4]
  wire  valid_8_42; // @[Switch.scala 30:36:@2713.4]
  wire  _T_20863; // @[Switch.scala 30:53:@2715.4]
  wire  valid_8_43; // @[Switch.scala 30:36:@2716.4]
  wire  _T_20866; // @[Switch.scala 30:53:@2718.4]
  wire  valid_8_44; // @[Switch.scala 30:36:@2719.4]
  wire  _T_20869; // @[Switch.scala 30:53:@2721.4]
  wire  valid_8_45; // @[Switch.scala 30:36:@2722.4]
  wire  _T_20872; // @[Switch.scala 30:53:@2724.4]
  wire  valid_8_46; // @[Switch.scala 30:36:@2725.4]
  wire  _T_20875; // @[Switch.scala 30:53:@2727.4]
  wire  valid_8_47; // @[Switch.scala 30:36:@2728.4]
  wire  _T_20878; // @[Switch.scala 30:53:@2730.4]
  wire  valid_8_48; // @[Switch.scala 30:36:@2731.4]
  wire  _T_20881; // @[Switch.scala 30:53:@2733.4]
  wire  valid_8_49; // @[Switch.scala 30:36:@2734.4]
  wire  _T_20884; // @[Switch.scala 30:53:@2736.4]
  wire  valid_8_50; // @[Switch.scala 30:36:@2737.4]
  wire  _T_20887; // @[Switch.scala 30:53:@2739.4]
  wire  valid_8_51; // @[Switch.scala 30:36:@2740.4]
  wire  _T_20890; // @[Switch.scala 30:53:@2742.4]
  wire  valid_8_52; // @[Switch.scala 30:36:@2743.4]
  wire  _T_20893; // @[Switch.scala 30:53:@2745.4]
  wire  valid_8_53; // @[Switch.scala 30:36:@2746.4]
  wire  _T_20896; // @[Switch.scala 30:53:@2748.4]
  wire  valid_8_54; // @[Switch.scala 30:36:@2749.4]
  wire  _T_20899; // @[Switch.scala 30:53:@2751.4]
  wire  valid_8_55; // @[Switch.scala 30:36:@2752.4]
  wire  _T_20902; // @[Switch.scala 30:53:@2754.4]
  wire  valid_8_56; // @[Switch.scala 30:36:@2755.4]
  wire  _T_20905; // @[Switch.scala 30:53:@2757.4]
  wire  valid_8_57; // @[Switch.scala 30:36:@2758.4]
  wire  _T_20908; // @[Switch.scala 30:53:@2760.4]
  wire  valid_8_58; // @[Switch.scala 30:36:@2761.4]
  wire  _T_20911; // @[Switch.scala 30:53:@2763.4]
  wire  valid_8_59; // @[Switch.scala 30:36:@2764.4]
  wire  _T_20914; // @[Switch.scala 30:53:@2766.4]
  wire  valid_8_60; // @[Switch.scala 30:36:@2767.4]
  wire  _T_20917; // @[Switch.scala 30:53:@2769.4]
  wire  valid_8_61; // @[Switch.scala 30:36:@2770.4]
  wire  _T_20920; // @[Switch.scala 30:53:@2772.4]
  wire  valid_8_62; // @[Switch.scala 30:36:@2773.4]
  wire  _T_20923; // @[Switch.scala 30:53:@2775.4]
  wire  valid_8_63; // @[Switch.scala 30:36:@2776.4]
  wire [5:0] _T_20989; // @[Mux.scala 31:69:@2778.4]
  wire [5:0] _T_20990; // @[Mux.scala 31:69:@2779.4]
  wire [5:0] _T_20991; // @[Mux.scala 31:69:@2780.4]
  wire [5:0] _T_20992; // @[Mux.scala 31:69:@2781.4]
  wire [5:0] _T_20993; // @[Mux.scala 31:69:@2782.4]
  wire [5:0] _T_20994; // @[Mux.scala 31:69:@2783.4]
  wire [5:0] _T_20995; // @[Mux.scala 31:69:@2784.4]
  wire [5:0] _T_20996; // @[Mux.scala 31:69:@2785.4]
  wire [5:0] _T_20997; // @[Mux.scala 31:69:@2786.4]
  wire [5:0] _T_20998; // @[Mux.scala 31:69:@2787.4]
  wire [5:0] _T_20999; // @[Mux.scala 31:69:@2788.4]
  wire [5:0] _T_21000; // @[Mux.scala 31:69:@2789.4]
  wire [5:0] _T_21001; // @[Mux.scala 31:69:@2790.4]
  wire [5:0] _T_21002; // @[Mux.scala 31:69:@2791.4]
  wire [5:0] _T_21003; // @[Mux.scala 31:69:@2792.4]
  wire [5:0] _T_21004; // @[Mux.scala 31:69:@2793.4]
  wire [5:0] _T_21005; // @[Mux.scala 31:69:@2794.4]
  wire [5:0] _T_21006; // @[Mux.scala 31:69:@2795.4]
  wire [5:0] _T_21007; // @[Mux.scala 31:69:@2796.4]
  wire [5:0] _T_21008; // @[Mux.scala 31:69:@2797.4]
  wire [5:0] _T_21009; // @[Mux.scala 31:69:@2798.4]
  wire [5:0] _T_21010; // @[Mux.scala 31:69:@2799.4]
  wire [5:0] _T_21011; // @[Mux.scala 31:69:@2800.4]
  wire [5:0] _T_21012; // @[Mux.scala 31:69:@2801.4]
  wire [5:0] _T_21013; // @[Mux.scala 31:69:@2802.4]
  wire [5:0] _T_21014; // @[Mux.scala 31:69:@2803.4]
  wire [5:0] _T_21015; // @[Mux.scala 31:69:@2804.4]
  wire [5:0] _T_21016; // @[Mux.scala 31:69:@2805.4]
  wire [5:0] _T_21017; // @[Mux.scala 31:69:@2806.4]
  wire [5:0] _T_21018; // @[Mux.scala 31:69:@2807.4]
  wire [5:0] _T_21019; // @[Mux.scala 31:69:@2808.4]
  wire [5:0] _T_21020; // @[Mux.scala 31:69:@2809.4]
  wire [5:0] _T_21021; // @[Mux.scala 31:69:@2810.4]
  wire [5:0] _T_21022; // @[Mux.scala 31:69:@2811.4]
  wire [5:0] _T_21023; // @[Mux.scala 31:69:@2812.4]
  wire [5:0] _T_21024; // @[Mux.scala 31:69:@2813.4]
  wire [5:0] _T_21025; // @[Mux.scala 31:69:@2814.4]
  wire [5:0] _T_21026; // @[Mux.scala 31:69:@2815.4]
  wire [5:0] _T_21027; // @[Mux.scala 31:69:@2816.4]
  wire [5:0] _T_21028; // @[Mux.scala 31:69:@2817.4]
  wire [5:0] _T_21029; // @[Mux.scala 31:69:@2818.4]
  wire [5:0] _T_21030; // @[Mux.scala 31:69:@2819.4]
  wire [5:0] _T_21031; // @[Mux.scala 31:69:@2820.4]
  wire [5:0] _T_21032; // @[Mux.scala 31:69:@2821.4]
  wire [5:0] _T_21033; // @[Mux.scala 31:69:@2822.4]
  wire [5:0] _T_21034; // @[Mux.scala 31:69:@2823.4]
  wire [5:0] _T_21035; // @[Mux.scala 31:69:@2824.4]
  wire [5:0] _T_21036; // @[Mux.scala 31:69:@2825.4]
  wire [5:0] _T_21037; // @[Mux.scala 31:69:@2826.4]
  wire [5:0] _T_21038; // @[Mux.scala 31:69:@2827.4]
  wire [5:0] _T_21039; // @[Mux.scala 31:69:@2828.4]
  wire [5:0] _T_21040; // @[Mux.scala 31:69:@2829.4]
  wire [5:0] _T_21041; // @[Mux.scala 31:69:@2830.4]
  wire [5:0] _T_21042; // @[Mux.scala 31:69:@2831.4]
  wire [5:0] _T_21043; // @[Mux.scala 31:69:@2832.4]
  wire [5:0] _T_21044; // @[Mux.scala 31:69:@2833.4]
  wire [5:0] _T_21045; // @[Mux.scala 31:69:@2834.4]
  wire [5:0] _T_21046; // @[Mux.scala 31:69:@2835.4]
  wire [5:0] _T_21047; // @[Mux.scala 31:69:@2836.4]
  wire [5:0] _T_21048; // @[Mux.scala 31:69:@2837.4]
  wire [5:0] _T_21049; // @[Mux.scala 31:69:@2838.4]
  wire [5:0] _T_21050; // @[Mux.scala 31:69:@2839.4]
  wire [5:0] select_8; // @[Mux.scala 31:69:@2840.4]
  wire [47:0] _GEN_513; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_514; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_515; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_516; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_517; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_518; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_519; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_520; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_521; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_522; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_523; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_524; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_525; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_526; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_527; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_528; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_529; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_530; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_531; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_532; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_533; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_534; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_535; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_536; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_537; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_538; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_539; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_540; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_541; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_542; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_543; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_544; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_545; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_546; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_547; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_548; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_549; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_550; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_551; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_552; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_553; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_554; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_555; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_556; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_557; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_558; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_559; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_560; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_561; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_562; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_563; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_564; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_565; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_566; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_567; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_568; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_569; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_570; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_571; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_572; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_573; // @[Switch.scala 33:19:@2842.4]
  wire [47:0] _GEN_574; // @[Switch.scala 33:19:@2842.4]
  wire [7:0] _T_21059; // @[Switch.scala 34:32:@2849.4]
  wire [15:0] _T_21067; // @[Switch.scala 34:32:@2857.4]
  wire [7:0] _T_21074; // @[Switch.scala 34:32:@2864.4]
  wire [31:0] _T_21083; // @[Switch.scala 34:32:@2873.4]
  wire [7:0] _T_21090; // @[Switch.scala 34:32:@2880.4]
  wire [15:0] _T_21098; // @[Switch.scala 34:32:@2888.4]
  wire [7:0] _T_21105; // @[Switch.scala 34:32:@2895.4]
  wire [31:0] _T_21114; // @[Switch.scala 34:32:@2904.4]
  wire [63:0] _T_21115; // @[Switch.scala 34:32:@2905.4]
  wire  _T_21119; // @[Switch.scala 30:53:@2908.4]
  wire  valid_9_0; // @[Switch.scala 30:36:@2909.4]
  wire  _T_21122; // @[Switch.scala 30:53:@2911.4]
  wire  valid_9_1; // @[Switch.scala 30:36:@2912.4]
  wire  _T_21125; // @[Switch.scala 30:53:@2914.4]
  wire  valid_9_2; // @[Switch.scala 30:36:@2915.4]
  wire  _T_21128; // @[Switch.scala 30:53:@2917.4]
  wire  valid_9_3; // @[Switch.scala 30:36:@2918.4]
  wire  _T_21131; // @[Switch.scala 30:53:@2920.4]
  wire  valid_9_4; // @[Switch.scala 30:36:@2921.4]
  wire  _T_21134; // @[Switch.scala 30:53:@2923.4]
  wire  valid_9_5; // @[Switch.scala 30:36:@2924.4]
  wire  _T_21137; // @[Switch.scala 30:53:@2926.4]
  wire  valid_9_6; // @[Switch.scala 30:36:@2927.4]
  wire  _T_21140; // @[Switch.scala 30:53:@2929.4]
  wire  valid_9_7; // @[Switch.scala 30:36:@2930.4]
  wire  _T_21143; // @[Switch.scala 30:53:@2932.4]
  wire  valid_9_8; // @[Switch.scala 30:36:@2933.4]
  wire  _T_21146; // @[Switch.scala 30:53:@2935.4]
  wire  valid_9_9; // @[Switch.scala 30:36:@2936.4]
  wire  _T_21149; // @[Switch.scala 30:53:@2938.4]
  wire  valid_9_10; // @[Switch.scala 30:36:@2939.4]
  wire  _T_21152; // @[Switch.scala 30:53:@2941.4]
  wire  valid_9_11; // @[Switch.scala 30:36:@2942.4]
  wire  _T_21155; // @[Switch.scala 30:53:@2944.4]
  wire  valid_9_12; // @[Switch.scala 30:36:@2945.4]
  wire  _T_21158; // @[Switch.scala 30:53:@2947.4]
  wire  valid_9_13; // @[Switch.scala 30:36:@2948.4]
  wire  _T_21161; // @[Switch.scala 30:53:@2950.4]
  wire  valid_9_14; // @[Switch.scala 30:36:@2951.4]
  wire  _T_21164; // @[Switch.scala 30:53:@2953.4]
  wire  valid_9_15; // @[Switch.scala 30:36:@2954.4]
  wire  _T_21167; // @[Switch.scala 30:53:@2956.4]
  wire  valid_9_16; // @[Switch.scala 30:36:@2957.4]
  wire  _T_21170; // @[Switch.scala 30:53:@2959.4]
  wire  valid_9_17; // @[Switch.scala 30:36:@2960.4]
  wire  _T_21173; // @[Switch.scala 30:53:@2962.4]
  wire  valid_9_18; // @[Switch.scala 30:36:@2963.4]
  wire  _T_21176; // @[Switch.scala 30:53:@2965.4]
  wire  valid_9_19; // @[Switch.scala 30:36:@2966.4]
  wire  _T_21179; // @[Switch.scala 30:53:@2968.4]
  wire  valid_9_20; // @[Switch.scala 30:36:@2969.4]
  wire  _T_21182; // @[Switch.scala 30:53:@2971.4]
  wire  valid_9_21; // @[Switch.scala 30:36:@2972.4]
  wire  _T_21185; // @[Switch.scala 30:53:@2974.4]
  wire  valid_9_22; // @[Switch.scala 30:36:@2975.4]
  wire  _T_21188; // @[Switch.scala 30:53:@2977.4]
  wire  valid_9_23; // @[Switch.scala 30:36:@2978.4]
  wire  _T_21191; // @[Switch.scala 30:53:@2980.4]
  wire  valid_9_24; // @[Switch.scala 30:36:@2981.4]
  wire  _T_21194; // @[Switch.scala 30:53:@2983.4]
  wire  valid_9_25; // @[Switch.scala 30:36:@2984.4]
  wire  _T_21197; // @[Switch.scala 30:53:@2986.4]
  wire  valid_9_26; // @[Switch.scala 30:36:@2987.4]
  wire  _T_21200; // @[Switch.scala 30:53:@2989.4]
  wire  valid_9_27; // @[Switch.scala 30:36:@2990.4]
  wire  _T_21203; // @[Switch.scala 30:53:@2992.4]
  wire  valid_9_28; // @[Switch.scala 30:36:@2993.4]
  wire  _T_21206; // @[Switch.scala 30:53:@2995.4]
  wire  valid_9_29; // @[Switch.scala 30:36:@2996.4]
  wire  _T_21209; // @[Switch.scala 30:53:@2998.4]
  wire  valid_9_30; // @[Switch.scala 30:36:@2999.4]
  wire  _T_21212; // @[Switch.scala 30:53:@3001.4]
  wire  valid_9_31; // @[Switch.scala 30:36:@3002.4]
  wire  _T_21215; // @[Switch.scala 30:53:@3004.4]
  wire  valid_9_32; // @[Switch.scala 30:36:@3005.4]
  wire  _T_21218; // @[Switch.scala 30:53:@3007.4]
  wire  valid_9_33; // @[Switch.scala 30:36:@3008.4]
  wire  _T_21221; // @[Switch.scala 30:53:@3010.4]
  wire  valid_9_34; // @[Switch.scala 30:36:@3011.4]
  wire  _T_21224; // @[Switch.scala 30:53:@3013.4]
  wire  valid_9_35; // @[Switch.scala 30:36:@3014.4]
  wire  _T_21227; // @[Switch.scala 30:53:@3016.4]
  wire  valid_9_36; // @[Switch.scala 30:36:@3017.4]
  wire  _T_21230; // @[Switch.scala 30:53:@3019.4]
  wire  valid_9_37; // @[Switch.scala 30:36:@3020.4]
  wire  _T_21233; // @[Switch.scala 30:53:@3022.4]
  wire  valid_9_38; // @[Switch.scala 30:36:@3023.4]
  wire  _T_21236; // @[Switch.scala 30:53:@3025.4]
  wire  valid_9_39; // @[Switch.scala 30:36:@3026.4]
  wire  _T_21239; // @[Switch.scala 30:53:@3028.4]
  wire  valid_9_40; // @[Switch.scala 30:36:@3029.4]
  wire  _T_21242; // @[Switch.scala 30:53:@3031.4]
  wire  valid_9_41; // @[Switch.scala 30:36:@3032.4]
  wire  _T_21245; // @[Switch.scala 30:53:@3034.4]
  wire  valid_9_42; // @[Switch.scala 30:36:@3035.4]
  wire  _T_21248; // @[Switch.scala 30:53:@3037.4]
  wire  valid_9_43; // @[Switch.scala 30:36:@3038.4]
  wire  _T_21251; // @[Switch.scala 30:53:@3040.4]
  wire  valid_9_44; // @[Switch.scala 30:36:@3041.4]
  wire  _T_21254; // @[Switch.scala 30:53:@3043.4]
  wire  valid_9_45; // @[Switch.scala 30:36:@3044.4]
  wire  _T_21257; // @[Switch.scala 30:53:@3046.4]
  wire  valid_9_46; // @[Switch.scala 30:36:@3047.4]
  wire  _T_21260; // @[Switch.scala 30:53:@3049.4]
  wire  valid_9_47; // @[Switch.scala 30:36:@3050.4]
  wire  _T_21263; // @[Switch.scala 30:53:@3052.4]
  wire  valid_9_48; // @[Switch.scala 30:36:@3053.4]
  wire  _T_21266; // @[Switch.scala 30:53:@3055.4]
  wire  valid_9_49; // @[Switch.scala 30:36:@3056.4]
  wire  _T_21269; // @[Switch.scala 30:53:@3058.4]
  wire  valid_9_50; // @[Switch.scala 30:36:@3059.4]
  wire  _T_21272; // @[Switch.scala 30:53:@3061.4]
  wire  valid_9_51; // @[Switch.scala 30:36:@3062.4]
  wire  _T_21275; // @[Switch.scala 30:53:@3064.4]
  wire  valid_9_52; // @[Switch.scala 30:36:@3065.4]
  wire  _T_21278; // @[Switch.scala 30:53:@3067.4]
  wire  valid_9_53; // @[Switch.scala 30:36:@3068.4]
  wire  _T_21281; // @[Switch.scala 30:53:@3070.4]
  wire  valid_9_54; // @[Switch.scala 30:36:@3071.4]
  wire  _T_21284; // @[Switch.scala 30:53:@3073.4]
  wire  valid_9_55; // @[Switch.scala 30:36:@3074.4]
  wire  _T_21287; // @[Switch.scala 30:53:@3076.4]
  wire  valid_9_56; // @[Switch.scala 30:36:@3077.4]
  wire  _T_21290; // @[Switch.scala 30:53:@3079.4]
  wire  valid_9_57; // @[Switch.scala 30:36:@3080.4]
  wire  _T_21293; // @[Switch.scala 30:53:@3082.4]
  wire  valid_9_58; // @[Switch.scala 30:36:@3083.4]
  wire  _T_21296; // @[Switch.scala 30:53:@3085.4]
  wire  valid_9_59; // @[Switch.scala 30:36:@3086.4]
  wire  _T_21299; // @[Switch.scala 30:53:@3088.4]
  wire  valid_9_60; // @[Switch.scala 30:36:@3089.4]
  wire  _T_21302; // @[Switch.scala 30:53:@3091.4]
  wire  valid_9_61; // @[Switch.scala 30:36:@3092.4]
  wire  _T_21305; // @[Switch.scala 30:53:@3094.4]
  wire  valid_9_62; // @[Switch.scala 30:36:@3095.4]
  wire  _T_21308; // @[Switch.scala 30:53:@3097.4]
  wire  valid_9_63; // @[Switch.scala 30:36:@3098.4]
  wire [5:0] _T_21374; // @[Mux.scala 31:69:@3100.4]
  wire [5:0] _T_21375; // @[Mux.scala 31:69:@3101.4]
  wire [5:0] _T_21376; // @[Mux.scala 31:69:@3102.4]
  wire [5:0] _T_21377; // @[Mux.scala 31:69:@3103.4]
  wire [5:0] _T_21378; // @[Mux.scala 31:69:@3104.4]
  wire [5:0] _T_21379; // @[Mux.scala 31:69:@3105.4]
  wire [5:0] _T_21380; // @[Mux.scala 31:69:@3106.4]
  wire [5:0] _T_21381; // @[Mux.scala 31:69:@3107.4]
  wire [5:0] _T_21382; // @[Mux.scala 31:69:@3108.4]
  wire [5:0] _T_21383; // @[Mux.scala 31:69:@3109.4]
  wire [5:0] _T_21384; // @[Mux.scala 31:69:@3110.4]
  wire [5:0] _T_21385; // @[Mux.scala 31:69:@3111.4]
  wire [5:0] _T_21386; // @[Mux.scala 31:69:@3112.4]
  wire [5:0] _T_21387; // @[Mux.scala 31:69:@3113.4]
  wire [5:0] _T_21388; // @[Mux.scala 31:69:@3114.4]
  wire [5:0] _T_21389; // @[Mux.scala 31:69:@3115.4]
  wire [5:0] _T_21390; // @[Mux.scala 31:69:@3116.4]
  wire [5:0] _T_21391; // @[Mux.scala 31:69:@3117.4]
  wire [5:0] _T_21392; // @[Mux.scala 31:69:@3118.4]
  wire [5:0] _T_21393; // @[Mux.scala 31:69:@3119.4]
  wire [5:0] _T_21394; // @[Mux.scala 31:69:@3120.4]
  wire [5:0] _T_21395; // @[Mux.scala 31:69:@3121.4]
  wire [5:0] _T_21396; // @[Mux.scala 31:69:@3122.4]
  wire [5:0] _T_21397; // @[Mux.scala 31:69:@3123.4]
  wire [5:0] _T_21398; // @[Mux.scala 31:69:@3124.4]
  wire [5:0] _T_21399; // @[Mux.scala 31:69:@3125.4]
  wire [5:0] _T_21400; // @[Mux.scala 31:69:@3126.4]
  wire [5:0] _T_21401; // @[Mux.scala 31:69:@3127.4]
  wire [5:0] _T_21402; // @[Mux.scala 31:69:@3128.4]
  wire [5:0] _T_21403; // @[Mux.scala 31:69:@3129.4]
  wire [5:0] _T_21404; // @[Mux.scala 31:69:@3130.4]
  wire [5:0] _T_21405; // @[Mux.scala 31:69:@3131.4]
  wire [5:0] _T_21406; // @[Mux.scala 31:69:@3132.4]
  wire [5:0] _T_21407; // @[Mux.scala 31:69:@3133.4]
  wire [5:0] _T_21408; // @[Mux.scala 31:69:@3134.4]
  wire [5:0] _T_21409; // @[Mux.scala 31:69:@3135.4]
  wire [5:0] _T_21410; // @[Mux.scala 31:69:@3136.4]
  wire [5:0] _T_21411; // @[Mux.scala 31:69:@3137.4]
  wire [5:0] _T_21412; // @[Mux.scala 31:69:@3138.4]
  wire [5:0] _T_21413; // @[Mux.scala 31:69:@3139.4]
  wire [5:0] _T_21414; // @[Mux.scala 31:69:@3140.4]
  wire [5:0] _T_21415; // @[Mux.scala 31:69:@3141.4]
  wire [5:0] _T_21416; // @[Mux.scala 31:69:@3142.4]
  wire [5:0] _T_21417; // @[Mux.scala 31:69:@3143.4]
  wire [5:0] _T_21418; // @[Mux.scala 31:69:@3144.4]
  wire [5:0] _T_21419; // @[Mux.scala 31:69:@3145.4]
  wire [5:0] _T_21420; // @[Mux.scala 31:69:@3146.4]
  wire [5:0] _T_21421; // @[Mux.scala 31:69:@3147.4]
  wire [5:0] _T_21422; // @[Mux.scala 31:69:@3148.4]
  wire [5:0] _T_21423; // @[Mux.scala 31:69:@3149.4]
  wire [5:0] _T_21424; // @[Mux.scala 31:69:@3150.4]
  wire [5:0] _T_21425; // @[Mux.scala 31:69:@3151.4]
  wire [5:0] _T_21426; // @[Mux.scala 31:69:@3152.4]
  wire [5:0] _T_21427; // @[Mux.scala 31:69:@3153.4]
  wire [5:0] _T_21428; // @[Mux.scala 31:69:@3154.4]
  wire [5:0] _T_21429; // @[Mux.scala 31:69:@3155.4]
  wire [5:0] _T_21430; // @[Mux.scala 31:69:@3156.4]
  wire [5:0] _T_21431; // @[Mux.scala 31:69:@3157.4]
  wire [5:0] _T_21432; // @[Mux.scala 31:69:@3158.4]
  wire [5:0] _T_21433; // @[Mux.scala 31:69:@3159.4]
  wire [5:0] _T_21434; // @[Mux.scala 31:69:@3160.4]
  wire [5:0] _T_21435; // @[Mux.scala 31:69:@3161.4]
  wire [5:0] select_9; // @[Mux.scala 31:69:@3162.4]
  wire [47:0] _GEN_577; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_578; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_579; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_580; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_581; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_582; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_583; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_584; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_585; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_586; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_587; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_588; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_589; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_590; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_591; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_592; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_593; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_594; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_595; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_596; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_597; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_598; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_599; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_600; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_601; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_602; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_603; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_604; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_605; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_606; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_607; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_608; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_609; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_610; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_611; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_612; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_613; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_614; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_615; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_616; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_617; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_618; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_619; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_620; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_621; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_622; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_623; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_624; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_625; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_626; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_627; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_628; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_629; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_630; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_631; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_632; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_633; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_634; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_635; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_636; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_637; // @[Switch.scala 33:19:@3164.4]
  wire [47:0] _GEN_638; // @[Switch.scala 33:19:@3164.4]
  wire [7:0] _T_21444; // @[Switch.scala 34:32:@3171.4]
  wire [15:0] _T_21452; // @[Switch.scala 34:32:@3179.4]
  wire [7:0] _T_21459; // @[Switch.scala 34:32:@3186.4]
  wire [31:0] _T_21468; // @[Switch.scala 34:32:@3195.4]
  wire [7:0] _T_21475; // @[Switch.scala 34:32:@3202.4]
  wire [15:0] _T_21483; // @[Switch.scala 34:32:@3210.4]
  wire [7:0] _T_21490; // @[Switch.scala 34:32:@3217.4]
  wire [31:0] _T_21499; // @[Switch.scala 34:32:@3226.4]
  wire [63:0] _T_21500; // @[Switch.scala 34:32:@3227.4]
  wire  _T_21504; // @[Switch.scala 30:53:@3230.4]
  wire  valid_10_0; // @[Switch.scala 30:36:@3231.4]
  wire  _T_21507; // @[Switch.scala 30:53:@3233.4]
  wire  valid_10_1; // @[Switch.scala 30:36:@3234.4]
  wire  _T_21510; // @[Switch.scala 30:53:@3236.4]
  wire  valid_10_2; // @[Switch.scala 30:36:@3237.4]
  wire  _T_21513; // @[Switch.scala 30:53:@3239.4]
  wire  valid_10_3; // @[Switch.scala 30:36:@3240.4]
  wire  _T_21516; // @[Switch.scala 30:53:@3242.4]
  wire  valid_10_4; // @[Switch.scala 30:36:@3243.4]
  wire  _T_21519; // @[Switch.scala 30:53:@3245.4]
  wire  valid_10_5; // @[Switch.scala 30:36:@3246.4]
  wire  _T_21522; // @[Switch.scala 30:53:@3248.4]
  wire  valid_10_6; // @[Switch.scala 30:36:@3249.4]
  wire  _T_21525; // @[Switch.scala 30:53:@3251.4]
  wire  valid_10_7; // @[Switch.scala 30:36:@3252.4]
  wire  _T_21528; // @[Switch.scala 30:53:@3254.4]
  wire  valid_10_8; // @[Switch.scala 30:36:@3255.4]
  wire  _T_21531; // @[Switch.scala 30:53:@3257.4]
  wire  valid_10_9; // @[Switch.scala 30:36:@3258.4]
  wire  _T_21534; // @[Switch.scala 30:53:@3260.4]
  wire  valid_10_10; // @[Switch.scala 30:36:@3261.4]
  wire  _T_21537; // @[Switch.scala 30:53:@3263.4]
  wire  valid_10_11; // @[Switch.scala 30:36:@3264.4]
  wire  _T_21540; // @[Switch.scala 30:53:@3266.4]
  wire  valid_10_12; // @[Switch.scala 30:36:@3267.4]
  wire  _T_21543; // @[Switch.scala 30:53:@3269.4]
  wire  valid_10_13; // @[Switch.scala 30:36:@3270.4]
  wire  _T_21546; // @[Switch.scala 30:53:@3272.4]
  wire  valid_10_14; // @[Switch.scala 30:36:@3273.4]
  wire  _T_21549; // @[Switch.scala 30:53:@3275.4]
  wire  valid_10_15; // @[Switch.scala 30:36:@3276.4]
  wire  _T_21552; // @[Switch.scala 30:53:@3278.4]
  wire  valid_10_16; // @[Switch.scala 30:36:@3279.4]
  wire  _T_21555; // @[Switch.scala 30:53:@3281.4]
  wire  valid_10_17; // @[Switch.scala 30:36:@3282.4]
  wire  _T_21558; // @[Switch.scala 30:53:@3284.4]
  wire  valid_10_18; // @[Switch.scala 30:36:@3285.4]
  wire  _T_21561; // @[Switch.scala 30:53:@3287.4]
  wire  valid_10_19; // @[Switch.scala 30:36:@3288.4]
  wire  _T_21564; // @[Switch.scala 30:53:@3290.4]
  wire  valid_10_20; // @[Switch.scala 30:36:@3291.4]
  wire  _T_21567; // @[Switch.scala 30:53:@3293.4]
  wire  valid_10_21; // @[Switch.scala 30:36:@3294.4]
  wire  _T_21570; // @[Switch.scala 30:53:@3296.4]
  wire  valid_10_22; // @[Switch.scala 30:36:@3297.4]
  wire  _T_21573; // @[Switch.scala 30:53:@3299.4]
  wire  valid_10_23; // @[Switch.scala 30:36:@3300.4]
  wire  _T_21576; // @[Switch.scala 30:53:@3302.4]
  wire  valid_10_24; // @[Switch.scala 30:36:@3303.4]
  wire  _T_21579; // @[Switch.scala 30:53:@3305.4]
  wire  valid_10_25; // @[Switch.scala 30:36:@3306.4]
  wire  _T_21582; // @[Switch.scala 30:53:@3308.4]
  wire  valid_10_26; // @[Switch.scala 30:36:@3309.4]
  wire  _T_21585; // @[Switch.scala 30:53:@3311.4]
  wire  valid_10_27; // @[Switch.scala 30:36:@3312.4]
  wire  _T_21588; // @[Switch.scala 30:53:@3314.4]
  wire  valid_10_28; // @[Switch.scala 30:36:@3315.4]
  wire  _T_21591; // @[Switch.scala 30:53:@3317.4]
  wire  valid_10_29; // @[Switch.scala 30:36:@3318.4]
  wire  _T_21594; // @[Switch.scala 30:53:@3320.4]
  wire  valid_10_30; // @[Switch.scala 30:36:@3321.4]
  wire  _T_21597; // @[Switch.scala 30:53:@3323.4]
  wire  valid_10_31; // @[Switch.scala 30:36:@3324.4]
  wire  _T_21600; // @[Switch.scala 30:53:@3326.4]
  wire  valid_10_32; // @[Switch.scala 30:36:@3327.4]
  wire  _T_21603; // @[Switch.scala 30:53:@3329.4]
  wire  valid_10_33; // @[Switch.scala 30:36:@3330.4]
  wire  _T_21606; // @[Switch.scala 30:53:@3332.4]
  wire  valid_10_34; // @[Switch.scala 30:36:@3333.4]
  wire  _T_21609; // @[Switch.scala 30:53:@3335.4]
  wire  valid_10_35; // @[Switch.scala 30:36:@3336.4]
  wire  _T_21612; // @[Switch.scala 30:53:@3338.4]
  wire  valid_10_36; // @[Switch.scala 30:36:@3339.4]
  wire  _T_21615; // @[Switch.scala 30:53:@3341.4]
  wire  valid_10_37; // @[Switch.scala 30:36:@3342.4]
  wire  _T_21618; // @[Switch.scala 30:53:@3344.4]
  wire  valid_10_38; // @[Switch.scala 30:36:@3345.4]
  wire  _T_21621; // @[Switch.scala 30:53:@3347.4]
  wire  valid_10_39; // @[Switch.scala 30:36:@3348.4]
  wire  _T_21624; // @[Switch.scala 30:53:@3350.4]
  wire  valid_10_40; // @[Switch.scala 30:36:@3351.4]
  wire  _T_21627; // @[Switch.scala 30:53:@3353.4]
  wire  valid_10_41; // @[Switch.scala 30:36:@3354.4]
  wire  _T_21630; // @[Switch.scala 30:53:@3356.4]
  wire  valid_10_42; // @[Switch.scala 30:36:@3357.4]
  wire  _T_21633; // @[Switch.scala 30:53:@3359.4]
  wire  valid_10_43; // @[Switch.scala 30:36:@3360.4]
  wire  _T_21636; // @[Switch.scala 30:53:@3362.4]
  wire  valid_10_44; // @[Switch.scala 30:36:@3363.4]
  wire  _T_21639; // @[Switch.scala 30:53:@3365.4]
  wire  valid_10_45; // @[Switch.scala 30:36:@3366.4]
  wire  _T_21642; // @[Switch.scala 30:53:@3368.4]
  wire  valid_10_46; // @[Switch.scala 30:36:@3369.4]
  wire  _T_21645; // @[Switch.scala 30:53:@3371.4]
  wire  valid_10_47; // @[Switch.scala 30:36:@3372.4]
  wire  _T_21648; // @[Switch.scala 30:53:@3374.4]
  wire  valid_10_48; // @[Switch.scala 30:36:@3375.4]
  wire  _T_21651; // @[Switch.scala 30:53:@3377.4]
  wire  valid_10_49; // @[Switch.scala 30:36:@3378.4]
  wire  _T_21654; // @[Switch.scala 30:53:@3380.4]
  wire  valid_10_50; // @[Switch.scala 30:36:@3381.4]
  wire  _T_21657; // @[Switch.scala 30:53:@3383.4]
  wire  valid_10_51; // @[Switch.scala 30:36:@3384.4]
  wire  _T_21660; // @[Switch.scala 30:53:@3386.4]
  wire  valid_10_52; // @[Switch.scala 30:36:@3387.4]
  wire  _T_21663; // @[Switch.scala 30:53:@3389.4]
  wire  valid_10_53; // @[Switch.scala 30:36:@3390.4]
  wire  _T_21666; // @[Switch.scala 30:53:@3392.4]
  wire  valid_10_54; // @[Switch.scala 30:36:@3393.4]
  wire  _T_21669; // @[Switch.scala 30:53:@3395.4]
  wire  valid_10_55; // @[Switch.scala 30:36:@3396.4]
  wire  _T_21672; // @[Switch.scala 30:53:@3398.4]
  wire  valid_10_56; // @[Switch.scala 30:36:@3399.4]
  wire  _T_21675; // @[Switch.scala 30:53:@3401.4]
  wire  valid_10_57; // @[Switch.scala 30:36:@3402.4]
  wire  _T_21678; // @[Switch.scala 30:53:@3404.4]
  wire  valid_10_58; // @[Switch.scala 30:36:@3405.4]
  wire  _T_21681; // @[Switch.scala 30:53:@3407.4]
  wire  valid_10_59; // @[Switch.scala 30:36:@3408.4]
  wire  _T_21684; // @[Switch.scala 30:53:@3410.4]
  wire  valid_10_60; // @[Switch.scala 30:36:@3411.4]
  wire  _T_21687; // @[Switch.scala 30:53:@3413.4]
  wire  valid_10_61; // @[Switch.scala 30:36:@3414.4]
  wire  _T_21690; // @[Switch.scala 30:53:@3416.4]
  wire  valid_10_62; // @[Switch.scala 30:36:@3417.4]
  wire  _T_21693; // @[Switch.scala 30:53:@3419.4]
  wire  valid_10_63; // @[Switch.scala 30:36:@3420.4]
  wire [5:0] _T_21759; // @[Mux.scala 31:69:@3422.4]
  wire [5:0] _T_21760; // @[Mux.scala 31:69:@3423.4]
  wire [5:0] _T_21761; // @[Mux.scala 31:69:@3424.4]
  wire [5:0] _T_21762; // @[Mux.scala 31:69:@3425.4]
  wire [5:0] _T_21763; // @[Mux.scala 31:69:@3426.4]
  wire [5:0] _T_21764; // @[Mux.scala 31:69:@3427.4]
  wire [5:0] _T_21765; // @[Mux.scala 31:69:@3428.4]
  wire [5:0] _T_21766; // @[Mux.scala 31:69:@3429.4]
  wire [5:0] _T_21767; // @[Mux.scala 31:69:@3430.4]
  wire [5:0] _T_21768; // @[Mux.scala 31:69:@3431.4]
  wire [5:0] _T_21769; // @[Mux.scala 31:69:@3432.4]
  wire [5:0] _T_21770; // @[Mux.scala 31:69:@3433.4]
  wire [5:0] _T_21771; // @[Mux.scala 31:69:@3434.4]
  wire [5:0] _T_21772; // @[Mux.scala 31:69:@3435.4]
  wire [5:0] _T_21773; // @[Mux.scala 31:69:@3436.4]
  wire [5:0] _T_21774; // @[Mux.scala 31:69:@3437.4]
  wire [5:0] _T_21775; // @[Mux.scala 31:69:@3438.4]
  wire [5:0] _T_21776; // @[Mux.scala 31:69:@3439.4]
  wire [5:0] _T_21777; // @[Mux.scala 31:69:@3440.4]
  wire [5:0] _T_21778; // @[Mux.scala 31:69:@3441.4]
  wire [5:0] _T_21779; // @[Mux.scala 31:69:@3442.4]
  wire [5:0] _T_21780; // @[Mux.scala 31:69:@3443.4]
  wire [5:0] _T_21781; // @[Mux.scala 31:69:@3444.4]
  wire [5:0] _T_21782; // @[Mux.scala 31:69:@3445.4]
  wire [5:0] _T_21783; // @[Mux.scala 31:69:@3446.4]
  wire [5:0] _T_21784; // @[Mux.scala 31:69:@3447.4]
  wire [5:0] _T_21785; // @[Mux.scala 31:69:@3448.4]
  wire [5:0] _T_21786; // @[Mux.scala 31:69:@3449.4]
  wire [5:0] _T_21787; // @[Mux.scala 31:69:@3450.4]
  wire [5:0] _T_21788; // @[Mux.scala 31:69:@3451.4]
  wire [5:0] _T_21789; // @[Mux.scala 31:69:@3452.4]
  wire [5:0] _T_21790; // @[Mux.scala 31:69:@3453.4]
  wire [5:0] _T_21791; // @[Mux.scala 31:69:@3454.4]
  wire [5:0] _T_21792; // @[Mux.scala 31:69:@3455.4]
  wire [5:0] _T_21793; // @[Mux.scala 31:69:@3456.4]
  wire [5:0] _T_21794; // @[Mux.scala 31:69:@3457.4]
  wire [5:0] _T_21795; // @[Mux.scala 31:69:@3458.4]
  wire [5:0] _T_21796; // @[Mux.scala 31:69:@3459.4]
  wire [5:0] _T_21797; // @[Mux.scala 31:69:@3460.4]
  wire [5:0] _T_21798; // @[Mux.scala 31:69:@3461.4]
  wire [5:0] _T_21799; // @[Mux.scala 31:69:@3462.4]
  wire [5:0] _T_21800; // @[Mux.scala 31:69:@3463.4]
  wire [5:0] _T_21801; // @[Mux.scala 31:69:@3464.4]
  wire [5:0] _T_21802; // @[Mux.scala 31:69:@3465.4]
  wire [5:0] _T_21803; // @[Mux.scala 31:69:@3466.4]
  wire [5:0] _T_21804; // @[Mux.scala 31:69:@3467.4]
  wire [5:0] _T_21805; // @[Mux.scala 31:69:@3468.4]
  wire [5:0] _T_21806; // @[Mux.scala 31:69:@3469.4]
  wire [5:0] _T_21807; // @[Mux.scala 31:69:@3470.4]
  wire [5:0] _T_21808; // @[Mux.scala 31:69:@3471.4]
  wire [5:0] _T_21809; // @[Mux.scala 31:69:@3472.4]
  wire [5:0] _T_21810; // @[Mux.scala 31:69:@3473.4]
  wire [5:0] _T_21811; // @[Mux.scala 31:69:@3474.4]
  wire [5:0] _T_21812; // @[Mux.scala 31:69:@3475.4]
  wire [5:0] _T_21813; // @[Mux.scala 31:69:@3476.4]
  wire [5:0] _T_21814; // @[Mux.scala 31:69:@3477.4]
  wire [5:0] _T_21815; // @[Mux.scala 31:69:@3478.4]
  wire [5:0] _T_21816; // @[Mux.scala 31:69:@3479.4]
  wire [5:0] _T_21817; // @[Mux.scala 31:69:@3480.4]
  wire [5:0] _T_21818; // @[Mux.scala 31:69:@3481.4]
  wire [5:0] _T_21819; // @[Mux.scala 31:69:@3482.4]
  wire [5:0] _T_21820; // @[Mux.scala 31:69:@3483.4]
  wire [5:0] select_10; // @[Mux.scala 31:69:@3484.4]
  wire [47:0] _GEN_641; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_642; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_643; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_644; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_645; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_646; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_647; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_648; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_649; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_650; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_651; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_652; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_653; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_654; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_655; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_656; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_657; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_658; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_659; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_660; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_661; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_662; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_663; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_664; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_665; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_666; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_667; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_668; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_669; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_670; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_671; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_672; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_673; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_674; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_675; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_676; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_677; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_678; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_679; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_680; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_681; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_682; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_683; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_684; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_685; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_686; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_687; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_688; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_689; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_690; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_691; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_692; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_693; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_694; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_695; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_696; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_697; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_698; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_699; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_700; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_701; // @[Switch.scala 33:19:@3486.4]
  wire [47:0] _GEN_702; // @[Switch.scala 33:19:@3486.4]
  wire [7:0] _T_21829; // @[Switch.scala 34:32:@3493.4]
  wire [15:0] _T_21837; // @[Switch.scala 34:32:@3501.4]
  wire [7:0] _T_21844; // @[Switch.scala 34:32:@3508.4]
  wire [31:0] _T_21853; // @[Switch.scala 34:32:@3517.4]
  wire [7:0] _T_21860; // @[Switch.scala 34:32:@3524.4]
  wire [15:0] _T_21868; // @[Switch.scala 34:32:@3532.4]
  wire [7:0] _T_21875; // @[Switch.scala 34:32:@3539.4]
  wire [31:0] _T_21884; // @[Switch.scala 34:32:@3548.4]
  wire [63:0] _T_21885; // @[Switch.scala 34:32:@3549.4]
  wire  _T_21889; // @[Switch.scala 30:53:@3552.4]
  wire  valid_11_0; // @[Switch.scala 30:36:@3553.4]
  wire  _T_21892; // @[Switch.scala 30:53:@3555.4]
  wire  valid_11_1; // @[Switch.scala 30:36:@3556.4]
  wire  _T_21895; // @[Switch.scala 30:53:@3558.4]
  wire  valid_11_2; // @[Switch.scala 30:36:@3559.4]
  wire  _T_21898; // @[Switch.scala 30:53:@3561.4]
  wire  valid_11_3; // @[Switch.scala 30:36:@3562.4]
  wire  _T_21901; // @[Switch.scala 30:53:@3564.4]
  wire  valid_11_4; // @[Switch.scala 30:36:@3565.4]
  wire  _T_21904; // @[Switch.scala 30:53:@3567.4]
  wire  valid_11_5; // @[Switch.scala 30:36:@3568.4]
  wire  _T_21907; // @[Switch.scala 30:53:@3570.4]
  wire  valid_11_6; // @[Switch.scala 30:36:@3571.4]
  wire  _T_21910; // @[Switch.scala 30:53:@3573.4]
  wire  valid_11_7; // @[Switch.scala 30:36:@3574.4]
  wire  _T_21913; // @[Switch.scala 30:53:@3576.4]
  wire  valid_11_8; // @[Switch.scala 30:36:@3577.4]
  wire  _T_21916; // @[Switch.scala 30:53:@3579.4]
  wire  valid_11_9; // @[Switch.scala 30:36:@3580.4]
  wire  _T_21919; // @[Switch.scala 30:53:@3582.4]
  wire  valid_11_10; // @[Switch.scala 30:36:@3583.4]
  wire  _T_21922; // @[Switch.scala 30:53:@3585.4]
  wire  valid_11_11; // @[Switch.scala 30:36:@3586.4]
  wire  _T_21925; // @[Switch.scala 30:53:@3588.4]
  wire  valid_11_12; // @[Switch.scala 30:36:@3589.4]
  wire  _T_21928; // @[Switch.scala 30:53:@3591.4]
  wire  valid_11_13; // @[Switch.scala 30:36:@3592.4]
  wire  _T_21931; // @[Switch.scala 30:53:@3594.4]
  wire  valid_11_14; // @[Switch.scala 30:36:@3595.4]
  wire  _T_21934; // @[Switch.scala 30:53:@3597.4]
  wire  valid_11_15; // @[Switch.scala 30:36:@3598.4]
  wire  _T_21937; // @[Switch.scala 30:53:@3600.4]
  wire  valid_11_16; // @[Switch.scala 30:36:@3601.4]
  wire  _T_21940; // @[Switch.scala 30:53:@3603.4]
  wire  valid_11_17; // @[Switch.scala 30:36:@3604.4]
  wire  _T_21943; // @[Switch.scala 30:53:@3606.4]
  wire  valid_11_18; // @[Switch.scala 30:36:@3607.4]
  wire  _T_21946; // @[Switch.scala 30:53:@3609.4]
  wire  valid_11_19; // @[Switch.scala 30:36:@3610.4]
  wire  _T_21949; // @[Switch.scala 30:53:@3612.4]
  wire  valid_11_20; // @[Switch.scala 30:36:@3613.4]
  wire  _T_21952; // @[Switch.scala 30:53:@3615.4]
  wire  valid_11_21; // @[Switch.scala 30:36:@3616.4]
  wire  _T_21955; // @[Switch.scala 30:53:@3618.4]
  wire  valid_11_22; // @[Switch.scala 30:36:@3619.4]
  wire  _T_21958; // @[Switch.scala 30:53:@3621.4]
  wire  valid_11_23; // @[Switch.scala 30:36:@3622.4]
  wire  _T_21961; // @[Switch.scala 30:53:@3624.4]
  wire  valid_11_24; // @[Switch.scala 30:36:@3625.4]
  wire  _T_21964; // @[Switch.scala 30:53:@3627.4]
  wire  valid_11_25; // @[Switch.scala 30:36:@3628.4]
  wire  _T_21967; // @[Switch.scala 30:53:@3630.4]
  wire  valid_11_26; // @[Switch.scala 30:36:@3631.4]
  wire  _T_21970; // @[Switch.scala 30:53:@3633.4]
  wire  valid_11_27; // @[Switch.scala 30:36:@3634.4]
  wire  _T_21973; // @[Switch.scala 30:53:@3636.4]
  wire  valid_11_28; // @[Switch.scala 30:36:@3637.4]
  wire  _T_21976; // @[Switch.scala 30:53:@3639.4]
  wire  valid_11_29; // @[Switch.scala 30:36:@3640.4]
  wire  _T_21979; // @[Switch.scala 30:53:@3642.4]
  wire  valid_11_30; // @[Switch.scala 30:36:@3643.4]
  wire  _T_21982; // @[Switch.scala 30:53:@3645.4]
  wire  valid_11_31; // @[Switch.scala 30:36:@3646.4]
  wire  _T_21985; // @[Switch.scala 30:53:@3648.4]
  wire  valid_11_32; // @[Switch.scala 30:36:@3649.4]
  wire  _T_21988; // @[Switch.scala 30:53:@3651.4]
  wire  valid_11_33; // @[Switch.scala 30:36:@3652.4]
  wire  _T_21991; // @[Switch.scala 30:53:@3654.4]
  wire  valid_11_34; // @[Switch.scala 30:36:@3655.4]
  wire  _T_21994; // @[Switch.scala 30:53:@3657.4]
  wire  valid_11_35; // @[Switch.scala 30:36:@3658.4]
  wire  _T_21997; // @[Switch.scala 30:53:@3660.4]
  wire  valid_11_36; // @[Switch.scala 30:36:@3661.4]
  wire  _T_22000; // @[Switch.scala 30:53:@3663.4]
  wire  valid_11_37; // @[Switch.scala 30:36:@3664.4]
  wire  _T_22003; // @[Switch.scala 30:53:@3666.4]
  wire  valid_11_38; // @[Switch.scala 30:36:@3667.4]
  wire  _T_22006; // @[Switch.scala 30:53:@3669.4]
  wire  valid_11_39; // @[Switch.scala 30:36:@3670.4]
  wire  _T_22009; // @[Switch.scala 30:53:@3672.4]
  wire  valid_11_40; // @[Switch.scala 30:36:@3673.4]
  wire  _T_22012; // @[Switch.scala 30:53:@3675.4]
  wire  valid_11_41; // @[Switch.scala 30:36:@3676.4]
  wire  _T_22015; // @[Switch.scala 30:53:@3678.4]
  wire  valid_11_42; // @[Switch.scala 30:36:@3679.4]
  wire  _T_22018; // @[Switch.scala 30:53:@3681.4]
  wire  valid_11_43; // @[Switch.scala 30:36:@3682.4]
  wire  _T_22021; // @[Switch.scala 30:53:@3684.4]
  wire  valid_11_44; // @[Switch.scala 30:36:@3685.4]
  wire  _T_22024; // @[Switch.scala 30:53:@3687.4]
  wire  valid_11_45; // @[Switch.scala 30:36:@3688.4]
  wire  _T_22027; // @[Switch.scala 30:53:@3690.4]
  wire  valid_11_46; // @[Switch.scala 30:36:@3691.4]
  wire  _T_22030; // @[Switch.scala 30:53:@3693.4]
  wire  valid_11_47; // @[Switch.scala 30:36:@3694.4]
  wire  _T_22033; // @[Switch.scala 30:53:@3696.4]
  wire  valid_11_48; // @[Switch.scala 30:36:@3697.4]
  wire  _T_22036; // @[Switch.scala 30:53:@3699.4]
  wire  valid_11_49; // @[Switch.scala 30:36:@3700.4]
  wire  _T_22039; // @[Switch.scala 30:53:@3702.4]
  wire  valid_11_50; // @[Switch.scala 30:36:@3703.4]
  wire  _T_22042; // @[Switch.scala 30:53:@3705.4]
  wire  valid_11_51; // @[Switch.scala 30:36:@3706.4]
  wire  _T_22045; // @[Switch.scala 30:53:@3708.4]
  wire  valid_11_52; // @[Switch.scala 30:36:@3709.4]
  wire  _T_22048; // @[Switch.scala 30:53:@3711.4]
  wire  valid_11_53; // @[Switch.scala 30:36:@3712.4]
  wire  _T_22051; // @[Switch.scala 30:53:@3714.4]
  wire  valid_11_54; // @[Switch.scala 30:36:@3715.4]
  wire  _T_22054; // @[Switch.scala 30:53:@3717.4]
  wire  valid_11_55; // @[Switch.scala 30:36:@3718.4]
  wire  _T_22057; // @[Switch.scala 30:53:@3720.4]
  wire  valid_11_56; // @[Switch.scala 30:36:@3721.4]
  wire  _T_22060; // @[Switch.scala 30:53:@3723.4]
  wire  valid_11_57; // @[Switch.scala 30:36:@3724.4]
  wire  _T_22063; // @[Switch.scala 30:53:@3726.4]
  wire  valid_11_58; // @[Switch.scala 30:36:@3727.4]
  wire  _T_22066; // @[Switch.scala 30:53:@3729.4]
  wire  valid_11_59; // @[Switch.scala 30:36:@3730.4]
  wire  _T_22069; // @[Switch.scala 30:53:@3732.4]
  wire  valid_11_60; // @[Switch.scala 30:36:@3733.4]
  wire  _T_22072; // @[Switch.scala 30:53:@3735.4]
  wire  valid_11_61; // @[Switch.scala 30:36:@3736.4]
  wire  _T_22075; // @[Switch.scala 30:53:@3738.4]
  wire  valid_11_62; // @[Switch.scala 30:36:@3739.4]
  wire  _T_22078; // @[Switch.scala 30:53:@3741.4]
  wire  valid_11_63; // @[Switch.scala 30:36:@3742.4]
  wire [5:0] _T_22144; // @[Mux.scala 31:69:@3744.4]
  wire [5:0] _T_22145; // @[Mux.scala 31:69:@3745.4]
  wire [5:0] _T_22146; // @[Mux.scala 31:69:@3746.4]
  wire [5:0] _T_22147; // @[Mux.scala 31:69:@3747.4]
  wire [5:0] _T_22148; // @[Mux.scala 31:69:@3748.4]
  wire [5:0] _T_22149; // @[Mux.scala 31:69:@3749.4]
  wire [5:0] _T_22150; // @[Mux.scala 31:69:@3750.4]
  wire [5:0] _T_22151; // @[Mux.scala 31:69:@3751.4]
  wire [5:0] _T_22152; // @[Mux.scala 31:69:@3752.4]
  wire [5:0] _T_22153; // @[Mux.scala 31:69:@3753.4]
  wire [5:0] _T_22154; // @[Mux.scala 31:69:@3754.4]
  wire [5:0] _T_22155; // @[Mux.scala 31:69:@3755.4]
  wire [5:0] _T_22156; // @[Mux.scala 31:69:@3756.4]
  wire [5:0] _T_22157; // @[Mux.scala 31:69:@3757.4]
  wire [5:0] _T_22158; // @[Mux.scala 31:69:@3758.4]
  wire [5:0] _T_22159; // @[Mux.scala 31:69:@3759.4]
  wire [5:0] _T_22160; // @[Mux.scala 31:69:@3760.4]
  wire [5:0] _T_22161; // @[Mux.scala 31:69:@3761.4]
  wire [5:0] _T_22162; // @[Mux.scala 31:69:@3762.4]
  wire [5:0] _T_22163; // @[Mux.scala 31:69:@3763.4]
  wire [5:0] _T_22164; // @[Mux.scala 31:69:@3764.4]
  wire [5:0] _T_22165; // @[Mux.scala 31:69:@3765.4]
  wire [5:0] _T_22166; // @[Mux.scala 31:69:@3766.4]
  wire [5:0] _T_22167; // @[Mux.scala 31:69:@3767.4]
  wire [5:0] _T_22168; // @[Mux.scala 31:69:@3768.4]
  wire [5:0] _T_22169; // @[Mux.scala 31:69:@3769.4]
  wire [5:0] _T_22170; // @[Mux.scala 31:69:@3770.4]
  wire [5:0] _T_22171; // @[Mux.scala 31:69:@3771.4]
  wire [5:0] _T_22172; // @[Mux.scala 31:69:@3772.4]
  wire [5:0] _T_22173; // @[Mux.scala 31:69:@3773.4]
  wire [5:0] _T_22174; // @[Mux.scala 31:69:@3774.4]
  wire [5:0] _T_22175; // @[Mux.scala 31:69:@3775.4]
  wire [5:0] _T_22176; // @[Mux.scala 31:69:@3776.4]
  wire [5:0] _T_22177; // @[Mux.scala 31:69:@3777.4]
  wire [5:0] _T_22178; // @[Mux.scala 31:69:@3778.4]
  wire [5:0] _T_22179; // @[Mux.scala 31:69:@3779.4]
  wire [5:0] _T_22180; // @[Mux.scala 31:69:@3780.4]
  wire [5:0] _T_22181; // @[Mux.scala 31:69:@3781.4]
  wire [5:0] _T_22182; // @[Mux.scala 31:69:@3782.4]
  wire [5:0] _T_22183; // @[Mux.scala 31:69:@3783.4]
  wire [5:0] _T_22184; // @[Mux.scala 31:69:@3784.4]
  wire [5:0] _T_22185; // @[Mux.scala 31:69:@3785.4]
  wire [5:0] _T_22186; // @[Mux.scala 31:69:@3786.4]
  wire [5:0] _T_22187; // @[Mux.scala 31:69:@3787.4]
  wire [5:0] _T_22188; // @[Mux.scala 31:69:@3788.4]
  wire [5:0] _T_22189; // @[Mux.scala 31:69:@3789.4]
  wire [5:0] _T_22190; // @[Mux.scala 31:69:@3790.4]
  wire [5:0] _T_22191; // @[Mux.scala 31:69:@3791.4]
  wire [5:0] _T_22192; // @[Mux.scala 31:69:@3792.4]
  wire [5:0] _T_22193; // @[Mux.scala 31:69:@3793.4]
  wire [5:0] _T_22194; // @[Mux.scala 31:69:@3794.4]
  wire [5:0] _T_22195; // @[Mux.scala 31:69:@3795.4]
  wire [5:0] _T_22196; // @[Mux.scala 31:69:@3796.4]
  wire [5:0] _T_22197; // @[Mux.scala 31:69:@3797.4]
  wire [5:0] _T_22198; // @[Mux.scala 31:69:@3798.4]
  wire [5:0] _T_22199; // @[Mux.scala 31:69:@3799.4]
  wire [5:0] _T_22200; // @[Mux.scala 31:69:@3800.4]
  wire [5:0] _T_22201; // @[Mux.scala 31:69:@3801.4]
  wire [5:0] _T_22202; // @[Mux.scala 31:69:@3802.4]
  wire [5:0] _T_22203; // @[Mux.scala 31:69:@3803.4]
  wire [5:0] _T_22204; // @[Mux.scala 31:69:@3804.4]
  wire [5:0] _T_22205; // @[Mux.scala 31:69:@3805.4]
  wire [5:0] select_11; // @[Mux.scala 31:69:@3806.4]
  wire [47:0] _GEN_705; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_706; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_707; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_708; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_709; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_710; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_711; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_712; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_713; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_714; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_715; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_716; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_717; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_718; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_719; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_720; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_721; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_722; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_723; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_724; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_725; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_726; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_727; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_728; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_729; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_730; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_731; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_732; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_733; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_734; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_735; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_736; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_737; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_738; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_739; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_740; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_741; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_742; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_743; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_744; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_745; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_746; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_747; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_748; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_749; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_750; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_751; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_752; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_753; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_754; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_755; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_756; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_757; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_758; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_759; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_760; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_761; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_762; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_763; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_764; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_765; // @[Switch.scala 33:19:@3808.4]
  wire [47:0] _GEN_766; // @[Switch.scala 33:19:@3808.4]
  wire [7:0] _T_22214; // @[Switch.scala 34:32:@3815.4]
  wire [15:0] _T_22222; // @[Switch.scala 34:32:@3823.4]
  wire [7:0] _T_22229; // @[Switch.scala 34:32:@3830.4]
  wire [31:0] _T_22238; // @[Switch.scala 34:32:@3839.4]
  wire [7:0] _T_22245; // @[Switch.scala 34:32:@3846.4]
  wire [15:0] _T_22253; // @[Switch.scala 34:32:@3854.4]
  wire [7:0] _T_22260; // @[Switch.scala 34:32:@3861.4]
  wire [31:0] _T_22269; // @[Switch.scala 34:32:@3870.4]
  wire [63:0] _T_22270; // @[Switch.scala 34:32:@3871.4]
  wire  _T_22274; // @[Switch.scala 30:53:@3874.4]
  wire  valid_12_0; // @[Switch.scala 30:36:@3875.4]
  wire  _T_22277; // @[Switch.scala 30:53:@3877.4]
  wire  valid_12_1; // @[Switch.scala 30:36:@3878.4]
  wire  _T_22280; // @[Switch.scala 30:53:@3880.4]
  wire  valid_12_2; // @[Switch.scala 30:36:@3881.4]
  wire  _T_22283; // @[Switch.scala 30:53:@3883.4]
  wire  valid_12_3; // @[Switch.scala 30:36:@3884.4]
  wire  _T_22286; // @[Switch.scala 30:53:@3886.4]
  wire  valid_12_4; // @[Switch.scala 30:36:@3887.4]
  wire  _T_22289; // @[Switch.scala 30:53:@3889.4]
  wire  valid_12_5; // @[Switch.scala 30:36:@3890.4]
  wire  _T_22292; // @[Switch.scala 30:53:@3892.4]
  wire  valid_12_6; // @[Switch.scala 30:36:@3893.4]
  wire  _T_22295; // @[Switch.scala 30:53:@3895.4]
  wire  valid_12_7; // @[Switch.scala 30:36:@3896.4]
  wire  _T_22298; // @[Switch.scala 30:53:@3898.4]
  wire  valid_12_8; // @[Switch.scala 30:36:@3899.4]
  wire  _T_22301; // @[Switch.scala 30:53:@3901.4]
  wire  valid_12_9; // @[Switch.scala 30:36:@3902.4]
  wire  _T_22304; // @[Switch.scala 30:53:@3904.4]
  wire  valid_12_10; // @[Switch.scala 30:36:@3905.4]
  wire  _T_22307; // @[Switch.scala 30:53:@3907.4]
  wire  valid_12_11; // @[Switch.scala 30:36:@3908.4]
  wire  _T_22310; // @[Switch.scala 30:53:@3910.4]
  wire  valid_12_12; // @[Switch.scala 30:36:@3911.4]
  wire  _T_22313; // @[Switch.scala 30:53:@3913.4]
  wire  valid_12_13; // @[Switch.scala 30:36:@3914.4]
  wire  _T_22316; // @[Switch.scala 30:53:@3916.4]
  wire  valid_12_14; // @[Switch.scala 30:36:@3917.4]
  wire  _T_22319; // @[Switch.scala 30:53:@3919.4]
  wire  valid_12_15; // @[Switch.scala 30:36:@3920.4]
  wire  _T_22322; // @[Switch.scala 30:53:@3922.4]
  wire  valid_12_16; // @[Switch.scala 30:36:@3923.4]
  wire  _T_22325; // @[Switch.scala 30:53:@3925.4]
  wire  valid_12_17; // @[Switch.scala 30:36:@3926.4]
  wire  _T_22328; // @[Switch.scala 30:53:@3928.4]
  wire  valid_12_18; // @[Switch.scala 30:36:@3929.4]
  wire  _T_22331; // @[Switch.scala 30:53:@3931.4]
  wire  valid_12_19; // @[Switch.scala 30:36:@3932.4]
  wire  _T_22334; // @[Switch.scala 30:53:@3934.4]
  wire  valid_12_20; // @[Switch.scala 30:36:@3935.4]
  wire  _T_22337; // @[Switch.scala 30:53:@3937.4]
  wire  valid_12_21; // @[Switch.scala 30:36:@3938.4]
  wire  _T_22340; // @[Switch.scala 30:53:@3940.4]
  wire  valid_12_22; // @[Switch.scala 30:36:@3941.4]
  wire  _T_22343; // @[Switch.scala 30:53:@3943.4]
  wire  valid_12_23; // @[Switch.scala 30:36:@3944.4]
  wire  _T_22346; // @[Switch.scala 30:53:@3946.4]
  wire  valid_12_24; // @[Switch.scala 30:36:@3947.4]
  wire  _T_22349; // @[Switch.scala 30:53:@3949.4]
  wire  valid_12_25; // @[Switch.scala 30:36:@3950.4]
  wire  _T_22352; // @[Switch.scala 30:53:@3952.4]
  wire  valid_12_26; // @[Switch.scala 30:36:@3953.4]
  wire  _T_22355; // @[Switch.scala 30:53:@3955.4]
  wire  valid_12_27; // @[Switch.scala 30:36:@3956.4]
  wire  _T_22358; // @[Switch.scala 30:53:@3958.4]
  wire  valid_12_28; // @[Switch.scala 30:36:@3959.4]
  wire  _T_22361; // @[Switch.scala 30:53:@3961.4]
  wire  valid_12_29; // @[Switch.scala 30:36:@3962.4]
  wire  _T_22364; // @[Switch.scala 30:53:@3964.4]
  wire  valid_12_30; // @[Switch.scala 30:36:@3965.4]
  wire  _T_22367; // @[Switch.scala 30:53:@3967.4]
  wire  valid_12_31; // @[Switch.scala 30:36:@3968.4]
  wire  _T_22370; // @[Switch.scala 30:53:@3970.4]
  wire  valid_12_32; // @[Switch.scala 30:36:@3971.4]
  wire  _T_22373; // @[Switch.scala 30:53:@3973.4]
  wire  valid_12_33; // @[Switch.scala 30:36:@3974.4]
  wire  _T_22376; // @[Switch.scala 30:53:@3976.4]
  wire  valid_12_34; // @[Switch.scala 30:36:@3977.4]
  wire  _T_22379; // @[Switch.scala 30:53:@3979.4]
  wire  valid_12_35; // @[Switch.scala 30:36:@3980.4]
  wire  _T_22382; // @[Switch.scala 30:53:@3982.4]
  wire  valid_12_36; // @[Switch.scala 30:36:@3983.4]
  wire  _T_22385; // @[Switch.scala 30:53:@3985.4]
  wire  valid_12_37; // @[Switch.scala 30:36:@3986.4]
  wire  _T_22388; // @[Switch.scala 30:53:@3988.4]
  wire  valid_12_38; // @[Switch.scala 30:36:@3989.4]
  wire  _T_22391; // @[Switch.scala 30:53:@3991.4]
  wire  valid_12_39; // @[Switch.scala 30:36:@3992.4]
  wire  _T_22394; // @[Switch.scala 30:53:@3994.4]
  wire  valid_12_40; // @[Switch.scala 30:36:@3995.4]
  wire  _T_22397; // @[Switch.scala 30:53:@3997.4]
  wire  valid_12_41; // @[Switch.scala 30:36:@3998.4]
  wire  _T_22400; // @[Switch.scala 30:53:@4000.4]
  wire  valid_12_42; // @[Switch.scala 30:36:@4001.4]
  wire  _T_22403; // @[Switch.scala 30:53:@4003.4]
  wire  valid_12_43; // @[Switch.scala 30:36:@4004.4]
  wire  _T_22406; // @[Switch.scala 30:53:@4006.4]
  wire  valid_12_44; // @[Switch.scala 30:36:@4007.4]
  wire  _T_22409; // @[Switch.scala 30:53:@4009.4]
  wire  valid_12_45; // @[Switch.scala 30:36:@4010.4]
  wire  _T_22412; // @[Switch.scala 30:53:@4012.4]
  wire  valid_12_46; // @[Switch.scala 30:36:@4013.4]
  wire  _T_22415; // @[Switch.scala 30:53:@4015.4]
  wire  valid_12_47; // @[Switch.scala 30:36:@4016.4]
  wire  _T_22418; // @[Switch.scala 30:53:@4018.4]
  wire  valid_12_48; // @[Switch.scala 30:36:@4019.4]
  wire  _T_22421; // @[Switch.scala 30:53:@4021.4]
  wire  valid_12_49; // @[Switch.scala 30:36:@4022.4]
  wire  _T_22424; // @[Switch.scala 30:53:@4024.4]
  wire  valid_12_50; // @[Switch.scala 30:36:@4025.4]
  wire  _T_22427; // @[Switch.scala 30:53:@4027.4]
  wire  valid_12_51; // @[Switch.scala 30:36:@4028.4]
  wire  _T_22430; // @[Switch.scala 30:53:@4030.4]
  wire  valid_12_52; // @[Switch.scala 30:36:@4031.4]
  wire  _T_22433; // @[Switch.scala 30:53:@4033.4]
  wire  valid_12_53; // @[Switch.scala 30:36:@4034.4]
  wire  _T_22436; // @[Switch.scala 30:53:@4036.4]
  wire  valid_12_54; // @[Switch.scala 30:36:@4037.4]
  wire  _T_22439; // @[Switch.scala 30:53:@4039.4]
  wire  valid_12_55; // @[Switch.scala 30:36:@4040.4]
  wire  _T_22442; // @[Switch.scala 30:53:@4042.4]
  wire  valid_12_56; // @[Switch.scala 30:36:@4043.4]
  wire  _T_22445; // @[Switch.scala 30:53:@4045.4]
  wire  valid_12_57; // @[Switch.scala 30:36:@4046.4]
  wire  _T_22448; // @[Switch.scala 30:53:@4048.4]
  wire  valid_12_58; // @[Switch.scala 30:36:@4049.4]
  wire  _T_22451; // @[Switch.scala 30:53:@4051.4]
  wire  valid_12_59; // @[Switch.scala 30:36:@4052.4]
  wire  _T_22454; // @[Switch.scala 30:53:@4054.4]
  wire  valid_12_60; // @[Switch.scala 30:36:@4055.4]
  wire  _T_22457; // @[Switch.scala 30:53:@4057.4]
  wire  valid_12_61; // @[Switch.scala 30:36:@4058.4]
  wire  _T_22460; // @[Switch.scala 30:53:@4060.4]
  wire  valid_12_62; // @[Switch.scala 30:36:@4061.4]
  wire  _T_22463; // @[Switch.scala 30:53:@4063.4]
  wire  valid_12_63; // @[Switch.scala 30:36:@4064.4]
  wire [5:0] _T_22529; // @[Mux.scala 31:69:@4066.4]
  wire [5:0] _T_22530; // @[Mux.scala 31:69:@4067.4]
  wire [5:0] _T_22531; // @[Mux.scala 31:69:@4068.4]
  wire [5:0] _T_22532; // @[Mux.scala 31:69:@4069.4]
  wire [5:0] _T_22533; // @[Mux.scala 31:69:@4070.4]
  wire [5:0] _T_22534; // @[Mux.scala 31:69:@4071.4]
  wire [5:0] _T_22535; // @[Mux.scala 31:69:@4072.4]
  wire [5:0] _T_22536; // @[Mux.scala 31:69:@4073.4]
  wire [5:0] _T_22537; // @[Mux.scala 31:69:@4074.4]
  wire [5:0] _T_22538; // @[Mux.scala 31:69:@4075.4]
  wire [5:0] _T_22539; // @[Mux.scala 31:69:@4076.4]
  wire [5:0] _T_22540; // @[Mux.scala 31:69:@4077.4]
  wire [5:0] _T_22541; // @[Mux.scala 31:69:@4078.4]
  wire [5:0] _T_22542; // @[Mux.scala 31:69:@4079.4]
  wire [5:0] _T_22543; // @[Mux.scala 31:69:@4080.4]
  wire [5:0] _T_22544; // @[Mux.scala 31:69:@4081.4]
  wire [5:0] _T_22545; // @[Mux.scala 31:69:@4082.4]
  wire [5:0] _T_22546; // @[Mux.scala 31:69:@4083.4]
  wire [5:0] _T_22547; // @[Mux.scala 31:69:@4084.4]
  wire [5:0] _T_22548; // @[Mux.scala 31:69:@4085.4]
  wire [5:0] _T_22549; // @[Mux.scala 31:69:@4086.4]
  wire [5:0] _T_22550; // @[Mux.scala 31:69:@4087.4]
  wire [5:0] _T_22551; // @[Mux.scala 31:69:@4088.4]
  wire [5:0] _T_22552; // @[Mux.scala 31:69:@4089.4]
  wire [5:0] _T_22553; // @[Mux.scala 31:69:@4090.4]
  wire [5:0] _T_22554; // @[Mux.scala 31:69:@4091.4]
  wire [5:0] _T_22555; // @[Mux.scala 31:69:@4092.4]
  wire [5:0] _T_22556; // @[Mux.scala 31:69:@4093.4]
  wire [5:0] _T_22557; // @[Mux.scala 31:69:@4094.4]
  wire [5:0] _T_22558; // @[Mux.scala 31:69:@4095.4]
  wire [5:0] _T_22559; // @[Mux.scala 31:69:@4096.4]
  wire [5:0] _T_22560; // @[Mux.scala 31:69:@4097.4]
  wire [5:0] _T_22561; // @[Mux.scala 31:69:@4098.4]
  wire [5:0] _T_22562; // @[Mux.scala 31:69:@4099.4]
  wire [5:0] _T_22563; // @[Mux.scala 31:69:@4100.4]
  wire [5:0] _T_22564; // @[Mux.scala 31:69:@4101.4]
  wire [5:0] _T_22565; // @[Mux.scala 31:69:@4102.4]
  wire [5:0] _T_22566; // @[Mux.scala 31:69:@4103.4]
  wire [5:0] _T_22567; // @[Mux.scala 31:69:@4104.4]
  wire [5:0] _T_22568; // @[Mux.scala 31:69:@4105.4]
  wire [5:0] _T_22569; // @[Mux.scala 31:69:@4106.4]
  wire [5:0] _T_22570; // @[Mux.scala 31:69:@4107.4]
  wire [5:0] _T_22571; // @[Mux.scala 31:69:@4108.4]
  wire [5:0] _T_22572; // @[Mux.scala 31:69:@4109.4]
  wire [5:0] _T_22573; // @[Mux.scala 31:69:@4110.4]
  wire [5:0] _T_22574; // @[Mux.scala 31:69:@4111.4]
  wire [5:0] _T_22575; // @[Mux.scala 31:69:@4112.4]
  wire [5:0] _T_22576; // @[Mux.scala 31:69:@4113.4]
  wire [5:0] _T_22577; // @[Mux.scala 31:69:@4114.4]
  wire [5:0] _T_22578; // @[Mux.scala 31:69:@4115.4]
  wire [5:0] _T_22579; // @[Mux.scala 31:69:@4116.4]
  wire [5:0] _T_22580; // @[Mux.scala 31:69:@4117.4]
  wire [5:0] _T_22581; // @[Mux.scala 31:69:@4118.4]
  wire [5:0] _T_22582; // @[Mux.scala 31:69:@4119.4]
  wire [5:0] _T_22583; // @[Mux.scala 31:69:@4120.4]
  wire [5:0] _T_22584; // @[Mux.scala 31:69:@4121.4]
  wire [5:0] _T_22585; // @[Mux.scala 31:69:@4122.4]
  wire [5:0] _T_22586; // @[Mux.scala 31:69:@4123.4]
  wire [5:0] _T_22587; // @[Mux.scala 31:69:@4124.4]
  wire [5:0] _T_22588; // @[Mux.scala 31:69:@4125.4]
  wire [5:0] _T_22589; // @[Mux.scala 31:69:@4126.4]
  wire [5:0] _T_22590; // @[Mux.scala 31:69:@4127.4]
  wire [5:0] select_12; // @[Mux.scala 31:69:@4128.4]
  wire [47:0] _GEN_769; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_770; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_771; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_772; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_773; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_774; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_775; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_776; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_777; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_778; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_779; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_780; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_781; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_782; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_783; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_784; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_785; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_786; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_787; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_788; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_789; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_790; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_791; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_792; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_793; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_794; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_795; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_796; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_797; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_798; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_799; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_800; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_801; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_802; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_803; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_804; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_805; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_806; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_807; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_808; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_809; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_810; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_811; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_812; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_813; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_814; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_815; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_816; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_817; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_818; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_819; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_820; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_821; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_822; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_823; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_824; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_825; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_826; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_827; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_828; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_829; // @[Switch.scala 33:19:@4130.4]
  wire [47:0] _GEN_830; // @[Switch.scala 33:19:@4130.4]
  wire [7:0] _T_22599; // @[Switch.scala 34:32:@4137.4]
  wire [15:0] _T_22607; // @[Switch.scala 34:32:@4145.4]
  wire [7:0] _T_22614; // @[Switch.scala 34:32:@4152.4]
  wire [31:0] _T_22623; // @[Switch.scala 34:32:@4161.4]
  wire [7:0] _T_22630; // @[Switch.scala 34:32:@4168.4]
  wire [15:0] _T_22638; // @[Switch.scala 34:32:@4176.4]
  wire [7:0] _T_22645; // @[Switch.scala 34:32:@4183.4]
  wire [31:0] _T_22654; // @[Switch.scala 34:32:@4192.4]
  wire [63:0] _T_22655; // @[Switch.scala 34:32:@4193.4]
  wire  _T_22659; // @[Switch.scala 30:53:@4196.4]
  wire  valid_13_0; // @[Switch.scala 30:36:@4197.4]
  wire  _T_22662; // @[Switch.scala 30:53:@4199.4]
  wire  valid_13_1; // @[Switch.scala 30:36:@4200.4]
  wire  _T_22665; // @[Switch.scala 30:53:@4202.4]
  wire  valid_13_2; // @[Switch.scala 30:36:@4203.4]
  wire  _T_22668; // @[Switch.scala 30:53:@4205.4]
  wire  valid_13_3; // @[Switch.scala 30:36:@4206.4]
  wire  _T_22671; // @[Switch.scala 30:53:@4208.4]
  wire  valid_13_4; // @[Switch.scala 30:36:@4209.4]
  wire  _T_22674; // @[Switch.scala 30:53:@4211.4]
  wire  valid_13_5; // @[Switch.scala 30:36:@4212.4]
  wire  _T_22677; // @[Switch.scala 30:53:@4214.4]
  wire  valid_13_6; // @[Switch.scala 30:36:@4215.4]
  wire  _T_22680; // @[Switch.scala 30:53:@4217.4]
  wire  valid_13_7; // @[Switch.scala 30:36:@4218.4]
  wire  _T_22683; // @[Switch.scala 30:53:@4220.4]
  wire  valid_13_8; // @[Switch.scala 30:36:@4221.4]
  wire  _T_22686; // @[Switch.scala 30:53:@4223.4]
  wire  valid_13_9; // @[Switch.scala 30:36:@4224.4]
  wire  _T_22689; // @[Switch.scala 30:53:@4226.4]
  wire  valid_13_10; // @[Switch.scala 30:36:@4227.4]
  wire  _T_22692; // @[Switch.scala 30:53:@4229.4]
  wire  valid_13_11; // @[Switch.scala 30:36:@4230.4]
  wire  _T_22695; // @[Switch.scala 30:53:@4232.4]
  wire  valid_13_12; // @[Switch.scala 30:36:@4233.4]
  wire  _T_22698; // @[Switch.scala 30:53:@4235.4]
  wire  valid_13_13; // @[Switch.scala 30:36:@4236.4]
  wire  _T_22701; // @[Switch.scala 30:53:@4238.4]
  wire  valid_13_14; // @[Switch.scala 30:36:@4239.4]
  wire  _T_22704; // @[Switch.scala 30:53:@4241.4]
  wire  valid_13_15; // @[Switch.scala 30:36:@4242.4]
  wire  _T_22707; // @[Switch.scala 30:53:@4244.4]
  wire  valid_13_16; // @[Switch.scala 30:36:@4245.4]
  wire  _T_22710; // @[Switch.scala 30:53:@4247.4]
  wire  valid_13_17; // @[Switch.scala 30:36:@4248.4]
  wire  _T_22713; // @[Switch.scala 30:53:@4250.4]
  wire  valid_13_18; // @[Switch.scala 30:36:@4251.4]
  wire  _T_22716; // @[Switch.scala 30:53:@4253.4]
  wire  valid_13_19; // @[Switch.scala 30:36:@4254.4]
  wire  _T_22719; // @[Switch.scala 30:53:@4256.4]
  wire  valid_13_20; // @[Switch.scala 30:36:@4257.4]
  wire  _T_22722; // @[Switch.scala 30:53:@4259.4]
  wire  valid_13_21; // @[Switch.scala 30:36:@4260.4]
  wire  _T_22725; // @[Switch.scala 30:53:@4262.4]
  wire  valid_13_22; // @[Switch.scala 30:36:@4263.4]
  wire  _T_22728; // @[Switch.scala 30:53:@4265.4]
  wire  valid_13_23; // @[Switch.scala 30:36:@4266.4]
  wire  _T_22731; // @[Switch.scala 30:53:@4268.4]
  wire  valid_13_24; // @[Switch.scala 30:36:@4269.4]
  wire  _T_22734; // @[Switch.scala 30:53:@4271.4]
  wire  valid_13_25; // @[Switch.scala 30:36:@4272.4]
  wire  _T_22737; // @[Switch.scala 30:53:@4274.4]
  wire  valid_13_26; // @[Switch.scala 30:36:@4275.4]
  wire  _T_22740; // @[Switch.scala 30:53:@4277.4]
  wire  valid_13_27; // @[Switch.scala 30:36:@4278.4]
  wire  _T_22743; // @[Switch.scala 30:53:@4280.4]
  wire  valid_13_28; // @[Switch.scala 30:36:@4281.4]
  wire  _T_22746; // @[Switch.scala 30:53:@4283.4]
  wire  valid_13_29; // @[Switch.scala 30:36:@4284.4]
  wire  _T_22749; // @[Switch.scala 30:53:@4286.4]
  wire  valid_13_30; // @[Switch.scala 30:36:@4287.4]
  wire  _T_22752; // @[Switch.scala 30:53:@4289.4]
  wire  valid_13_31; // @[Switch.scala 30:36:@4290.4]
  wire  _T_22755; // @[Switch.scala 30:53:@4292.4]
  wire  valid_13_32; // @[Switch.scala 30:36:@4293.4]
  wire  _T_22758; // @[Switch.scala 30:53:@4295.4]
  wire  valid_13_33; // @[Switch.scala 30:36:@4296.4]
  wire  _T_22761; // @[Switch.scala 30:53:@4298.4]
  wire  valid_13_34; // @[Switch.scala 30:36:@4299.4]
  wire  _T_22764; // @[Switch.scala 30:53:@4301.4]
  wire  valid_13_35; // @[Switch.scala 30:36:@4302.4]
  wire  _T_22767; // @[Switch.scala 30:53:@4304.4]
  wire  valid_13_36; // @[Switch.scala 30:36:@4305.4]
  wire  _T_22770; // @[Switch.scala 30:53:@4307.4]
  wire  valid_13_37; // @[Switch.scala 30:36:@4308.4]
  wire  _T_22773; // @[Switch.scala 30:53:@4310.4]
  wire  valid_13_38; // @[Switch.scala 30:36:@4311.4]
  wire  _T_22776; // @[Switch.scala 30:53:@4313.4]
  wire  valid_13_39; // @[Switch.scala 30:36:@4314.4]
  wire  _T_22779; // @[Switch.scala 30:53:@4316.4]
  wire  valid_13_40; // @[Switch.scala 30:36:@4317.4]
  wire  _T_22782; // @[Switch.scala 30:53:@4319.4]
  wire  valid_13_41; // @[Switch.scala 30:36:@4320.4]
  wire  _T_22785; // @[Switch.scala 30:53:@4322.4]
  wire  valid_13_42; // @[Switch.scala 30:36:@4323.4]
  wire  _T_22788; // @[Switch.scala 30:53:@4325.4]
  wire  valid_13_43; // @[Switch.scala 30:36:@4326.4]
  wire  _T_22791; // @[Switch.scala 30:53:@4328.4]
  wire  valid_13_44; // @[Switch.scala 30:36:@4329.4]
  wire  _T_22794; // @[Switch.scala 30:53:@4331.4]
  wire  valid_13_45; // @[Switch.scala 30:36:@4332.4]
  wire  _T_22797; // @[Switch.scala 30:53:@4334.4]
  wire  valid_13_46; // @[Switch.scala 30:36:@4335.4]
  wire  _T_22800; // @[Switch.scala 30:53:@4337.4]
  wire  valid_13_47; // @[Switch.scala 30:36:@4338.4]
  wire  _T_22803; // @[Switch.scala 30:53:@4340.4]
  wire  valid_13_48; // @[Switch.scala 30:36:@4341.4]
  wire  _T_22806; // @[Switch.scala 30:53:@4343.4]
  wire  valid_13_49; // @[Switch.scala 30:36:@4344.4]
  wire  _T_22809; // @[Switch.scala 30:53:@4346.4]
  wire  valid_13_50; // @[Switch.scala 30:36:@4347.4]
  wire  _T_22812; // @[Switch.scala 30:53:@4349.4]
  wire  valid_13_51; // @[Switch.scala 30:36:@4350.4]
  wire  _T_22815; // @[Switch.scala 30:53:@4352.4]
  wire  valid_13_52; // @[Switch.scala 30:36:@4353.4]
  wire  _T_22818; // @[Switch.scala 30:53:@4355.4]
  wire  valid_13_53; // @[Switch.scala 30:36:@4356.4]
  wire  _T_22821; // @[Switch.scala 30:53:@4358.4]
  wire  valid_13_54; // @[Switch.scala 30:36:@4359.4]
  wire  _T_22824; // @[Switch.scala 30:53:@4361.4]
  wire  valid_13_55; // @[Switch.scala 30:36:@4362.4]
  wire  _T_22827; // @[Switch.scala 30:53:@4364.4]
  wire  valid_13_56; // @[Switch.scala 30:36:@4365.4]
  wire  _T_22830; // @[Switch.scala 30:53:@4367.4]
  wire  valid_13_57; // @[Switch.scala 30:36:@4368.4]
  wire  _T_22833; // @[Switch.scala 30:53:@4370.4]
  wire  valid_13_58; // @[Switch.scala 30:36:@4371.4]
  wire  _T_22836; // @[Switch.scala 30:53:@4373.4]
  wire  valid_13_59; // @[Switch.scala 30:36:@4374.4]
  wire  _T_22839; // @[Switch.scala 30:53:@4376.4]
  wire  valid_13_60; // @[Switch.scala 30:36:@4377.4]
  wire  _T_22842; // @[Switch.scala 30:53:@4379.4]
  wire  valid_13_61; // @[Switch.scala 30:36:@4380.4]
  wire  _T_22845; // @[Switch.scala 30:53:@4382.4]
  wire  valid_13_62; // @[Switch.scala 30:36:@4383.4]
  wire  _T_22848; // @[Switch.scala 30:53:@4385.4]
  wire  valid_13_63; // @[Switch.scala 30:36:@4386.4]
  wire [5:0] _T_22914; // @[Mux.scala 31:69:@4388.4]
  wire [5:0] _T_22915; // @[Mux.scala 31:69:@4389.4]
  wire [5:0] _T_22916; // @[Mux.scala 31:69:@4390.4]
  wire [5:0] _T_22917; // @[Mux.scala 31:69:@4391.4]
  wire [5:0] _T_22918; // @[Mux.scala 31:69:@4392.4]
  wire [5:0] _T_22919; // @[Mux.scala 31:69:@4393.4]
  wire [5:0] _T_22920; // @[Mux.scala 31:69:@4394.4]
  wire [5:0] _T_22921; // @[Mux.scala 31:69:@4395.4]
  wire [5:0] _T_22922; // @[Mux.scala 31:69:@4396.4]
  wire [5:0] _T_22923; // @[Mux.scala 31:69:@4397.4]
  wire [5:0] _T_22924; // @[Mux.scala 31:69:@4398.4]
  wire [5:0] _T_22925; // @[Mux.scala 31:69:@4399.4]
  wire [5:0] _T_22926; // @[Mux.scala 31:69:@4400.4]
  wire [5:0] _T_22927; // @[Mux.scala 31:69:@4401.4]
  wire [5:0] _T_22928; // @[Mux.scala 31:69:@4402.4]
  wire [5:0] _T_22929; // @[Mux.scala 31:69:@4403.4]
  wire [5:0] _T_22930; // @[Mux.scala 31:69:@4404.4]
  wire [5:0] _T_22931; // @[Mux.scala 31:69:@4405.4]
  wire [5:0] _T_22932; // @[Mux.scala 31:69:@4406.4]
  wire [5:0] _T_22933; // @[Mux.scala 31:69:@4407.4]
  wire [5:0] _T_22934; // @[Mux.scala 31:69:@4408.4]
  wire [5:0] _T_22935; // @[Mux.scala 31:69:@4409.4]
  wire [5:0] _T_22936; // @[Mux.scala 31:69:@4410.4]
  wire [5:0] _T_22937; // @[Mux.scala 31:69:@4411.4]
  wire [5:0] _T_22938; // @[Mux.scala 31:69:@4412.4]
  wire [5:0] _T_22939; // @[Mux.scala 31:69:@4413.4]
  wire [5:0] _T_22940; // @[Mux.scala 31:69:@4414.4]
  wire [5:0] _T_22941; // @[Mux.scala 31:69:@4415.4]
  wire [5:0] _T_22942; // @[Mux.scala 31:69:@4416.4]
  wire [5:0] _T_22943; // @[Mux.scala 31:69:@4417.4]
  wire [5:0] _T_22944; // @[Mux.scala 31:69:@4418.4]
  wire [5:0] _T_22945; // @[Mux.scala 31:69:@4419.4]
  wire [5:0] _T_22946; // @[Mux.scala 31:69:@4420.4]
  wire [5:0] _T_22947; // @[Mux.scala 31:69:@4421.4]
  wire [5:0] _T_22948; // @[Mux.scala 31:69:@4422.4]
  wire [5:0] _T_22949; // @[Mux.scala 31:69:@4423.4]
  wire [5:0] _T_22950; // @[Mux.scala 31:69:@4424.4]
  wire [5:0] _T_22951; // @[Mux.scala 31:69:@4425.4]
  wire [5:0] _T_22952; // @[Mux.scala 31:69:@4426.4]
  wire [5:0] _T_22953; // @[Mux.scala 31:69:@4427.4]
  wire [5:0] _T_22954; // @[Mux.scala 31:69:@4428.4]
  wire [5:0] _T_22955; // @[Mux.scala 31:69:@4429.4]
  wire [5:0] _T_22956; // @[Mux.scala 31:69:@4430.4]
  wire [5:0] _T_22957; // @[Mux.scala 31:69:@4431.4]
  wire [5:0] _T_22958; // @[Mux.scala 31:69:@4432.4]
  wire [5:0] _T_22959; // @[Mux.scala 31:69:@4433.4]
  wire [5:0] _T_22960; // @[Mux.scala 31:69:@4434.4]
  wire [5:0] _T_22961; // @[Mux.scala 31:69:@4435.4]
  wire [5:0] _T_22962; // @[Mux.scala 31:69:@4436.4]
  wire [5:0] _T_22963; // @[Mux.scala 31:69:@4437.4]
  wire [5:0] _T_22964; // @[Mux.scala 31:69:@4438.4]
  wire [5:0] _T_22965; // @[Mux.scala 31:69:@4439.4]
  wire [5:0] _T_22966; // @[Mux.scala 31:69:@4440.4]
  wire [5:0] _T_22967; // @[Mux.scala 31:69:@4441.4]
  wire [5:0] _T_22968; // @[Mux.scala 31:69:@4442.4]
  wire [5:0] _T_22969; // @[Mux.scala 31:69:@4443.4]
  wire [5:0] _T_22970; // @[Mux.scala 31:69:@4444.4]
  wire [5:0] _T_22971; // @[Mux.scala 31:69:@4445.4]
  wire [5:0] _T_22972; // @[Mux.scala 31:69:@4446.4]
  wire [5:0] _T_22973; // @[Mux.scala 31:69:@4447.4]
  wire [5:0] _T_22974; // @[Mux.scala 31:69:@4448.4]
  wire [5:0] _T_22975; // @[Mux.scala 31:69:@4449.4]
  wire [5:0] select_13; // @[Mux.scala 31:69:@4450.4]
  wire [47:0] _GEN_833; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_834; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_835; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_836; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_837; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_838; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_839; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_840; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_841; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_842; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_843; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_844; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_845; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_846; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_847; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_848; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_849; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_850; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_851; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_852; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_853; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_854; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_855; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_856; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_857; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_858; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_859; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_860; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_861; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_862; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_863; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_864; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_865; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_866; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_867; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_868; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_869; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_870; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_871; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_872; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_873; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_874; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_875; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_876; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_877; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_878; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_879; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_880; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_881; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_882; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_883; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_884; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_885; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_886; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_887; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_888; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_889; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_890; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_891; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_892; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_893; // @[Switch.scala 33:19:@4452.4]
  wire [47:0] _GEN_894; // @[Switch.scala 33:19:@4452.4]
  wire [7:0] _T_22984; // @[Switch.scala 34:32:@4459.4]
  wire [15:0] _T_22992; // @[Switch.scala 34:32:@4467.4]
  wire [7:0] _T_22999; // @[Switch.scala 34:32:@4474.4]
  wire [31:0] _T_23008; // @[Switch.scala 34:32:@4483.4]
  wire [7:0] _T_23015; // @[Switch.scala 34:32:@4490.4]
  wire [15:0] _T_23023; // @[Switch.scala 34:32:@4498.4]
  wire [7:0] _T_23030; // @[Switch.scala 34:32:@4505.4]
  wire [31:0] _T_23039; // @[Switch.scala 34:32:@4514.4]
  wire [63:0] _T_23040; // @[Switch.scala 34:32:@4515.4]
  wire  _T_23044; // @[Switch.scala 30:53:@4518.4]
  wire  valid_14_0; // @[Switch.scala 30:36:@4519.4]
  wire  _T_23047; // @[Switch.scala 30:53:@4521.4]
  wire  valid_14_1; // @[Switch.scala 30:36:@4522.4]
  wire  _T_23050; // @[Switch.scala 30:53:@4524.4]
  wire  valid_14_2; // @[Switch.scala 30:36:@4525.4]
  wire  _T_23053; // @[Switch.scala 30:53:@4527.4]
  wire  valid_14_3; // @[Switch.scala 30:36:@4528.4]
  wire  _T_23056; // @[Switch.scala 30:53:@4530.4]
  wire  valid_14_4; // @[Switch.scala 30:36:@4531.4]
  wire  _T_23059; // @[Switch.scala 30:53:@4533.4]
  wire  valid_14_5; // @[Switch.scala 30:36:@4534.4]
  wire  _T_23062; // @[Switch.scala 30:53:@4536.4]
  wire  valid_14_6; // @[Switch.scala 30:36:@4537.4]
  wire  _T_23065; // @[Switch.scala 30:53:@4539.4]
  wire  valid_14_7; // @[Switch.scala 30:36:@4540.4]
  wire  _T_23068; // @[Switch.scala 30:53:@4542.4]
  wire  valid_14_8; // @[Switch.scala 30:36:@4543.4]
  wire  _T_23071; // @[Switch.scala 30:53:@4545.4]
  wire  valid_14_9; // @[Switch.scala 30:36:@4546.4]
  wire  _T_23074; // @[Switch.scala 30:53:@4548.4]
  wire  valid_14_10; // @[Switch.scala 30:36:@4549.4]
  wire  _T_23077; // @[Switch.scala 30:53:@4551.4]
  wire  valid_14_11; // @[Switch.scala 30:36:@4552.4]
  wire  _T_23080; // @[Switch.scala 30:53:@4554.4]
  wire  valid_14_12; // @[Switch.scala 30:36:@4555.4]
  wire  _T_23083; // @[Switch.scala 30:53:@4557.4]
  wire  valid_14_13; // @[Switch.scala 30:36:@4558.4]
  wire  _T_23086; // @[Switch.scala 30:53:@4560.4]
  wire  valid_14_14; // @[Switch.scala 30:36:@4561.4]
  wire  _T_23089; // @[Switch.scala 30:53:@4563.4]
  wire  valid_14_15; // @[Switch.scala 30:36:@4564.4]
  wire  _T_23092; // @[Switch.scala 30:53:@4566.4]
  wire  valid_14_16; // @[Switch.scala 30:36:@4567.4]
  wire  _T_23095; // @[Switch.scala 30:53:@4569.4]
  wire  valid_14_17; // @[Switch.scala 30:36:@4570.4]
  wire  _T_23098; // @[Switch.scala 30:53:@4572.4]
  wire  valid_14_18; // @[Switch.scala 30:36:@4573.4]
  wire  _T_23101; // @[Switch.scala 30:53:@4575.4]
  wire  valid_14_19; // @[Switch.scala 30:36:@4576.4]
  wire  _T_23104; // @[Switch.scala 30:53:@4578.4]
  wire  valid_14_20; // @[Switch.scala 30:36:@4579.4]
  wire  _T_23107; // @[Switch.scala 30:53:@4581.4]
  wire  valid_14_21; // @[Switch.scala 30:36:@4582.4]
  wire  _T_23110; // @[Switch.scala 30:53:@4584.4]
  wire  valid_14_22; // @[Switch.scala 30:36:@4585.4]
  wire  _T_23113; // @[Switch.scala 30:53:@4587.4]
  wire  valid_14_23; // @[Switch.scala 30:36:@4588.4]
  wire  _T_23116; // @[Switch.scala 30:53:@4590.4]
  wire  valid_14_24; // @[Switch.scala 30:36:@4591.4]
  wire  _T_23119; // @[Switch.scala 30:53:@4593.4]
  wire  valid_14_25; // @[Switch.scala 30:36:@4594.4]
  wire  _T_23122; // @[Switch.scala 30:53:@4596.4]
  wire  valid_14_26; // @[Switch.scala 30:36:@4597.4]
  wire  _T_23125; // @[Switch.scala 30:53:@4599.4]
  wire  valid_14_27; // @[Switch.scala 30:36:@4600.4]
  wire  _T_23128; // @[Switch.scala 30:53:@4602.4]
  wire  valid_14_28; // @[Switch.scala 30:36:@4603.4]
  wire  _T_23131; // @[Switch.scala 30:53:@4605.4]
  wire  valid_14_29; // @[Switch.scala 30:36:@4606.4]
  wire  _T_23134; // @[Switch.scala 30:53:@4608.4]
  wire  valid_14_30; // @[Switch.scala 30:36:@4609.4]
  wire  _T_23137; // @[Switch.scala 30:53:@4611.4]
  wire  valid_14_31; // @[Switch.scala 30:36:@4612.4]
  wire  _T_23140; // @[Switch.scala 30:53:@4614.4]
  wire  valid_14_32; // @[Switch.scala 30:36:@4615.4]
  wire  _T_23143; // @[Switch.scala 30:53:@4617.4]
  wire  valid_14_33; // @[Switch.scala 30:36:@4618.4]
  wire  _T_23146; // @[Switch.scala 30:53:@4620.4]
  wire  valid_14_34; // @[Switch.scala 30:36:@4621.4]
  wire  _T_23149; // @[Switch.scala 30:53:@4623.4]
  wire  valid_14_35; // @[Switch.scala 30:36:@4624.4]
  wire  _T_23152; // @[Switch.scala 30:53:@4626.4]
  wire  valid_14_36; // @[Switch.scala 30:36:@4627.4]
  wire  _T_23155; // @[Switch.scala 30:53:@4629.4]
  wire  valid_14_37; // @[Switch.scala 30:36:@4630.4]
  wire  _T_23158; // @[Switch.scala 30:53:@4632.4]
  wire  valid_14_38; // @[Switch.scala 30:36:@4633.4]
  wire  _T_23161; // @[Switch.scala 30:53:@4635.4]
  wire  valid_14_39; // @[Switch.scala 30:36:@4636.4]
  wire  _T_23164; // @[Switch.scala 30:53:@4638.4]
  wire  valid_14_40; // @[Switch.scala 30:36:@4639.4]
  wire  _T_23167; // @[Switch.scala 30:53:@4641.4]
  wire  valid_14_41; // @[Switch.scala 30:36:@4642.4]
  wire  _T_23170; // @[Switch.scala 30:53:@4644.4]
  wire  valid_14_42; // @[Switch.scala 30:36:@4645.4]
  wire  _T_23173; // @[Switch.scala 30:53:@4647.4]
  wire  valid_14_43; // @[Switch.scala 30:36:@4648.4]
  wire  _T_23176; // @[Switch.scala 30:53:@4650.4]
  wire  valid_14_44; // @[Switch.scala 30:36:@4651.4]
  wire  _T_23179; // @[Switch.scala 30:53:@4653.4]
  wire  valid_14_45; // @[Switch.scala 30:36:@4654.4]
  wire  _T_23182; // @[Switch.scala 30:53:@4656.4]
  wire  valid_14_46; // @[Switch.scala 30:36:@4657.4]
  wire  _T_23185; // @[Switch.scala 30:53:@4659.4]
  wire  valid_14_47; // @[Switch.scala 30:36:@4660.4]
  wire  _T_23188; // @[Switch.scala 30:53:@4662.4]
  wire  valid_14_48; // @[Switch.scala 30:36:@4663.4]
  wire  _T_23191; // @[Switch.scala 30:53:@4665.4]
  wire  valid_14_49; // @[Switch.scala 30:36:@4666.4]
  wire  _T_23194; // @[Switch.scala 30:53:@4668.4]
  wire  valid_14_50; // @[Switch.scala 30:36:@4669.4]
  wire  _T_23197; // @[Switch.scala 30:53:@4671.4]
  wire  valid_14_51; // @[Switch.scala 30:36:@4672.4]
  wire  _T_23200; // @[Switch.scala 30:53:@4674.4]
  wire  valid_14_52; // @[Switch.scala 30:36:@4675.4]
  wire  _T_23203; // @[Switch.scala 30:53:@4677.4]
  wire  valid_14_53; // @[Switch.scala 30:36:@4678.4]
  wire  _T_23206; // @[Switch.scala 30:53:@4680.4]
  wire  valid_14_54; // @[Switch.scala 30:36:@4681.4]
  wire  _T_23209; // @[Switch.scala 30:53:@4683.4]
  wire  valid_14_55; // @[Switch.scala 30:36:@4684.4]
  wire  _T_23212; // @[Switch.scala 30:53:@4686.4]
  wire  valid_14_56; // @[Switch.scala 30:36:@4687.4]
  wire  _T_23215; // @[Switch.scala 30:53:@4689.4]
  wire  valid_14_57; // @[Switch.scala 30:36:@4690.4]
  wire  _T_23218; // @[Switch.scala 30:53:@4692.4]
  wire  valid_14_58; // @[Switch.scala 30:36:@4693.4]
  wire  _T_23221; // @[Switch.scala 30:53:@4695.4]
  wire  valid_14_59; // @[Switch.scala 30:36:@4696.4]
  wire  _T_23224; // @[Switch.scala 30:53:@4698.4]
  wire  valid_14_60; // @[Switch.scala 30:36:@4699.4]
  wire  _T_23227; // @[Switch.scala 30:53:@4701.4]
  wire  valid_14_61; // @[Switch.scala 30:36:@4702.4]
  wire  _T_23230; // @[Switch.scala 30:53:@4704.4]
  wire  valid_14_62; // @[Switch.scala 30:36:@4705.4]
  wire  _T_23233; // @[Switch.scala 30:53:@4707.4]
  wire  valid_14_63; // @[Switch.scala 30:36:@4708.4]
  wire [5:0] _T_23299; // @[Mux.scala 31:69:@4710.4]
  wire [5:0] _T_23300; // @[Mux.scala 31:69:@4711.4]
  wire [5:0] _T_23301; // @[Mux.scala 31:69:@4712.4]
  wire [5:0] _T_23302; // @[Mux.scala 31:69:@4713.4]
  wire [5:0] _T_23303; // @[Mux.scala 31:69:@4714.4]
  wire [5:0] _T_23304; // @[Mux.scala 31:69:@4715.4]
  wire [5:0] _T_23305; // @[Mux.scala 31:69:@4716.4]
  wire [5:0] _T_23306; // @[Mux.scala 31:69:@4717.4]
  wire [5:0] _T_23307; // @[Mux.scala 31:69:@4718.4]
  wire [5:0] _T_23308; // @[Mux.scala 31:69:@4719.4]
  wire [5:0] _T_23309; // @[Mux.scala 31:69:@4720.4]
  wire [5:0] _T_23310; // @[Mux.scala 31:69:@4721.4]
  wire [5:0] _T_23311; // @[Mux.scala 31:69:@4722.4]
  wire [5:0] _T_23312; // @[Mux.scala 31:69:@4723.4]
  wire [5:0] _T_23313; // @[Mux.scala 31:69:@4724.4]
  wire [5:0] _T_23314; // @[Mux.scala 31:69:@4725.4]
  wire [5:0] _T_23315; // @[Mux.scala 31:69:@4726.4]
  wire [5:0] _T_23316; // @[Mux.scala 31:69:@4727.4]
  wire [5:0] _T_23317; // @[Mux.scala 31:69:@4728.4]
  wire [5:0] _T_23318; // @[Mux.scala 31:69:@4729.4]
  wire [5:0] _T_23319; // @[Mux.scala 31:69:@4730.4]
  wire [5:0] _T_23320; // @[Mux.scala 31:69:@4731.4]
  wire [5:0] _T_23321; // @[Mux.scala 31:69:@4732.4]
  wire [5:0] _T_23322; // @[Mux.scala 31:69:@4733.4]
  wire [5:0] _T_23323; // @[Mux.scala 31:69:@4734.4]
  wire [5:0] _T_23324; // @[Mux.scala 31:69:@4735.4]
  wire [5:0] _T_23325; // @[Mux.scala 31:69:@4736.4]
  wire [5:0] _T_23326; // @[Mux.scala 31:69:@4737.4]
  wire [5:0] _T_23327; // @[Mux.scala 31:69:@4738.4]
  wire [5:0] _T_23328; // @[Mux.scala 31:69:@4739.4]
  wire [5:0] _T_23329; // @[Mux.scala 31:69:@4740.4]
  wire [5:0] _T_23330; // @[Mux.scala 31:69:@4741.4]
  wire [5:0] _T_23331; // @[Mux.scala 31:69:@4742.4]
  wire [5:0] _T_23332; // @[Mux.scala 31:69:@4743.4]
  wire [5:0] _T_23333; // @[Mux.scala 31:69:@4744.4]
  wire [5:0] _T_23334; // @[Mux.scala 31:69:@4745.4]
  wire [5:0] _T_23335; // @[Mux.scala 31:69:@4746.4]
  wire [5:0] _T_23336; // @[Mux.scala 31:69:@4747.4]
  wire [5:0] _T_23337; // @[Mux.scala 31:69:@4748.4]
  wire [5:0] _T_23338; // @[Mux.scala 31:69:@4749.4]
  wire [5:0] _T_23339; // @[Mux.scala 31:69:@4750.4]
  wire [5:0] _T_23340; // @[Mux.scala 31:69:@4751.4]
  wire [5:0] _T_23341; // @[Mux.scala 31:69:@4752.4]
  wire [5:0] _T_23342; // @[Mux.scala 31:69:@4753.4]
  wire [5:0] _T_23343; // @[Mux.scala 31:69:@4754.4]
  wire [5:0] _T_23344; // @[Mux.scala 31:69:@4755.4]
  wire [5:0] _T_23345; // @[Mux.scala 31:69:@4756.4]
  wire [5:0] _T_23346; // @[Mux.scala 31:69:@4757.4]
  wire [5:0] _T_23347; // @[Mux.scala 31:69:@4758.4]
  wire [5:0] _T_23348; // @[Mux.scala 31:69:@4759.4]
  wire [5:0] _T_23349; // @[Mux.scala 31:69:@4760.4]
  wire [5:0] _T_23350; // @[Mux.scala 31:69:@4761.4]
  wire [5:0] _T_23351; // @[Mux.scala 31:69:@4762.4]
  wire [5:0] _T_23352; // @[Mux.scala 31:69:@4763.4]
  wire [5:0] _T_23353; // @[Mux.scala 31:69:@4764.4]
  wire [5:0] _T_23354; // @[Mux.scala 31:69:@4765.4]
  wire [5:0] _T_23355; // @[Mux.scala 31:69:@4766.4]
  wire [5:0] _T_23356; // @[Mux.scala 31:69:@4767.4]
  wire [5:0] _T_23357; // @[Mux.scala 31:69:@4768.4]
  wire [5:0] _T_23358; // @[Mux.scala 31:69:@4769.4]
  wire [5:0] _T_23359; // @[Mux.scala 31:69:@4770.4]
  wire [5:0] _T_23360; // @[Mux.scala 31:69:@4771.4]
  wire [5:0] select_14; // @[Mux.scala 31:69:@4772.4]
  wire [47:0] _GEN_897; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_898; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_899; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_900; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_901; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_902; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_903; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_904; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_905; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_906; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_907; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_908; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_909; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_910; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_911; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_912; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_913; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_914; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_915; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_916; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_917; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_918; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_919; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_920; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_921; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_922; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_923; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_924; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_925; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_926; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_927; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_928; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_929; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_930; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_931; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_932; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_933; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_934; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_935; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_936; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_937; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_938; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_939; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_940; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_941; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_942; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_943; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_944; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_945; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_946; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_947; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_948; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_949; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_950; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_951; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_952; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_953; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_954; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_955; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_956; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_957; // @[Switch.scala 33:19:@4774.4]
  wire [47:0] _GEN_958; // @[Switch.scala 33:19:@4774.4]
  wire [7:0] _T_23369; // @[Switch.scala 34:32:@4781.4]
  wire [15:0] _T_23377; // @[Switch.scala 34:32:@4789.4]
  wire [7:0] _T_23384; // @[Switch.scala 34:32:@4796.4]
  wire [31:0] _T_23393; // @[Switch.scala 34:32:@4805.4]
  wire [7:0] _T_23400; // @[Switch.scala 34:32:@4812.4]
  wire [15:0] _T_23408; // @[Switch.scala 34:32:@4820.4]
  wire [7:0] _T_23415; // @[Switch.scala 34:32:@4827.4]
  wire [31:0] _T_23424; // @[Switch.scala 34:32:@4836.4]
  wire [63:0] _T_23425; // @[Switch.scala 34:32:@4837.4]
  wire  _T_23429; // @[Switch.scala 30:53:@4840.4]
  wire  valid_15_0; // @[Switch.scala 30:36:@4841.4]
  wire  _T_23432; // @[Switch.scala 30:53:@4843.4]
  wire  valid_15_1; // @[Switch.scala 30:36:@4844.4]
  wire  _T_23435; // @[Switch.scala 30:53:@4846.4]
  wire  valid_15_2; // @[Switch.scala 30:36:@4847.4]
  wire  _T_23438; // @[Switch.scala 30:53:@4849.4]
  wire  valid_15_3; // @[Switch.scala 30:36:@4850.4]
  wire  _T_23441; // @[Switch.scala 30:53:@4852.4]
  wire  valid_15_4; // @[Switch.scala 30:36:@4853.4]
  wire  _T_23444; // @[Switch.scala 30:53:@4855.4]
  wire  valid_15_5; // @[Switch.scala 30:36:@4856.4]
  wire  _T_23447; // @[Switch.scala 30:53:@4858.4]
  wire  valid_15_6; // @[Switch.scala 30:36:@4859.4]
  wire  _T_23450; // @[Switch.scala 30:53:@4861.4]
  wire  valid_15_7; // @[Switch.scala 30:36:@4862.4]
  wire  _T_23453; // @[Switch.scala 30:53:@4864.4]
  wire  valid_15_8; // @[Switch.scala 30:36:@4865.4]
  wire  _T_23456; // @[Switch.scala 30:53:@4867.4]
  wire  valid_15_9; // @[Switch.scala 30:36:@4868.4]
  wire  _T_23459; // @[Switch.scala 30:53:@4870.4]
  wire  valid_15_10; // @[Switch.scala 30:36:@4871.4]
  wire  _T_23462; // @[Switch.scala 30:53:@4873.4]
  wire  valid_15_11; // @[Switch.scala 30:36:@4874.4]
  wire  _T_23465; // @[Switch.scala 30:53:@4876.4]
  wire  valid_15_12; // @[Switch.scala 30:36:@4877.4]
  wire  _T_23468; // @[Switch.scala 30:53:@4879.4]
  wire  valid_15_13; // @[Switch.scala 30:36:@4880.4]
  wire  _T_23471; // @[Switch.scala 30:53:@4882.4]
  wire  valid_15_14; // @[Switch.scala 30:36:@4883.4]
  wire  _T_23474; // @[Switch.scala 30:53:@4885.4]
  wire  valid_15_15; // @[Switch.scala 30:36:@4886.4]
  wire  _T_23477; // @[Switch.scala 30:53:@4888.4]
  wire  valid_15_16; // @[Switch.scala 30:36:@4889.4]
  wire  _T_23480; // @[Switch.scala 30:53:@4891.4]
  wire  valid_15_17; // @[Switch.scala 30:36:@4892.4]
  wire  _T_23483; // @[Switch.scala 30:53:@4894.4]
  wire  valid_15_18; // @[Switch.scala 30:36:@4895.4]
  wire  _T_23486; // @[Switch.scala 30:53:@4897.4]
  wire  valid_15_19; // @[Switch.scala 30:36:@4898.4]
  wire  _T_23489; // @[Switch.scala 30:53:@4900.4]
  wire  valid_15_20; // @[Switch.scala 30:36:@4901.4]
  wire  _T_23492; // @[Switch.scala 30:53:@4903.4]
  wire  valid_15_21; // @[Switch.scala 30:36:@4904.4]
  wire  _T_23495; // @[Switch.scala 30:53:@4906.4]
  wire  valid_15_22; // @[Switch.scala 30:36:@4907.4]
  wire  _T_23498; // @[Switch.scala 30:53:@4909.4]
  wire  valid_15_23; // @[Switch.scala 30:36:@4910.4]
  wire  _T_23501; // @[Switch.scala 30:53:@4912.4]
  wire  valid_15_24; // @[Switch.scala 30:36:@4913.4]
  wire  _T_23504; // @[Switch.scala 30:53:@4915.4]
  wire  valid_15_25; // @[Switch.scala 30:36:@4916.4]
  wire  _T_23507; // @[Switch.scala 30:53:@4918.4]
  wire  valid_15_26; // @[Switch.scala 30:36:@4919.4]
  wire  _T_23510; // @[Switch.scala 30:53:@4921.4]
  wire  valid_15_27; // @[Switch.scala 30:36:@4922.4]
  wire  _T_23513; // @[Switch.scala 30:53:@4924.4]
  wire  valid_15_28; // @[Switch.scala 30:36:@4925.4]
  wire  _T_23516; // @[Switch.scala 30:53:@4927.4]
  wire  valid_15_29; // @[Switch.scala 30:36:@4928.4]
  wire  _T_23519; // @[Switch.scala 30:53:@4930.4]
  wire  valid_15_30; // @[Switch.scala 30:36:@4931.4]
  wire  _T_23522; // @[Switch.scala 30:53:@4933.4]
  wire  valid_15_31; // @[Switch.scala 30:36:@4934.4]
  wire  _T_23525; // @[Switch.scala 30:53:@4936.4]
  wire  valid_15_32; // @[Switch.scala 30:36:@4937.4]
  wire  _T_23528; // @[Switch.scala 30:53:@4939.4]
  wire  valid_15_33; // @[Switch.scala 30:36:@4940.4]
  wire  _T_23531; // @[Switch.scala 30:53:@4942.4]
  wire  valid_15_34; // @[Switch.scala 30:36:@4943.4]
  wire  _T_23534; // @[Switch.scala 30:53:@4945.4]
  wire  valid_15_35; // @[Switch.scala 30:36:@4946.4]
  wire  _T_23537; // @[Switch.scala 30:53:@4948.4]
  wire  valid_15_36; // @[Switch.scala 30:36:@4949.4]
  wire  _T_23540; // @[Switch.scala 30:53:@4951.4]
  wire  valid_15_37; // @[Switch.scala 30:36:@4952.4]
  wire  _T_23543; // @[Switch.scala 30:53:@4954.4]
  wire  valid_15_38; // @[Switch.scala 30:36:@4955.4]
  wire  _T_23546; // @[Switch.scala 30:53:@4957.4]
  wire  valid_15_39; // @[Switch.scala 30:36:@4958.4]
  wire  _T_23549; // @[Switch.scala 30:53:@4960.4]
  wire  valid_15_40; // @[Switch.scala 30:36:@4961.4]
  wire  _T_23552; // @[Switch.scala 30:53:@4963.4]
  wire  valid_15_41; // @[Switch.scala 30:36:@4964.4]
  wire  _T_23555; // @[Switch.scala 30:53:@4966.4]
  wire  valid_15_42; // @[Switch.scala 30:36:@4967.4]
  wire  _T_23558; // @[Switch.scala 30:53:@4969.4]
  wire  valid_15_43; // @[Switch.scala 30:36:@4970.4]
  wire  _T_23561; // @[Switch.scala 30:53:@4972.4]
  wire  valid_15_44; // @[Switch.scala 30:36:@4973.4]
  wire  _T_23564; // @[Switch.scala 30:53:@4975.4]
  wire  valid_15_45; // @[Switch.scala 30:36:@4976.4]
  wire  _T_23567; // @[Switch.scala 30:53:@4978.4]
  wire  valid_15_46; // @[Switch.scala 30:36:@4979.4]
  wire  _T_23570; // @[Switch.scala 30:53:@4981.4]
  wire  valid_15_47; // @[Switch.scala 30:36:@4982.4]
  wire  _T_23573; // @[Switch.scala 30:53:@4984.4]
  wire  valid_15_48; // @[Switch.scala 30:36:@4985.4]
  wire  _T_23576; // @[Switch.scala 30:53:@4987.4]
  wire  valid_15_49; // @[Switch.scala 30:36:@4988.4]
  wire  _T_23579; // @[Switch.scala 30:53:@4990.4]
  wire  valid_15_50; // @[Switch.scala 30:36:@4991.4]
  wire  _T_23582; // @[Switch.scala 30:53:@4993.4]
  wire  valid_15_51; // @[Switch.scala 30:36:@4994.4]
  wire  _T_23585; // @[Switch.scala 30:53:@4996.4]
  wire  valid_15_52; // @[Switch.scala 30:36:@4997.4]
  wire  _T_23588; // @[Switch.scala 30:53:@4999.4]
  wire  valid_15_53; // @[Switch.scala 30:36:@5000.4]
  wire  _T_23591; // @[Switch.scala 30:53:@5002.4]
  wire  valid_15_54; // @[Switch.scala 30:36:@5003.4]
  wire  _T_23594; // @[Switch.scala 30:53:@5005.4]
  wire  valid_15_55; // @[Switch.scala 30:36:@5006.4]
  wire  _T_23597; // @[Switch.scala 30:53:@5008.4]
  wire  valid_15_56; // @[Switch.scala 30:36:@5009.4]
  wire  _T_23600; // @[Switch.scala 30:53:@5011.4]
  wire  valid_15_57; // @[Switch.scala 30:36:@5012.4]
  wire  _T_23603; // @[Switch.scala 30:53:@5014.4]
  wire  valid_15_58; // @[Switch.scala 30:36:@5015.4]
  wire  _T_23606; // @[Switch.scala 30:53:@5017.4]
  wire  valid_15_59; // @[Switch.scala 30:36:@5018.4]
  wire  _T_23609; // @[Switch.scala 30:53:@5020.4]
  wire  valid_15_60; // @[Switch.scala 30:36:@5021.4]
  wire  _T_23612; // @[Switch.scala 30:53:@5023.4]
  wire  valid_15_61; // @[Switch.scala 30:36:@5024.4]
  wire  _T_23615; // @[Switch.scala 30:53:@5026.4]
  wire  valid_15_62; // @[Switch.scala 30:36:@5027.4]
  wire  _T_23618; // @[Switch.scala 30:53:@5029.4]
  wire  valid_15_63; // @[Switch.scala 30:36:@5030.4]
  wire [5:0] _T_23684; // @[Mux.scala 31:69:@5032.4]
  wire [5:0] _T_23685; // @[Mux.scala 31:69:@5033.4]
  wire [5:0] _T_23686; // @[Mux.scala 31:69:@5034.4]
  wire [5:0] _T_23687; // @[Mux.scala 31:69:@5035.4]
  wire [5:0] _T_23688; // @[Mux.scala 31:69:@5036.4]
  wire [5:0] _T_23689; // @[Mux.scala 31:69:@5037.4]
  wire [5:0] _T_23690; // @[Mux.scala 31:69:@5038.4]
  wire [5:0] _T_23691; // @[Mux.scala 31:69:@5039.4]
  wire [5:0] _T_23692; // @[Mux.scala 31:69:@5040.4]
  wire [5:0] _T_23693; // @[Mux.scala 31:69:@5041.4]
  wire [5:0] _T_23694; // @[Mux.scala 31:69:@5042.4]
  wire [5:0] _T_23695; // @[Mux.scala 31:69:@5043.4]
  wire [5:0] _T_23696; // @[Mux.scala 31:69:@5044.4]
  wire [5:0] _T_23697; // @[Mux.scala 31:69:@5045.4]
  wire [5:0] _T_23698; // @[Mux.scala 31:69:@5046.4]
  wire [5:0] _T_23699; // @[Mux.scala 31:69:@5047.4]
  wire [5:0] _T_23700; // @[Mux.scala 31:69:@5048.4]
  wire [5:0] _T_23701; // @[Mux.scala 31:69:@5049.4]
  wire [5:0] _T_23702; // @[Mux.scala 31:69:@5050.4]
  wire [5:0] _T_23703; // @[Mux.scala 31:69:@5051.4]
  wire [5:0] _T_23704; // @[Mux.scala 31:69:@5052.4]
  wire [5:0] _T_23705; // @[Mux.scala 31:69:@5053.4]
  wire [5:0] _T_23706; // @[Mux.scala 31:69:@5054.4]
  wire [5:0] _T_23707; // @[Mux.scala 31:69:@5055.4]
  wire [5:0] _T_23708; // @[Mux.scala 31:69:@5056.4]
  wire [5:0] _T_23709; // @[Mux.scala 31:69:@5057.4]
  wire [5:0] _T_23710; // @[Mux.scala 31:69:@5058.4]
  wire [5:0] _T_23711; // @[Mux.scala 31:69:@5059.4]
  wire [5:0] _T_23712; // @[Mux.scala 31:69:@5060.4]
  wire [5:0] _T_23713; // @[Mux.scala 31:69:@5061.4]
  wire [5:0] _T_23714; // @[Mux.scala 31:69:@5062.4]
  wire [5:0] _T_23715; // @[Mux.scala 31:69:@5063.4]
  wire [5:0] _T_23716; // @[Mux.scala 31:69:@5064.4]
  wire [5:0] _T_23717; // @[Mux.scala 31:69:@5065.4]
  wire [5:0] _T_23718; // @[Mux.scala 31:69:@5066.4]
  wire [5:0] _T_23719; // @[Mux.scala 31:69:@5067.4]
  wire [5:0] _T_23720; // @[Mux.scala 31:69:@5068.4]
  wire [5:0] _T_23721; // @[Mux.scala 31:69:@5069.4]
  wire [5:0] _T_23722; // @[Mux.scala 31:69:@5070.4]
  wire [5:0] _T_23723; // @[Mux.scala 31:69:@5071.4]
  wire [5:0] _T_23724; // @[Mux.scala 31:69:@5072.4]
  wire [5:0] _T_23725; // @[Mux.scala 31:69:@5073.4]
  wire [5:0] _T_23726; // @[Mux.scala 31:69:@5074.4]
  wire [5:0] _T_23727; // @[Mux.scala 31:69:@5075.4]
  wire [5:0] _T_23728; // @[Mux.scala 31:69:@5076.4]
  wire [5:0] _T_23729; // @[Mux.scala 31:69:@5077.4]
  wire [5:0] _T_23730; // @[Mux.scala 31:69:@5078.4]
  wire [5:0] _T_23731; // @[Mux.scala 31:69:@5079.4]
  wire [5:0] _T_23732; // @[Mux.scala 31:69:@5080.4]
  wire [5:0] _T_23733; // @[Mux.scala 31:69:@5081.4]
  wire [5:0] _T_23734; // @[Mux.scala 31:69:@5082.4]
  wire [5:0] _T_23735; // @[Mux.scala 31:69:@5083.4]
  wire [5:0] _T_23736; // @[Mux.scala 31:69:@5084.4]
  wire [5:0] _T_23737; // @[Mux.scala 31:69:@5085.4]
  wire [5:0] _T_23738; // @[Mux.scala 31:69:@5086.4]
  wire [5:0] _T_23739; // @[Mux.scala 31:69:@5087.4]
  wire [5:0] _T_23740; // @[Mux.scala 31:69:@5088.4]
  wire [5:0] _T_23741; // @[Mux.scala 31:69:@5089.4]
  wire [5:0] _T_23742; // @[Mux.scala 31:69:@5090.4]
  wire [5:0] _T_23743; // @[Mux.scala 31:69:@5091.4]
  wire [5:0] _T_23744; // @[Mux.scala 31:69:@5092.4]
  wire [5:0] _T_23745; // @[Mux.scala 31:69:@5093.4]
  wire [5:0] select_15; // @[Mux.scala 31:69:@5094.4]
  wire [47:0] _GEN_961; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_962; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_963; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_964; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_965; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_966; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_967; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_968; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_969; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_970; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_971; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_972; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_973; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_974; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_975; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_976; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_977; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_978; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_979; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_980; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_981; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_982; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_983; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_984; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_985; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_986; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_987; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_988; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_989; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_990; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_991; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_992; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_993; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_994; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_995; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_996; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_997; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_998; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_999; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_1000; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_1001; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_1002; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_1003; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_1004; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_1005; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_1006; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_1007; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_1008; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_1009; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_1010; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_1011; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_1012; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_1013; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_1014; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_1015; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_1016; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_1017; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_1018; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_1019; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_1020; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_1021; // @[Switch.scala 33:19:@5096.4]
  wire [47:0] _GEN_1022; // @[Switch.scala 33:19:@5096.4]
  wire [7:0] _T_23754; // @[Switch.scala 34:32:@5103.4]
  wire [15:0] _T_23762; // @[Switch.scala 34:32:@5111.4]
  wire [7:0] _T_23769; // @[Switch.scala 34:32:@5118.4]
  wire [31:0] _T_23778; // @[Switch.scala 34:32:@5127.4]
  wire [7:0] _T_23785; // @[Switch.scala 34:32:@5134.4]
  wire [15:0] _T_23793; // @[Switch.scala 34:32:@5142.4]
  wire [7:0] _T_23800; // @[Switch.scala 34:32:@5149.4]
  wire [31:0] _T_23809; // @[Switch.scala 34:32:@5158.4]
  wire [63:0] _T_23810; // @[Switch.scala 34:32:@5159.4]
  wire  _T_23814; // @[Switch.scala 30:53:@5162.4]
  wire  valid_16_0; // @[Switch.scala 30:36:@5163.4]
  wire  _T_23817; // @[Switch.scala 30:53:@5165.4]
  wire  valid_16_1; // @[Switch.scala 30:36:@5166.4]
  wire  _T_23820; // @[Switch.scala 30:53:@5168.4]
  wire  valid_16_2; // @[Switch.scala 30:36:@5169.4]
  wire  _T_23823; // @[Switch.scala 30:53:@5171.4]
  wire  valid_16_3; // @[Switch.scala 30:36:@5172.4]
  wire  _T_23826; // @[Switch.scala 30:53:@5174.4]
  wire  valid_16_4; // @[Switch.scala 30:36:@5175.4]
  wire  _T_23829; // @[Switch.scala 30:53:@5177.4]
  wire  valid_16_5; // @[Switch.scala 30:36:@5178.4]
  wire  _T_23832; // @[Switch.scala 30:53:@5180.4]
  wire  valid_16_6; // @[Switch.scala 30:36:@5181.4]
  wire  _T_23835; // @[Switch.scala 30:53:@5183.4]
  wire  valid_16_7; // @[Switch.scala 30:36:@5184.4]
  wire  _T_23838; // @[Switch.scala 30:53:@5186.4]
  wire  valid_16_8; // @[Switch.scala 30:36:@5187.4]
  wire  _T_23841; // @[Switch.scala 30:53:@5189.4]
  wire  valid_16_9; // @[Switch.scala 30:36:@5190.4]
  wire  _T_23844; // @[Switch.scala 30:53:@5192.4]
  wire  valid_16_10; // @[Switch.scala 30:36:@5193.4]
  wire  _T_23847; // @[Switch.scala 30:53:@5195.4]
  wire  valid_16_11; // @[Switch.scala 30:36:@5196.4]
  wire  _T_23850; // @[Switch.scala 30:53:@5198.4]
  wire  valid_16_12; // @[Switch.scala 30:36:@5199.4]
  wire  _T_23853; // @[Switch.scala 30:53:@5201.4]
  wire  valid_16_13; // @[Switch.scala 30:36:@5202.4]
  wire  _T_23856; // @[Switch.scala 30:53:@5204.4]
  wire  valid_16_14; // @[Switch.scala 30:36:@5205.4]
  wire  _T_23859; // @[Switch.scala 30:53:@5207.4]
  wire  valid_16_15; // @[Switch.scala 30:36:@5208.4]
  wire  _T_23862; // @[Switch.scala 30:53:@5210.4]
  wire  valid_16_16; // @[Switch.scala 30:36:@5211.4]
  wire  _T_23865; // @[Switch.scala 30:53:@5213.4]
  wire  valid_16_17; // @[Switch.scala 30:36:@5214.4]
  wire  _T_23868; // @[Switch.scala 30:53:@5216.4]
  wire  valid_16_18; // @[Switch.scala 30:36:@5217.4]
  wire  _T_23871; // @[Switch.scala 30:53:@5219.4]
  wire  valid_16_19; // @[Switch.scala 30:36:@5220.4]
  wire  _T_23874; // @[Switch.scala 30:53:@5222.4]
  wire  valid_16_20; // @[Switch.scala 30:36:@5223.4]
  wire  _T_23877; // @[Switch.scala 30:53:@5225.4]
  wire  valid_16_21; // @[Switch.scala 30:36:@5226.4]
  wire  _T_23880; // @[Switch.scala 30:53:@5228.4]
  wire  valid_16_22; // @[Switch.scala 30:36:@5229.4]
  wire  _T_23883; // @[Switch.scala 30:53:@5231.4]
  wire  valid_16_23; // @[Switch.scala 30:36:@5232.4]
  wire  _T_23886; // @[Switch.scala 30:53:@5234.4]
  wire  valid_16_24; // @[Switch.scala 30:36:@5235.4]
  wire  _T_23889; // @[Switch.scala 30:53:@5237.4]
  wire  valid_16_25; // @[Switch.scala 30:36:@5238.4]
  wire  _T_23892; // @[Switch.scala 30:53:@5240.4]
  wire  valid_16_26; // @[Switch.scala 30:36:@5241.4]
  wire  _T_23895; // @[Switch.scala 30:53:@5243.4]
  wire  valid_16_27; // @[Switch.scala 30:36:@5244.4]
  wire  _T_23898; // @[Switch.scala 30:53:@5246.4]
  wire  valid_16_28; // @[Switch.scala 30:36:@5247.4]
  wire  _T_23901; // @[Switch.scala 30:53:@5249.4]
  wire  valid_16_29; // @[Switch.scala 30:36:@5250.4]
  wire  _T_23904; // @[Switch.scala 30:53:@5252.4]
  wire  valid_16_30; // @[Switch.scala 30:36:@5253.4]
  wire  _T_23907; // @[Switch.scala 30:53:@5255.4]
  wire  valid_16_31; // @[Switch.scala 30:36:@5256.4]
  wire  _T_23910; // @[Switch.scala 30:53:@5258.4]
  wire  valid_16_32; // @[Switch.scala 30:36:@5259.4]
  wire  _T_23913; // @[Switch.scala 30:53:@5261.4]
  wire  valid_16_33; // @[Switch.scala 30:36:@5262.4]
  wire  _T_23916; // @[Switch.scala 30:53:@5264.4]
  wire  valid_16_34; // @[Switch.scala 30:36:@5265.4]
  wire  _T_23919; // @[Switch.scala 30:53:@5267.4]
  wire  valid_16_35; // @[Switch.scala 30:36:@5268.4]
  wire  _T_23922; // @[Switch.scala 30:53:@5270.4]
  wire  valid_16_36; // @[Switch.scala 30:36:@5271.4]
  wire  _T_23925; // @[Switch.scala 30:53:@5273.4]
  wire  valid_16_37; // @[Switch.scala 30:36:@5274.4]
  wire  _T_23928; // @[Switch.scala 30:53:@5276.4]
  wire  valid_16_38; // @[Switch.scala 30:36:@5277.4]
  wire  _T_23931; // @[Switch.scala 30:53:@5279.4]
  wire  valid_16_39; // @[Switch.scala 30:36:@5280.4]
  wire  _T_23934; // @[Switch.scala 30:53:@5282.4]
  wire  valid_16_40; // @[Switch.scala 30:36:@5283.4]
  wire  _T_23937; // @[Switch.scala 30:53:@5285.4]
  wire  valid_16_41; // @[Switch.scala 30:36:@5286.4]
  wire  _T_23940; // @[Switch.scala 30:53:@5288.4]
  wire  valid_16_42; // @[Switch.scala 30:36:@5289.4]
  wire  _T_23943; // @[Switch.scala 30:53:@5291.4]
  wire  valid_16_43; // @[Switch.scala 30:36:@5292.4]
  wire  _T_23946; // @[Switch.scala 30:53:@5294.4]
  wire  valid_16_44; // @[Switch.scala 30:36:@5295.4]
  wire  _T_23949; // @[Switch.scala 30:53:@5297.4]
  wire  valid_16_45; // @[Switch.scala 30:36:@5298.4]
  wire  _T_23952; // @[Switch.scala 30:53:@5300.4]
  wire  valid_16_46; // @[Switch.scala 30:36:@5301.4]
  wire  _T_23955; // @[Switch.scala 30:53:@5303.4]
  wire  valid_16_47; // @[Switch.scala 30:36:@5304.4]
  wire  _T_23958; // @[Switch.scala 30:53:@5306.4]
  wire  valid_16_48; // @[Switch.scala 30:36:@5307.4]
  wire  _T_23961; // @[Switch.scala 30:53:@5309.4]
  wire  valid_16_49; // @[Switch.scala 30:36:@5310.4]
  wire  _T_23964; // @[Switch.scala 30:53:@5312.4]
  wire  valid_16_50; // @[Switch.scala 30:36:@5313.4]
  wire  _T_23967; // @[Switch.scala 30:53:@5315.4]
  wire  valid_16_51; // @[Switch.scala 30:36:@5316.4]
  wire  _T_23970; // @[Switch.scala 30:53:@5318.4]
  wire  valid_16_52; // @[Switch.scala 30:36:@5319.4]
  wire  _T_23973; // @[Switch.scala 30:53:@5321.4]
  wire  valid_16_53; // @[Switch.scala 30:36:@5322.4]
  wire  _T_23976; // @[Switch.scala 30:53:@5324.4]
  wire  valid_16_54; // @[Switch.scala 30:36:@5325.4]
  wire  _T_23979; // @[Switch.scala 30:53:@5327.4]
  wire  valid_16_55; // @[Switch.scala 30:36:@5328.4]
  wire  _T_23982; // @[Switch.scala 30:53:@5330.4]
  wire  valid_16_56; // @[Switch.scala 30:36:@5331.4]
  wire  _T_23985; // @[Switch.scala 30:53:@5333.4]
  wire  valid_16_57; // @[Switch.scala 30:36:@5334.4]
  wire  _T_23988; // @[Switch.scala 30:53:@5336.4]
  wire  valid_16_58; // @[Switch.scala 30:36:@5337.4]
  wire  _T_23991; // @[Switch.scala 30:53:@5339.4]
  wire  valid_16_59; // @[Switch.scala 30:36:@5340.4]
  wire  _T_23994; // @[Switch.scala 30:53:@5342.4]
  wire  valid_16_60; // @[Switch.scala 30:36:@5343.4]
  wire  _T_23997; // @[Switch.scala 30:53:@5345.4]
  wire  valid_16_61; // @[Switch.scala 30:36:@5346.4]
  wire  _T_24000; // @[Switch.scala 30:53:@5348.4]
  wire  valid_16_62; // @[Switch.scala 30:36:@5349.4]
  wire  _T_24003; // @[Switch.scala 30:53:@5351.4]
  wire  valid_16_63; // @[Switch.scala 30:36:@5352.4]
  wire [5:0] _T_24069; // @[Mux.scala 31:69:@5354.4]
  wire [5:0] _T_24070; // @[Mux.scala 31:69:@5355.4]
  wire [5:0] _T_24071; // @[Mux.scala 31:69:@5356.4]
  wire [5:0] _T_24072; // @[Mux.scala 31:69:@5357.4]
  wire [5:0] _T_24073; // @[Mux.scala 31:69:@5358.4]
  wire [5:0] _T_24074; // @[Mux.scala 31:69:@5359.4]
  wire [5:0] _T_24075; // @[Mux.scala 31:69:@5360.4]
  wire [5:0] _T_24076; // @[Mux.scala 31:69:@5361.4]
  wire [5:0] _T_24077; // @[Mux.scala 31:69:@5362.4]
  wire [5:0] _T_24078; // @[Mux.scala 31:69:@5363.4]
  wire [5:0] _T_24079; // @[Mux.scala 31:69:@5364.4]
  wire [5:0] _T_24080; // @[Mux.scala 31:69:@5365.4]
  wire [5:0] _T_24081; // @[Mux.scala 31:69:@5366.4]
  wire [5:0] _T_24082; // @[Mux.scala 31:69:@5367.4]
  wire [5:0] _T_24083; // @[Mux.scala 31:69:@5368.4]
  wire [5:0] _T_24084; // @[Mux.scala 31:69:@5369.4]
  wire [5:0] _T_24085; // @[Mux.scala 31:69:@5370.4]
  wire [5:0] _T_24086; // @[Mux.scala 31:69:@5371.4]
  wire [5:0] _T_24087; // @[Mux.scala 31:69:@5372.4]
  wire [5:0] _T_24088; // @[Mux.scala 31:69:@5373.4]
  wire [5:0] _T_24089; // @[Mux.scala 31:69:@5374.4]
  wire [5:0] _T_24090; // @[Mux.scala 31:69:@5375.4]
  wire [5:0] _T_24091; // @[Mux.scala 31:69:@5376.4]
  wire [5:0] _T_24092; // @[Mux.scala 31:69:@5377.4]
  wire [5:0] _T_24093; // @[Mux.scala 31:69:@5378.4]
  wire [5:0] _T_24094; // @[Mux.scala 31:69:@5379.4]
  wire [5:0] _T_24095; // @[Mux.scala 31:69:@5380.4]
  wire [5:0] _T_24096; // @[Mux.scala 31:69:@5381.4]
  wire [5:0] _T_24097; // @[Mux.scala 31:69:@5382.4]
  wire [5:0] _T_24098; // @[Mux.scala 31:69:@5383.4]
  wire [5:0] _T_24099; // @[Mux.scala 31:69:@5384.4]
  wire [5:0] _T_24100; // @[Mux.scala 31:69:@5385.4]
  wire [5:0] _T_24101; // @[Mux.scala 31:69:@5386.4]
  wire [5:0] _T_24102; // @[Mux.scala 31:69:@5387.4]
  wire [5:0] _T_24103; // @[Mux.scala 31:69:@5388.4]
  wire [5:0] _T_24104; // @[Mux.scala 31:69:@5389.4]
  wire [5:0] _T_24105; // @[Mux.scala 31:69:@5390.4]
  wire [5:0] _T_24106; // @[Mux.scala 31:69:@5391.4]
  wire [5:0] _T_24107; // @[Mux.scala 31:69:@5392.4]
  wire [5:0] _T_24108; // @[Mux.scala 31:69:@5393.4]
  wire [5:0] _T_24109; // @[Mux.scala 31:69:@5394.4]
  wire [5:0] _T_24110; // @[Mux.scala 31:69:@5395.4]
  wire [5:0] _T_24111; // @[Mux.scala 31:69:@5396.4]
  wire [5:0] _T_24112; // @[Mux.scala 31:69:@5397.4]
  wire [5:0] _T_24113; // @[Mux.scala 31:69:@5398.4]
  wire [5:0] _T_24114; // @[Mux.scala 31:69:@5399.4]
  wire [5:0] _T_24115; // @[Mux.scala 31:69:@5400.4]
  wire [5:0] _T_24116; // @[Mux.scala 31:69:@5401.4]
  wire [5:0] _T_24117; // @[Mux.scala 31:69:@5402.4]
  wire [5:0] _T_24118; // @[Mux.scala 31:69:@5403.4]
  wire [5:0] _T_24119; // @[Mux.scala 31:69:@5404.4]
  wire [5:0] _T_24120; // @[Mux.scala 31:69:@5405.4]
  wire [5:0] _T_24121; // @[Mux.scala 31:69:@5406.4]
  wire [5:0] _T_24122; // @[Mux.scala 31:69:@5407.4]
  wire [5:0] _T_24123; // @[Mux.scala 31:69:@5408.4]
  wire [5:0] _T_24124; // @[Mux.scala 31:69:@5409.4]
  wire [5:0] _T_24125; // @[Mux.scala 31:69:@5410.4]
  wire [5:0] _T_24126; // @[Mux.scala 31:69:@5411.4]
  wire [5:0] _T_24127; // @[Mux.scala 31:69:@5412.4]
  wire [5:0] _T_24128; // @[Mux.scala 31:69:@5413.4]
  wire [5:0] _T_24129; // @[Mux.scala 31:69:@5414.4]
  wire [5:0] _T_24130; // @[Mux.scala 31:69:@5415.4]
  wire [5:0] select_16; // @[Mux.scala 31:69:@5416.4]
  wire [47:0] _GEN_1025; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1026; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1027; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1028; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1029; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1030; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1031; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1032; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1033; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1034; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1035; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1036; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1037; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1038; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1039; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1040; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1041; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1042; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1043; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1044; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1045; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1046; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1047; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1048; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1049; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1050; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1051; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1052; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1053; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1054; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1055; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1056; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1057; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1058; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1059; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1060; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1061; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1062; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1063; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1064; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1065; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1066; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1067; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1068; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1069; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1070; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1071; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1072; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1073; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1074; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1075; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1076; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1077; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1078; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1079; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1080; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1081; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1082; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1083; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1084; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1085; // @[Switch.scala 33:19:@5418.4]
  wire [47:0] _GEN_1086; // @[Switch.scala 33:19:@5418.4]
  wire [7:0] _T_24139; // @[Switch.scala 34:32:@5425.4]
  wire [15:0] _T_24147; // @[Switch.scala 34:32:@5433.4]
  wire [7:0] _T_24154; // @[Switch.scala 34:32:@5440.4]
  wire [31:0] _T_24163; // @[Switch.scala 34:32:@5449.4]
  wire [7:0] _T_24170; // @[Switch.scala 34:32:@5456.4]
  wire [15:0] _T_24178; // @[Switch.scala 34:32:@5464.4]
  wire [7:0] _T_24185; // @[Switch.scala 34:32:@5471.4]
  wire [31:0] _T_24194; // @[Switch.scala 34:32:@5480.4]
  wire [63:0] _T_24195; // @[Switch.scala 34:32:@5481.4]
  wire  _T_24199; // @[Switch.scala 30:53:@5484.4]
  wire  valid_17_0; // @[Switch.scala 30:36:@5485.4]
  wire  _T_24202; // @[Switch.scala 30:53:@5487.4]
  wire  valid_17_1; // @[Switch.scala 30:36:@5488.4]
  wire  _T_24205; // @[Switch.scala 30:53:@5490.4]
  wire  valid_17_2; // @[Switch.scala 30:36:@5491.4]
  wire  _T_24208; // @[Switch.scala 30:53:@5493.4]
  wire  valid_17_3; // @[Switch.scala 30:36:@5494.4]
  wire  _T_24211; // @[Switch.scala 30:53:@5496.4]
  wire  valid_17_4; // @[Switch.scala 30:36:@5497.4]
  wire  _T_24214; // @[Switch.scala 30:53:@5499.4]
  wire  valid_17_5; // @[Switch.scala 30:36:@5500.4]
  wire  _T_24217; // @[Switch.scala 30:53:@5502.4]
  wire  valid_17_6; // @[Switch.scala 30:36:@5503.4]
  wire  _T_24220; // @[Switch.scala 30:53:@5505.4]
  wire  valid_17_7; // @[Switch.scala 30:36:@5506.4]
  wire  _T_24223; // @[Switch.scala 30:53:@5508.4]
  wire  valid_17_8; // @[Switch.scala 30:36:@5509.4]
  wire  _T_24226; // @[Switch.scala 30:53:@5511.4]
  wire  valid_17_9; // @[Switch.scala 30:36:@5512.4]
  wire  _T_24229; // @[Switch.scala 30:53:@5514.4]
  wire  valid_17_10; // @[Switch.scala 30:36:@5515.4]
  wire  _T_24232; // @[Switch.scala 30:53:@5517.4]
  wire  valid_17_11; // @[Switch.scala 30:36:@5518.4]
  wire  _T_24235; // @[Switch.scala 30:53:@5520.4]
  wire  valid_17_12; // @[Switch.scala 30:36:@5521.4]
  wire  _T_24238; // @[Switch.scala 30:53:@5523.4]
  wire  valid_17_13; // @[Switch.scala 30:36:@5524.4]
  wire  _T_24241; // @[Switch.scala 30:53:@5526.4]
  wire  valid_17_14; // @[Switch.scala 30:36:@5527.4]
  wire  _T_24244; // @[Switch.scala 30:53:@5529.4]
  wire  valid_17_15; // @[Switch.scala 30:36:@5530.4]
  wire  _T_24247; // @[Switch.scala 30:53:@5532.4]
  wire  valid_17_16; // @[Switch.scala 30:36:@5533.4]
  wire  _T_24250; // @[Switch.scala 30:53:@5535.4]
  wire  valid_17_17; // @[Switch.scala 30:36:@5536.4]
  wire  _T_24253; // @[Switch.scala 30:53:@5538.4]
  wire  valid_17_18; // @[Switch.scala 30:36:@5539.4]
  wire  _T_24256; // @[Switch.scala 30:53:@5541.4]
  wire  valid_17_19; // @[Switch.scala 30:36:@5542.4]
  wire  _T_24259; // @[Switch.scala 30:53:@5544.4]
  wire  valid_17_20; // @[Switch.scala 30:36:@5545.4]
  wire  _T_24262; // @[Switch.scala 30:53:@5547.4]
  wire  valid_17_21; // @[Switch.scala 30:36:@5548.4]
  wire  _T_24265; // @[Switch.scala 30:53:@5550.4]
  wire  valid_17_22; // @[Switch.scala 30:36:@5551.4]
  wire  _T_24268; // @[Switch.scala 30:53:@5553.4]
  wire  valid_17_23; // @[Switch.scala 30:36:@5554.4]
  wire  _T_24271; // @[Switch.scala 30:53:@5556.4]
  wire  valid_17_24; // @[Switch.scala 30:36:@5557.4]
  wire  _T_24274; // @[Switch.scala 30:53:@5559.4]
  wire  valid_17_25; // @[Switch.scala 30:36:@5560.4]
  wire  _T_24277; // @[Switch.scala 30:53:@5562.4]
  wire  valid_17_26; // @[Switch.scala 30:36:@5563.4]
  wire  _T_24280; // @[Switch.scala 30:53:@5565.4]
  wire  valid_17_27; // @[Switch.scala 30:36:@5566.4]
  wire  _T_24283; // @[Switch.scala 30:53:@5568.4]
  wire  valid_17_28; // @[Switch.scala 30:36:@5569.4]
  wire  _T_24286; // @[Switch.scala 30:53:@5571.4]
  wire  valid_17_29; // @[Switch.scala 30:36:@5572.4]
  wire  _T_24289; // @[Switch.scala 30:53:@5574.4]
  wire  valid_17_30; // @[Switch.scala 30:36:@5575.4]
  wire  _T_24292; // @[Switch.scala 30:53:@5577.4]
  wire  valid_17_31; // @[Switch.scala 30:36:@5578.4]
  wire  _T_24295; // @[Switch.scala 30:53:@5580.4]
  wire  valid_17_32; // @[Switch.scala 30:36:@5581.4]
  wire  _T_24298; // @[Switch.scala 30:53:@5583.4]
  wire  valid_17_33; // @[Switch.scala 30:36:@5584.4]
  wire  _T_24301; // @[Switch.scala 30:53:@5586.4]
  wire  valid_17_34; // @[Switch.scala 30:36:@5587.4]
  wire  _T_24304; // @[Switch.scala 30:53:@5589.4]
  wire  valid_17_35; // @[Switch.scala 30:36:@5590.4]
  wire  _T_24307; // @[Switch.scala 30:53:@5592.4]
  wire  valid_17_36; // @[Switch.scala 30:36:@5593.4]
  wire  _T_24310; // @[Switch.scala 30:53:@5595.4]
  wire  valid_17_37; // @[Switch.scala 30:36:@5596.4]
  wire  _T_24313; // @[Switch.scala 30:53:@5598.4]
  wire  valid_17_38; // @[Switch.scala 30:36:@5599.4]
  wire  _T_24316; // @[Switch.scala 30:53:@5601.4]
  wire  valid_17_39; // @[Switch.scala 30:36:@5602.4]
  wire  _T_24319; // @[Switch.scala 30:53:@5604.4]
  wire  valid_17_40; // @[Switch.scala 30:36:@5605.4]
  wire  _T_24322; // @[Switch.scala 30:53:@5607.4]
  wire  valid_17_41; // @[Switch.scala 30:36:@5608.4]
  wire  _T_24325; // @[Switch.scala 30:53:@5610.4]
  wire  valid_17_42; // @[Switch.scala 30:36:@5611.4]
  wire  _T_24328; // @[Switch.scala 30:53:@5613.4]
  wire  valid_17_43; // @[Switch.scala 30:36:@5614.4]
  wire  _T_24331; // @[Switch.scala 30:53:@5616.4]
  wire  valid_17_44; // @[Switch.scala 30:36:@5617.4]
  wire  _T_24334; // @[Switch.scala 30:53:@5619.4]
  wire  valid_17_45; // @[Switch.scala 30:36:@5620.4]
  wire  _T_24337; // @[Switch.scala 30:53:@5622.4]
  wire  valid_17_46; // @[Switch.scala 30:36:@5623.4]
  wire  _T_24340; // @[Switch.scala 30:53:@5625.4]
  wire  valid_17_47; // @[Switch.scala 30:36:@5626.4]
  wire  _T_24343; // @[Switch.scala 30:53:@5628.4]
  wire  valid_17_48; // @[Switch.scala 30:36:@5629.4]
  wire  _T_24346; // @[Switch.scala 30:53:@5631.4]
  wire  valid_17_49; // @[Switch.scala 30:36:@5632.4]
  wire  _T_24349; // @[Switch.scala 30:53:@5634.4]
  wire  valid_17_50; // @[Switch.scala 30:36:@5635.4]
  wire  _T_24352; // @[Switch.scala 30:53:@5637.4]
  wire  valid_17_51; // @[Switch.scala 30:36:@5638.4]
  wire  _T_24355; // @[Switch.scala 30:53:@5640.4]
  wire  valid_17_52; // @[Switch.scala 30:36:@5641.4]
  wire  _T_24358; // @[Switch.scala 30:53:@5643.4]
  wire  valid_17_53; // @[Switch.scala 30:36:@5644.4]
  wire  _T_24361; // @[Switch.scala 30:53:@5646.4]
  wire  valid_17_54; // @[Switch.scala 30:36:@5647.4]
  wire  _T_24364; // @[Switch.scala 30:53:@5649.4]
  wire  valid_17_55; // @[Switch.scala 30:36:@5650.4]
  wire  _T_24367; // @[Switch.scala 30:53:@5652.4]
  wire  valid_17_56; // @[Switch.scala 30:36:@5653.4]
  wire  _T_24370; // @[Switch.scala 30:53:@5655.4]
  wire  valid_17_57; // @[Switch.scala 30:36:@5656.4]
  wire  _T_24373; // @[Switch.scala 30:53:@5658.4]
  wire  valid_17_58; // @[Switch.scala 30:36:@5659.4]
  wire  _T_24376; // @[Switch.scala 30:53:@5661.4]
  wire  valid_17_59; // @[Switch.scala 30:36:@5662.4]
  wire  _T_24379; // @[Switch.scala 30:53:@5664.4]
  wire  valid_17_60; // @[Switch.scala 30:36:@5665.4]
  wire  _T_24382; // @[Switch.scala 30:53:@5667.4]
  wire  valid_17_61; // @[Switch.scala 30:36:@5668.4]
  wire  _T_24385; // @[Switch.scala 30:53:@5670.4]
  wire  valid_17_62; // @[Switch.scala 30:36:@5671.4]
  wire  _T_24388; // @[Switch.scala 30:53:@5673.4]
  wire  valid_17_63; // @[Switch.scala 30:36:@5674.4]
  wire [5:0] _T_24454; // @[Mux.scala 31:69:@5676.4]
  wire [5:0] _T_24455; // @[Mux.scala 31:69:@5677.4]
  wire [5:0] _T_24456; // @[Mux.scala 31:69:@5678.4]
  wire [5:0] _T_24457; // @[Mux.scala 31:69:@5679.4]
  wire [5:0] _T_24458; // @[Mux.scala 31:69:@5680.4]
  wire [5:0] _T_24459; // @[Mux.scala 31:69:@5681.4]
  wire [5:0] _T_24460; // @[Mux.scala 31:69:@5682.4]
  wire [5:0] _T_24461; // @[Mux.scala 31:69:@5683.4]
  wire [5:0] _T_24462; // @[Mux.scala 31:69:@5684.4]
  wire [5:0] _T_24463; // @[Mux.scala 31:69:@5685.4]
  wire [5:0] _T_24464; // @[Mux.scala 31:69:@5686.4]
  wire [5:0] _T_24465; // @[Mux.scala 31:69:@5687.4]
  wire [5:0] _T_24466; // @[Mux.scala 31:69:@5688.4]
  wire [5:0] _T_24467; // @[Mux.scala 31:69:@5689.4]
  wire [5:0] _T_24468; // @[Mux.scala 31:69:@5690.4]
  wire [5:0] _T_24469; // @[Mux.scala 31:69:@5691.4]
  wire [5:0] _T_24470; // @[Mux.scala 31:69:@5692.4]
  wire [5:0] _T_24471; // @[Mux.scala 31:69:@5693.4]
  wire [5:0] _T_24472; // @[Mux.scala 31:69:@5694.4]
  wire [5:0] _T_24473; // @[Mux.scala 31:69:@5695.4]
  wire [5:0] _T_24474; // @[Mux.scala 31:69:@5696.4]
  wire [5:0] _T_24475; // @[Mux.scala 31:69:@5697.4]
  wire [5:0] _T_24476; // @[Mux.scala 31:69:@5698.4]
  wire [5:0] _T_24477; // @[Mux.scala 31:69:@5699.4]
  wire [5:0] _T_24478; // @[Mux.scala 31:69:@5700.4]
  wire [5:0] _T_24479; // @[Mux.scala 31:69:@5701.4]
  wire [5:0] _T_24480; // @[Mux.scala 31:69:@5702.4]
  wire [5:0] _T_24481; // @[Mux.scala 31:69:@5703.4]
  wire [5:0] _T_24482; // @[Mux.scala 31:69:@5704.4]
  wire [5:0] _T_24483; // @[Mux.scala 31:69:@5705.4]
  wire [5:0] _T_24484; // @[Mux.scala 31:69:@5706.4]
  wire [5:0] _T_24485; // @[Mux.scala 31:69:@5707.4]
  wire [5:0] _T_24486; // @[Mux.scala 31:69:@5708.4]
  wire [5:0] _T_24487; // @[Mux.scala 31:69:@5709.4]
  wire [5:0] _T_24488; // @[Mux.scala 31:69:@5710.4]
  wire [5:0] _T_24489; // @[Mux.scala 31:69:@5711.4]
  wire [5:0] _T_24490; // @[Mux.scala 31:69:@5712.4]
  wire [5:0] _T_24491; // @[Mux.scala 31:69:@5713.4]
  wire [5:0] _T_24492; // @[Mux.scala 31:69:@5714.4]
  wire [5:0] _T_24493; // @[Mux.scala 31:69:@5715.4]
  wire [5:0] _T_24494; // @[Mux.scala 31:69:@5716.4]
  wire [5:0] _T_24495; // @[Mux.scala 31:69:@5717.4]
  wire [5:0] _T_24496; // @[Mux.scala 31:69:@5718.4]
  wire [5:0] _T_24497; // @[Mux.scala 31:69:@5719.4]
  wire [5:0] _T_24498; // @[Mux.scala 31:69:@5720.4]
  wire [5:0] _T_24499; // @[Mux.scala 31:69:@5721.4]
  wire [5:0] _T_24500; // @[Mux.scala 31:69:@5722.4]
  wire [5:0] _T_24501; // @[Mux.scala 31:69:@5723.4]
  wire [5:0] _T_24502; // @[Mux.scala 31:69:@5724.4]
  wire [5:0] _T_24503; // @[Mux.scala 31:69:@5725.4]
  wire [5:0] _T_24504; // @[Mux.scala 31:69:@5726.4]
  wire [5:0] _T_24505; // @[Mux.scala 31:69:@5727.4]
  wire [5:0] _T_24506; // @[Mux.scala 31:69:@5728.4]
  wire [5:0] _T_24507; // @[Mux.scala 31:69:@5729.4]
  wire [5:0] _T_24508; // @[Mux.scala 31:69:@5730.4]
  wire [5:0] _T_24509; // @[Mux.scala 31:69:@5731.4]
  wire [5:0] _T_24510; // @[Mux.scala 31:69:@5732.4]
  wire [5:0] _T_24511; // @[Mux.scala 31:69:@5733.4]
  wire [5:0] _T_24512; // @[Mux.scala 31:69:@5734.4]
  wire [5:0] _T_24513; // @[Mux.scala 31:69:@5735.4]
  wire [5:0] _T_24514; // @[Mux.scala 31:69:@5736.4]
  wire [5:0] _T_24515; // @[Mux.scala 31:69:@5737.4]
  wire [5:0] select_17; // @[Mux.scala 31:69:@5738.4]
  wire [47:0] _GEN_1089; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1090; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1091; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1092; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1093; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1094; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1095; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1096; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1097; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1098; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1099; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1100; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1101; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1102; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1103; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1104; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1105; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1106; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1107; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1108; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1109; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1110; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1111; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1112; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1113; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1114; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1115; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1116; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1117; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1118; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1119; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1120; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1121; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1122; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1123; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1124; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1125; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1126; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1127; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1128; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1129; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1130; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1131; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1132; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1133; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1134; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1135; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1136; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1137; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1138; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1139; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1140; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1141; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1142; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1143; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1144; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1145; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1146; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1147; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1148; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1149; // @[Switch.scala 33:19:@5740.4]
  wire [47:0] _GEN_1150; // @[Switch.scala 33:19:@5740.4]
  wire [7:0] _T_24524; // @[Switch.scala 34:32:@5747.4]
  wire [15:0] _T_24532; // @[Switch.scala 34:32:@5755.4]
  wire [7:0] _T_24539; // @[Switch.scala 34:32:@5762.4]
  wire [31:0] _T_24548; // @[Switch.scala 34:32:@5771.4]
  wire [7:0] _T_24555; // @[Switch.scala 34:32:@5778.4]
  wire [15:0] _T_24563; // @[Switch.scala 34:32:@5786.4]
  wire [7:0] _T_24570; // @[Switch.scala 34:32:@5793.4]
  wire [31:0] _T_24579; // @[Switch.scala 34:32:@5802.4]
  wire [63:0] _T_24580; // @[Switch.scala 34:32:@5803.4]
  wire  _T_24584; // @[Switch.scala 30:53:@5806.4]
  wire  valid_18_0; // @[Switch.scala 30:36:@5807.4]
  wire  _T_24587; // @[Switch.scala 30:53:@5809.4]
  wire  valid_18_1; // @[Switch.scala 30:36:@5810.4]
  wire  _T_24590; // @[Switch.scala 30:53:@5812.4]
  wire  valid_18_2; // @[Switch.scala 30:36:@5813.4]
  wire  _T_24593; // @[Switch.scala 30:53:@5815.4]
  wire  valid_18_3; // @[Switch.scala 30:36:@5816.4]
  wire  _T_24596; // @[Switch.scala 30:53:@5818.4]
  wire  valid_18_4; // @[Switch.scala 30:36:@5819.4]
  wire  _T_24599; // @[Switch.scala 30:53:@5821.4]
  wire  valid_18_5; // @[Switch.scala 30:36:@5822.4]
  wire  _T_24602; // @[Switch.scala 30:53:@5824.4]
  wire  valid_18_6; // @[Switch.scala 30:36:@5825.4]
  wire  _T_24605; // @[Switch.scala 30:53:@5827.4]
  wire  valid_18_7; // @[Switch.scala 30:36:@5828.4]
  wire  _T_24608; // @[Switch.scala 30:53:@5830.4]
  wire  valid_18_8; // @[Switch.scala 30:36:@5831.4]
  wire  _T_24611; // @[Switch.scala 30:53:@5833.4]
  wire  valid_18_9; // @[Switch.scala 30:36:@5834.4]
  wire  _T_24614; // @[Switch.scala 30:53:@5836.4]
  wire  valid_18_10; // @[Switch.scala 30:36:@5837.4]
  wire  _T_24617; // @[Switch.scala 30:53:@5839.4]
  wire  valid_18_11; // @[Switch.scala 30:36:@5840.4]
  wire  _T_24620; // @[Switch.scala 30:53:@5842.4]
  wire  valid_18_12; // @[Switch.scala 30:36:@5843.4]
  wire  _T_24623; // @[Switch.scala 30:53:@5845.4]
  wire  valid_18_13; // @[Switch.scala 30:36:@5846.4]
  wire  _T_24626; // @[Switch.scala 30:53:@5848.4]
  wire  valid_18_14; // @[Switch.scala 30:36:@5849.4]
  wire  _T_24629; // @[Switch.scala 30:53:@5851.4]
  wire  valid_18_15; // @[Switch.scala 30:36:@5852.4]
  wire  _T_24632; // @[Switch.scala 30:53:@5854.4]
  wire  valid_18_16; // @[Switch.scala 30:36:@5855.4]
  wire  _T_24635; // @[Switch.scala 30:53:@5857.4]
  wire  valid_18_17; // @[Switch.scala 30:36:@5858.4]
  wire  _T_24638; // @[Switch.scala 30:53:@5860.4]
  wire  valid_18_18; // @[Switch.scala 30:36:@5861.4]
  wire  _T_24641; // @[Switch.scala 30:53:@5863.4]
  wire  valid_18_19; // @[Switch.scala 30:36:@5864.4]
  wire  _T_24644; // @[Switch.scala 30:53:@5866.4]
  wire  valid_18_20; // @[Switch.scala 30:36:@5867.4]
  wire  _T_24647; // @[Switch.scala 30:53:@5869.4]
  wire  valid_18_21; // @[Switch.scala 30:36:@5870.4]
  wire  _T_24650; // @[Switch.scala 30:53:@5872.4]
  wire  valid_18_22; // @[Switch.scala 30:36:@5873.4]
  wire  _T_24653; // @[Switch.scala 30:53:@5875.4]
  wire  valid_18_23; // @[Switch.scala 30:36:@5876.4]
  wire  _T_24656; // @[Switch.scala 30:53:@5878.4]
  wire  valid_18_24; // @[Switch.scala 30:36:@5879.4]
  wire  _T_24659; // @[Switch.scala 30:53:@5881.4]
  wire  valid_18_25; // @[Switch.scala 30:36:@5882.4]
  wire  _T_24662; // @[Switch.scala 30:53:@5884.4]
  wire  valid_18_26; // @[Switch.scala 30:36:@5885.4]
  wire  _T_24665; // @[Switch.scala 30:53:@5887.4]
  wire  valid_18_27; // @[Switch.scala 30:36:@5888.4]
  wire  _T_24668; // @[Switch.scala 30:53:@5890.4]
  wire  valid_18_28; // @[Switch.scala 30:36:@5891.4]
  wire  _T_24671; // @[Switch.scala 30:53:@5893.4]
  wire  valid_18_29; // @[Switch.scala 30:36:@5894.4]
  wire  _T_24674; // @[Switch.scala 30:53:@5896.4]
  wire  valid_18_30; // @[Switch.scala 30:36:@5897.4]
  wire  _T_24677; // @[Switch.scala 30:53:@5899.4]
  wire  valid_18_31; // @[Switch.scala 30:36:@5900.4]
  wire  _T_24680; // @[Switch.scala 30:53:@5902.4]
  wire  valid_18_32; // @[Switch.scala 30:36:@5903.4]
  wire  _T_24683; // @[Switch.scala 30:53:@5905.4]
  wire  valid_18_33; // @[Switch.scala 30:36:@5906.4]
  wire  _T_24686; // @[Switch.scala 30:53:@5908.4]
  wire  valid_18_34; // @[Switch.scala 30:36:@5909.4]
  wire  _T_24689; // @[Switch.scala 30:53:@5911.4]
  wire  valid_18_35; // @[Switch.scala 30:36:@5912.4]
  wire  _T_24692; // @[Switch.scala 30:53:@5914.4]
  wire  valid_18_36; // @[Switch.scala 30:36:@5915.4]
  wire  _T_24695; // @[Switch.scala 30:53:@5917.4]
  wire  valid_18_37; // @[Switch.scala 30:36:@5918.4]
  wire  _T_24698; // @[Switch.scala 30:53:@5920.4]
  wire  valid_18_38; // @[Switch.scala 30:36:@5921.4]
  wire  _T_24701; // @[Switch.scala 30:53:@5923.4]
  wire  valid_18_39; // @[Switch.scala 30:36:@5924.4]
  wire  _T_24704; // @[Switch.scala 30:53:@5926.4]
  wire  valid_18_40; // @[Switch.scala 30:36:@5927.4]
  wire  _T_24707; // @[Switch.scala 30:53:@5929.4]
  wire  valid_18_41; // @[Switch.scala 30:36:@5930.4]
  wire  _T_24710; // @[Switch.scala 30:53:@5932.4]
  wire  valid_18_42; // @[Switch.scala 30:36:@5933.4]
  wire  _T_24713; // @[Switch.scala 30:53:@5935.4]
  wire  valid_18_43; // @[Switch.scala 30:36:@5936.4]
  wire  _T_24716; // @[Switch.scala 30:53:@5938.4]
  wire  valid_18_44; // @[Switch.scala 30:36:@5939.4]
  wire  _T_24719; // @[Switch.scala 30:53:@5941.4]
  wire  valid_18_45; // @[Switch.scala 30:36:@5942.4]
  wire  _T_24722; // @[Switch.scala 30:53:@5944.4]
  wire  valid_18_46; // @[Switch.scala 30:36:@5945.4]
  wire  _T_24725; // @[Switch.scala 30:53:@5947.4]
  wire  valid_18_47; // @[Switch.scala 30:36:@5948.4]
  wire  _T_24728; // @[Switch.scala 30:53:@5950.4]
  wire  valid_18_48; // @[Switch.scala 30:36:@5951.4]
  wire  _T_24731; // @[Switch.scala 30:53:@5953.4]
  wire  valid_18_49; // @[Switch.scala 30:36:@5954.4]
  wire  _T_24734; // @[Switch.scala 30:53:@5956.4]
  wire  valid_18_50; // @[Switch.scala 30:36:@5957.4]
  wire  _T_24737; // @[Switch.scala 30:53:@5959.4]
  wire  valid_18_51; // @[Switch.scala 30:36:@5960.4]
  wire  _T_24740; // @[Switch.scala 30:53:@5962.4]
  wire  valid_18_52; // @[Switch.scala 30:36:@5963.4]
  wire  _T_24743; // @[Switch.scala 30:53:@5965.4]
  wire  valid_18_53; // @[Switch.scala 30:36:@5966.4]
  wire  _T_24746; // @[Switch.scala 30:53:@5968.4]
  wire  valid_18_54; // @[Switch.scala 30:36:@5969.4]
  wire  _T_24749; // @[Switch.scala 30:53:@5971.4]
  wire  valid_18_55; // @[Switch.scala 30:36:@5972.4]
  wire  _T_24752; // @[Switch.scala 30:53:@5974.4]
  wire  valid_18_56; // @[Switch.scala 30:36:@5975.4]
  wire  _T_24755; // @[Switch.scala 30:53:@5977.4]
  wire  valid_18_57; // @[Switch.scala 30:36:@5978.4]
  wire  _T_24758; // @[Switch.scala 30:53:@5980.4]
  wire  valid_18_58; // @[Switch.scala 30:36:@5981.4]
  wire  _T_24761; // @[Switch.scala 30:53:@5983.4]
  wire  valid_18_59; // @[Switch.scala 30:36:@5984.4]
  wire  _T_24764; // @[Switch.scala 30:53:@5986.4]
  wire  valid_18_60; // @[Switch.scala 30:36:@5987.4]
  wire  _T_24767; // @[Switch.scala 30:53:@5989.4]
  wire  valid_18_61; // @[Switch.scala 30:36:@5990.4]
  wire  _T_24770; // @[Switch.scala 30:53:@5992.4]
  wire  valid_18_62; // @[Switch.scala 30:36:@5993.4]
  wire  _T_24773; // @[Switch.scala 30:53:@5995.4]
  wire  valid_18_63; // @[Switch.scala 30:36:@5996.4]
  wire [5:0] _T_24839; // @[Mux.scala 31:69:@5998.4]
  wire [5:0] _T_24840; // @[Mux.scala 31:69:@5999.4]
  wire [5:0] _T_24841; // @[Mux.scala 31:69:@6000.4]
  wire [5:0] _T_24842; // @[Mux.scala 31:69:@6001.4]
  wire [5:0] _T_24843; // @[Mux.scala 31:69:@6002.4]
  wire [5:0] _T_24844; // @[Mux.scala 31:69:@6003.4]
  wire [5:0] _T_24845; // @[Mux.scala 31:69:@6004.4]
  wire [5:0] _T_24846; // @[Mux.scala 31:69:@6005.4]
  wire [5:0] _T_24847; // @[Mux.scala 31:69:@6006.4]
  wire [5:0] _T_24848; // @[Mux.scala 31:69:@6007.4]
  wire [5:0] _T_24849; // @[Mux.scala 31:69:@6008.4]
  wire [5:0] _T_24850; // @[Mux.scala 31:69:@6009.4]
  wire [5:0] _T_24851; // @[Mux.scala 31:69:@6010.4]
  wire [5:0] _T_24852; // @[Mux.scala 31:69:@6011.4]
  wire [5:0] _T_24853; // @[Mux.scala 31:69:@6012.4]
  wire [5:0] _T_24854; // @[Mux.scala 31:69:@6013.4]
  wire [5:0] _T_24855; // @[Mux.scala 31:69:@6014.4]
  wire [5:0] _T_24856; // @[Mux.scala 31:69:@6015.4]
  wire [5:0] _T_24857; // @[Mux.scala 31:69:@6016.4]
  wire [5:0] _T_24858; // @[Mux.scala 31:69:@6017.4]
  wire [5:0] _T_24859; // @[Mux.scala 31:69:@6018.4]
  wire [5:0] _T_24860; // @[Mux.scala 31:69:@6019.4]
  wire [5:0] _T_24861; // @[Mux.scala 31:69:@6020.4]
  wire [5:0] _T_24862; // @[Mux.scala 31:69:@6021.4]
  wire [5:0] _T_24863; // @[Mux.scala 31:69:@6022.4]
  wire [5:0] _T_24864; // @[Mux.scala 31:69:@6023.4]
  wire [5:0] _T_24865; // @[Mux.scala 31:69:@6024.4]
  wire [5:0] _T_24866; // @[Mux.scala 31:69:@6025.4]
  wire [5:0] _T_24867; // @[Mux.scala 31:69:@6026.4]
  wire [5:0] _T_24868; // @[Mux.scala 31:69:@6027.4]
  wire [5:0] _T_24869; // @[Mux.scala 31:69:@6028.4]
  wire [5:0] _T_24870; // @[Mux.scala 31:69:@6029.4]
  wire [5:0] _T_24871; // @[Mux.scala 31:69:@6030.4]
  wire [5:0] _T_24872; // @[Mux.scala 31:69:@6031.4]
  wire [5:0] _T_24873; // @[Mux.scala 31:69:@6032.4]
  wire [5:0] _T_24874; // @[Mux.scala 31:69:@6033.4]
  wire [5:0] _T_24875; // @[Mux.scala 31:69:@6034.4]
  wire [5:0] _T_24876; // @[Mux.scala 31:69:@6035.4]
  wire [5:0] _T_24877; // @[Mux.scala 31:69:@6036.4]
  wire [5:0] _T_24878; // @[Mux.scala 31:69:@6037.4]
  wire [5:0] _T_24879; // @[Mux.scala 31:69:@6038.4]
  wire [5:0] _T_24880; // @[Mux.scala 31:69:@6039.4]
  wire [5:0] _T_24881; // @[Mux.scala 31:69:@6040.4]
  wire [5:0] _T_24882; // @[Mux.scala 31:69:@6041.4]
  wire [5:0] _T_24883; // @[Mux.scala 31:69:@6042.4]
  wire [5:0] _T_24884; // @[Mux.scala 31:69:@6043.4]
  wire [5:0] _T_24885; // @[Mux.scala 31:69:@6044.4]
  wire [5:0] _T_24886; // @[Mux.scala 31:69:@6045.4]
  wire [5:0] _T_24887; // @[Mux.scala 31:69:@6046.4]
  wire [5:0] _T_24888; // @[Mux.scala 31:69:@6047.4]
  wire [5:0] _T_24889; // @[Mux.scala 31:69:@6048.4]
  wire [5:0] _T_24890; // @[Mux.scala 31:69:@6049.4]
  wire [5:0] _T_24891; // @[Mux.scala 31:69:@6050.4]
  wire [5:0] _T_24892; // @[Mux.scala 31:69:@6051.4]
  wire [5:0] _T_24893; // @[Mux.scala 31:69:@6052.4]
  wire [5:0] _T_24894; // @[Mux.scala 31:69:@6053.4]
  wire [5:0] _T_24895; // @[Mux.scala 31:69:@6054.4]
  wire [5:0] _T_24896; // @[Mux.scala 31:69:@6055.4]
  wire [5:0] _T_24897; // @[Mux.scala 31:69:@6056.4]
  wire [5:0] _T_24898; // @[Mux.scala 31:69:@6057.4]
  wire [5:0] _T_24899; // @[Mux.scala 31:69:@6058.4]
  wire [5:0] _T_24900; // @[Mux.scala 31:69:@6059.4]
  wire [5:0] select_18; // @[Mux.scala 31:69:@6060.4]
  wire [47:0] _GEN_1153; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1154; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1155; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1156; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1157; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1158; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1159; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1160; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1161; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1162; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1163; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1164; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1165; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1166; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1167; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1168; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1169; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1170; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1171; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1172; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1173; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1174; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1175; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1176; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1177; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1178; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1179; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1180; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1181; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1182; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1183; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1184; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1185; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1186; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1187; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1188; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1189; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1190; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1191; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1192; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1193; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1194; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1195; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1196; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1197; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1198; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1199; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1200; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1201; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1202; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1203; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1204; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1205; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1206; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1207; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1208; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1209; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1210; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1211; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1212; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1213; // @[Switch.scala 33:19:@6062.4]
  wire [47:0] _GEN_1214; // @[Switch.scala 33:19:@6062.4]
  wire [7:0] _T_24909; // @[Switch.scala 34:32:@6069.4]
  wire [15:0] _T_24917; // @[Switch.scala 34:32:@6077.4]
  wire [7:0] _T_24924; // @[Switch.scala 34:32:@6084.4]
  wire [31:0] _T_24933; // @[Switch.scala 34:32:@6093.4]
  wire [7:0] _T_24940; // @[Switch.scala 34:32:@6100.4]
  wire [15:0] _T_24948; // @[Switch.scala 34:32:@6108.4]
  wire [7:0] _T_24955; // @[Switch.scala 34:32:@6115.4]
  wire [31:0] _T_24964; // @[Switch.scala 34:32:@6124.4]
  wire [63:0] _T_24965; // @[Switch.scala 34:32:@6125.4]
  wire  _T_24969; // @[Switch.scala 30:53:@6128.4]
  wire  valid_19_0; // @[Switch.scala 30:36:@6129.4]
  wire  _T_24972; // @[Switch.scala 30:53:@6131.4]
  wire  valid_19_1; // @[Switch.scala 30:36:@6132.4]
  wire  _T_24975; // @[Switch.scala 30:53:@6134.4]
  wire  valid_19_2; // @[Switch.scala 30:36:@6135.4]
  wire  _T_24978; // @[Switch.scala 30:53:@6137.4]
  wire  valid_19_3; // @[Switch.scala 30:36:@6138.4]
  wire  _T_24981; // @[Switch.scala 30:53:@6140.4]
  wire  valid_19_4; // @[Switch.scala 30:36:@6141.4]
  wire  _T_24984; // @[Switch.scala 30:53:@6143.4]
  wire  valid_19_5; // @[Switch.scala 30:36:@6144.4]
  wire  _T_24987; // @[Switch.scala 30:53:@6146.4]
  wire  valid_19_6; // @[Switch.scala 30:36:@6147.4]
  wire  _T_24990; // @[Switch.scala 30:53:@6149.4]
  wire  valid_19_7; // @[Switch.scala 30:36:@6150.4]
  wire  _T_24993; // @[Switch.scala 30:53:@6152.4]
  wire  valid_19_8; // @[Switch.scala 30:36:@6153.4]
  wire  _T_24996; // @[Switch.scala 30:53:@6155.4]
  wire  valid_19_9; // @[Switch.scala 30:36:@6156.4]
  wire  _T_24999; // @[Switch.scala 30:53:@6158.4]
  wire  valid_19_10; // @[Switch.scala 30:36:@6159.4]
  wire  _T_25002; // @[Switch.scala 30:53:@6161.4]
  wire  valid_19_11; // @[Switch.scala 30:36:@6162.4]
  wire  _T_25005; // @[Switch.scala 30:53:@6164.4]
  wire  valid_19_12; // @[Switch.scala 30:36:@6165.4]
  wire  _T_25008; // @[Switch.scala 30:53:@6167.4]
  wire  valid_19_13; // @[Switch.scala 30:36:@6168.4]
  wire  _T_25011; // @[Switch.scala 30:53:@6170.4]
  wire  valid_19_14; // @[Switch.scala 30:36:@6171.4]
  wire  _T_25014; // @[Switch.scala 30:53:@6173.4]
  wire  valid_19_15; // @[Switch.scala 30:36:@6174.4]
  wire  _T_25017; // @[Switch.scala 30:53:@6176.4]
  wire  valid_19_16; // @[Switch.scala 30:36:@6177.4]
  wire  _T_25020; // @[Switch.scala 30:53:@6179.4]
  wire  valid_19_17; // @[Switch.scala 30:36:@6180.4]
  wire  _T_25023; // @[Switch.scala 30:53:@6182.4]
  wire  valid_19_18; // @[Switch.scala 30:36:@6183.4]
  wire  _T_25026; // @[Switch.scala 30:53:@6185.4]
  wire  valid_19_19; // @[Switch.scala 30:36:@6186.4]
  wire  _T_25029; // @[Switch.scala 30:53:@6188.4]
  wire  valid_19_20; // @[Switch.scala 30:36:@6189.4]
  wire  _T_25032; // @[Switch.scala 30:53:@6191.4]
  wire  valid_19_21; // @[Switch.scala 30:36:@6192.4]
  wire  _T_25035; // @[Switch.scala 30:53:@6194.4]
  wire  valid_19_22; // @[Switch.scala 30:36:@6195.4]
  wire  _T_25038; // @[Switch.scala 30:53:@6197.4]
  wire  valid_19_23; // @[Switch.scala 30:36:@6198.4]
  wire  _T_25041; // @[Switch.scala 30:53:@6200.4]
  wire  valid_19_24; // @[Switch.scala 30:36:@6201.4]
  wire  _T_25044; // @[Switch.scala 30:53:@6203.4]
  wire  valid_19_25; // @[Switch.scala 30:36:@6204.4]
  wire  _T_25047; // @[Switch.scala 30:53:@6206.4]
  wire  valid_19_26; // @[Switch.scala 30:36:@6207.4]
  wire  _T_25050; // @[Switch.scala 30:53:@6209.4]
  wire  valid_19_27; // @[Switch.scala 30:36:@6210.4]
  wire  _T_25053; // @[Switch.scala 30:53:@6212.4]
  wire  valid_19_28; // @[Switch.scala 30:36:@6213.4]
  wire  _T_25056; // @[Switch.scala 30:53:@6215.4]
  wire  valid_19_29; // @[Switch.scala 30:36:@6216.4]
  wire  _T_25059; // @[Switch.scala 30:53:@6218.4]
  wire  valid_19_30; // @[Switch.scala 30:36:@6219.4]
  wire  _T_25062; // @[Switch.scala 30:53:@6221.4]
  wire  valid_19_31; // @[Switch.scala 30:36:@6222.4]
  wire  _T_25065; // @[Switch.scala 30:53:@6224.4]
  wire  valid_19_32; // @[Switch.scala 30:36:@6225.4]
  wire  _T_25068; // @[Switch.scala 30:53:@6227.4]
  wire  valid_19_33; // @[Switch.scala 30:36:@6228.4]
  wire  _T_25071; // @[Switch.scala 30:53:@6230.4]
  wire  valid_19_34; // @[Switch.scala 30:36:@6231.4]
  wire  _T_25074; // @[Switch.scala 30:53:@6233.4]
  wire  valid_19_35; // @[Switch.scala 30:36:@6234.4]
  wire  _T_25077; // @[Switch.scala 30:53:@6236.4]
  wire  valid_19_36; // @[Switch.scala 30:36:@6237.4]
  wire  _T_25080; // @[Switch.scala 30:53:@6239.4]
  wire  valid_19_37; // @[Switch.scala 30:36:@6240.4]
  wire  _T_25083; // @[Switch.scala 30:53:@6242.4]
  wire  valid_19_38; // @[Switch.scala 30:36:@6243.4]
  wire  _T_25086; // @[Switch.scala 30:53:@6245.4]
  wire  valid_19_39; // @[Switch.scala 30:36:@6246.4]
  wire  _T_25089; // @[Switch.scala 30:53:@6248.4]
  wire  valid_19_40; // @[Switch.scala 30:36:@6249.4]
  wire  _T_25092; // @[Switch.scala 30:53:@6251.4]
  wire  valid_19_41; // @[Switch.scala 30:36:@6252.4]
  wire  _T_25095; // @[Switch.scala 30:53:@6254.4]
  wire  valid_19_42; // @[Switch.scala 30:36:@6255.4]
  wire  _T_25098; // @[Switch.scala 30:53:@6257.4]
  wire  valid_19_43; // @[Switch.scala 30:36:@6258.4]
  wire  _T_25101; // @[Switch.scala 30:53:@6260.4]
  wire  valid_19_44; // @[Switch.scala 30:36:@6261.4]
  wire  _T_25104; // @[Switch.scala 30:53:@6263.4]
  wire  valid_19_45; // @[Switch.scala 30:36:@6264.4]
  wire  _T_25107; // @[Switch.scala 30:53:@6266.4]
  wire  valid_19_46; // @[Switch.scala 30:36:@6267.4]
  wire  _T_25110; // @[Switch.scala 30:53:@6269.4]
  wire  valid_19_47; // @[Switch.scala 30:36:@6270.4]
  wire  _T_25113; // @[Switch.scala 30:53:@6272.4]
  wire  valid_19_48; // @[Switch.scala 30:36:@6273.4]
  wire  _T_25116; // @[Switch.scala 30:53:@6275.4]
  wire  valid_19_49; // @[Switch.scala 30:36:@6276.4]
  wire  _T_25119; // @[Switch.scala 30:53:@6278.4]
  wire  valid_19_50; // @[Switch.scala 30:36:@6279.4]
  wire  _T_25122; // @[Switch.scala 30:53:@6281.4]
  wire  valid_19_51; // @[Switch.scala 30:36:@6282.4]
  wire  _T_25125; // @[Switch.scala 30:53:@6284.4]
  wire  valid_19_52; // @[Switch.scala 30:36:@6285.4]
  wire  _T_25128; // @[Switch.scala 30:53:@6287.4]
  wire  valid_19_53; // @[Switch.scala 30:36:@6288.4]
  wire  _T_25131; // @[Switch.scala 30:53:@6290.4]
  wire  valid_19_54; // @[Switch.scala 30:36:@6291.4]
  wire  _T_25134; // @[Switch.scala 30:53:@6293.4]
  wire  valid_19_55; // @[Switch.scala 30:36:@6294.4]
  wire  _T_25137; // @[Switch.scala 30:53:@6296.4]
  wire  valid_19_56; // @[Switch.scala 30:36:@6297.4]
  wire  _T_25140; // @[Switch.scala 30:53:@6299.4]
  wire  valid_19_57; // @[Switch.scala 30:36:@6300.4]
  wire  _T_25143; // @[Switch.scala 30:53:@6302.4]
  wire  valid_19_58; // @[Switch.scala 30:36:@6303.4]
  wire  _T_25146; // @[Switch.scala 30:53:@6305.4]
  wire  valid_19_59; // @[Switch.scala 30:36:@6306.4]
  wire  _T_25149; // @[Switch.scala 30:53:@6308.4]
  wire  valid_19_60; // @[Switch.scala 30:36:@6309.4]
  wire  _T_25152; // @[Switch.scala 30:53:@6311.4]
  wire  valid_19_61; // @[Switch.scala 30:36:@6312.4]
  wire  _T_25155; // @[Switch.scala 30:53:@6314.4]
  wire  valid_19_62; // @[Switch.scala 30:36:@6315.4]
  wire  _T_25158; // @[Switch.scala 30:53:@6317.4]
  wire  valid_19_63; // @[Switch.scala 30:36:@6318.4]
  wire [5:0] _T_25224; // @[Mux.scala 31:69:@6320.4]
  wire [5:0] _T_25225; // @[Mux.scala 31:69:@6321.4]
  wire [5:0] _T_25226; // @[Mux.scala 31:69:@6322.4]
  wire [5:0] _T_25227; // @[Mux.scala 31:69:@6323.4]
  wire [5:0] _T_25228; // @[Mux.scala 31:69:@6324.4]
  wire [5:0] _T_25229; // @[Mux.scala 31:69:@6325.4]
  wire [5:0] _T_25230; // @[Mux.scala 31:69:@6326.4]
  wire [5:0] _T_25231; // @[Mux.scala 31:69:@6327.4]
  wire [5:0] _T_25232; // @[Mux.scala 31:69:@6328.4]
  wire [5:0] _T_25233; // @[Mux.scala 31:69:@6329.4]
  wire [5:0] _T_25234; // @[Mux.scala 31:69:@6330.4]
  wire [5:0] _T_25235; // @[Mux.scala 31:69:@6331.4]
  wire [5:0] _T_25236; // @[Mux.scala 31:69:@6332.4]
  wire [5:0] _T_25237; // @[Mux.scala 31:69:@6333.4]
  wire [5:0] _T_25238; // @[Mux.scala 31:69:@6334.4]
  wire [5:0] _T_25239; // @[Mux.scala 31:69:@6335.4]
  wire [5:0] _T_25240; // @[Mux.scala 31:69:@6336.4]
  wire [5:0] _T_25241; // @[Mux.scala 31:69:@6337.4]
  wire [5:0] _T_25242; // @[Mux.scala 31:69:@6338.4]
  wire [5:0] _T_25243; // @[Mux.scala 31:69:@6339.4]
  wire [5:0] _T_25244; // @[Mux.scala 31:69:@6340.4]
  wire [5:0] _T_25245; // @[Mux.scala 31:69:@6341.4]
  wire [5:0] _T_25246; // @[Mux.scala 31:69:@6342.4]
  wire [5:0] _T_25247; // @[Mux.scala 31:69:@6343.4]
  wire [5:0] _T_25248; // @[Mux.scala 31:69:@6344.4]
  wire [5:0] _T_25249; // @[Mux.scala 31:69:@6345.4]
  wire [5:0] _T_25250; // @[Mux.scala 31:69:@6346.4]
  wire [5:0] _T_25251; // @[Mux.scala 31:69:@6347.4]
  wire [5:0] _T_25252; // @[Mux.scala 31:69:@6348.4]
  wire [5:0] _T_25253; // @[Mux.scala 31:69:@6349.4]
  wire [5:0] _T_25254; // @[Mux.scala 31:69:@6350.4]
  wire [5:0] _T_25255; // @[Mux.scala 31:69:@6351.4]
  wire [5:0] _T_25256; // @[Mux.scala 31:69:@6352.4]
  wire [5:0] _T_25257; // @[Mux.scala 31:69:@6353.4]
  wire [5:0] _T_25258; // @[Mux.scala 31:69:@6354.4]
  wire [5:0] _T_25259; // @[Mux.scala 31:69:@6355.4]
  wire [5:0] _T_25260; // @[Mux.scala 31:69:@6356.4]
  wire [5:0] _T_25261; // @[Mux.scala 31:69:@6357.4]
  wire [5:0] _T_25262; // @[Mux.scala 31:69:@6358.4]
  wire [5:0] _T_25263; // @[Mux.scala 31:69:@6359.4]
  wire [5:0] _T_25264; // @[Mux.scala 31:69:@6360.4]
  wire [5:0] _T_25265; // @[Mux.scala 31:69:@6361.4]
  wire [5:0] _T_25266; // @[Mux.scala 31:69:@6362.4]
  wire [5:0] _T_25267; // @[Mux.scala 31:69:@6363.4]
  wire [5:0] _T_25268; // @[Mux.scala 31:69:@6364.4]
  wire [5:0] _T_25269; // @[Mux.scala 31:69:@6365.4]
  wire [5:0] _T_25270; // @[Mux.scala 31:69:@6366.4]
  wire [5:0] _T_25271; // @[Mux.scala 31:69:@6367.4]
  wire [5:0] _T_25272; // @[Mux.scala 31:69:@6368.4]
  wire [5:0] _T_25273; // @[Mux.scala 31:69:@6369.4]
  wire [5:0] _T_25274; // @[Mux.scala 31:69:@6370.4]
  wire [5:0] _T_25275; // @[Mux.scala 31:69:@6371.4]
  wire [5:0] _T_25276; // @[Mux.scala 31:69:@6372.4]
  wire [5:0] _T_25277; // @[Mux.scala 31:69:@6373.4]
  wire [5:0] _T_25278; // @[Mux.scala 31:69:@6374.4]
  wire [5:0] _T_25279; // @[Mux.scala 31:69:@6375.4]
  wire [5:0] _T_25280; // @[Mux.scala 31:69:@6376.4]
  wire [5:0] _T_25281; // @[Mux.scala 31:69:@6377.4]
  wire [5:0] _T_25282; // @[Mux.scala 31:69:@6378.4]
  wire [5:0] _T_25283; // @[Mux.scala 31:69:@6379.4]
  wire [5:0] _T_25284; // @[Mux.scala 31:69:@6380.4]
  wire [5:0] _T_25285; // @[Mux.scala 31:69:@6381.4]
  wire [5:0] select_19; // @[Mux.scala 31:69:@6382.4]
  wire [47:0] _GEN_1217; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1218; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1219; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1220; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1221; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1222; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1223; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1224; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1225; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1226; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1227; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1228; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1229; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1230; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1231; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1232; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1233; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1234; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1235; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1236; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1237; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1238; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1239; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1240; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1241; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1242; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1243; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1244; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1245; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1246; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1247; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1248; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1249; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1250; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1251; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1252; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1253; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1254; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1255; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1256; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1257; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1258; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1259; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1260; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1261; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1262; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1263; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1264; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1265; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1266; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1267; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1268; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1269; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1270; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1271; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1272; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1273; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1274; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1275; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1276; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1277; // @[Switch.scala 33:19:@6384.4]
  wire [47:0] _GEN_1278; // @[Switch.scala 33:19:@6384.4]
  wire [7:0] _T_25294; // @[Switch.scala 34:32:@6391.4]
  wire [15:0] _T_25302; // @[Switch.scala 34:32:@6399.4]
  wire [7:0] _T_25309; // @[Switch.scala 34:32:@6406.4]
  wire [31:0] _T_25318; // @[Switch.scala 34:32:@6415.4]
  wire [7:0] _T_25325; // @[Switch.scala 34:32:@6422.4]
  wire [15:0] _T_25333; // @[Switch.scala 34:32:@6430.4]
  wire [7:0] _T_25340; // @[Switch.scala 34:32:@6437.4]
  wire [31:0] _T_25349; // @[Switch.scala 34:32:@6446.4]
  wire [63:0] _T_25350; // @[Switch.scala 34:32:@6447.4]
  wire  _T_25354; // @[Switch.scala 30:53:@6450.4]
  wire  valid_20_0; // @[Switch.scala 30:36:@6451.4]
  wire  _T_25357; // @[Switch.scala 30:53:@6453.4]
  wire  valid_20_1; // @[Switch.scala 30:36:@6454.4]
  wire  _T_25360; // @[Switch.scala 30:53:@6456.4]
  wire  valid_20_2; // @[Switch.scala 30:36:@6457.4]
  wire  _T_25363; // @[Switch.scala 30:53:@6459.4]
  wire  valid_20_3; // @[Switch.scala 30:36:@6460.4]
  wire  _T_25366; // @[Switch.scala 30:53:@6462.4]
  wire  valid_20_4; // @[Switch.scala 30:36:@6463.4]
  wire  _T_25369; // @[Switch.scala 30:53:@6465.4]
  wire  valid_20_5; // @[Switch.scala 30:36:@6466.4]
  wire  _T_25372; // @[Switch.scala 30:53:@6468.4]
  wire  valid_20_6; // @[Switch.scala 30:36:@6469.4]
  wire  _T_25375; // @[Switch.scala 30:53:@6471.4]
  wire  valid_20_7; // @[Switch.scala 30:36:@6472.4]
  wire  _T_25378; // @[Switch.scala 30:53:@6474.4]
  wire  valid_20_8; // @[Switch.scala 30:36:@6475.4]
  wire  _T_25381; // @[Switch.scala 30:53:@6477.4]
  wire  valid_20_9; // @[Switch.scala 30:36:@6478.4]
  wire  _T_25384; // @[Switch.scala 30:53:@6480.4]
  wire  valid_20_10; // @[Switch.scala 30:36:@6481.4]
  wire  _T_25387; // @[Switch.scala 30:53:@6483.4]
  wire  valid_20_11; // @[Switch.scala 30:36:@6484.4]
  wire  _T_25390; // @[Switch.scala 30:53:@6486.4]
  wire  valid_20_12; // @[Switch.scala 30:36:@6487.4]
  wire  _T_25393; // @[Switch.scala 30:53:@6489.4]
  wire  valid_20_13; // @[Switch.scala 30:36:@6490.4]
  wire  _T_25396; // @[Switch.scala 30:53:@6492.4]
  wire  valid_20_14; // @[Switch.scala 30:36:@6493.4]
  wire  _T_25399; // @[Switch.scala 30:53:@6495.4]
  wire  valid_20_15; // @[Switch.scala 30:36:@6496.4]
  wire  _T_25402; // @[Switch.scala 30:53:@6498.4]
  wire  valid_20_16; // @[Switch.scala 30:36:@6499.4]
  wire  _T_25405; // @[Switch.scala 30:53:@6501.4]
  wire  valid_20_17; // @[Switch.scala 30:36:@6502.4]
  wire  _T_25408; // @[Switch.scala 30:53:@6504.4]
  wire  valid_20_18; // @[Switch.scala 30:36:@6505.4]
  wire  _T_25411; // @[Switch.scala 30:53:@6507.4]
  wire  valid_20_19; // @[Switch.scala 30:36:@6508.4]
  wire  _T_25414; // @[Switch.scala 30:53:@6510.4]
  wire  valid_20_20; // @[Switch.scala 30:36:@6511.4]
  wire  _T_25417; // @[Switch.scala 30:53:@6513.4]
  wire  valid_20_21; // @[Switch.scala 30:36:@6514.4]
  wire  _T_25420; // @[Switch.scala 30:53:@6516.4]
  wire  valid_20_22; // @[Switch.scala 30:36:@6517.4]
  wire  _T_25423; // @[Switch.scala 30:53:@6519.4]
  wire  valid_20_23; // @[Switch.scala 30:36:@6520.4]
  wire  _T_25426; // @[Switch.scala 30:53:@6522.4]
  wire  valid_20_24; // @[Switch.scala 30:36:@6523.4]
  wire  _T_25429; // @[Switch.scala 30:53:@6525.4]
  wire  valid_20_25; // @[Switch.scala 30:36:@6526.4]
  wire  _T_25432; // @[Switch.scala 30:53:@6528.4]
  wire  valid_20_26; // @[Switch.scala 30:36:@6529.4]
  wire  _T_25435; // @[Switch.scala 30:53:@6531.4]
  wire  valid_20_27; // @[Switch.scala 30:36:@6532.4]
  wire  _T_25438; // @[Switch.scala 30:53:@6534.4]
  wire  valid_20_28; // @[Switch.scala 30:36:@6535.4]
  wire  _T_25441; // @[Switch.scala 30:53:@6537.4]
  wire  valid_20_29; // @[Switch.scala 30:36:@6538.4]
  wire  _T_25444; // @[Switch.scala 30:53:@6540.4]
  wire  valid_20_30; // @[Switch.scala 30:36:@6541.4]
  wire  _T_25447; // @[Switch.scala 30:53:@6543.4]
  wire  valid_20_31; // @[Switch.scala 30:36:@6544.4]
  wire  _T_25450; // @[Switch.scala 30:53:@6546.4]
  wire  valid_20_32; // @[Switch.scala 30:36:@6547.4]
  wire  _T_25453; // @[Switch.scala 30:53:@6549.4]
  wire  valid_20_33; // @[Switch.scala 30:36:@6550.4]
  wire  _T_25456; // @[Switch.scala 30:53:@6552.4]
  wire  valid_20_34; // @[Switch.scala 30:36:@6553.4]
  wire  _T_25459; // @[Switch.scala 30:53:@6555.4]
  wire  valid_20_35; // @[Switch.scala 30:36:@6556.4]
  wire  _T_25462; // @[Switch.scala 30:53:@6558.4]
  wire  valid_20_36; // @[Switch.scala 30:36:@6559.4]
  wire  _T_25465; // @[Switch.scala 30:53:@6561.4]
  wire  valid_20_37; // @[Switch.scala 30:36:@6562.4]
  wire  _T_25468; // @[Switch.scala 30:53:@6564.4]
  wire  valid_20_38; // @[Switch.scala 30:36:@6565.4]
  wire  _T_25471; // @[Switch.scala 30:53:@6567.4]
  wire  valid_20_39; // @[Switch.scala 30:36:@6568.4]
  wire  _T_25474; // @[Switch.scala 30:53:@6570.4]
  wire  valid_20_40; // @[Switch.scala 30:36:@6571.4]
  wire  _T_25477; // @[Switch.scala 30:53:@6573.4]
  wire  valid_20_41; // @[Switch.scala 30:36:@6574.4]
  wire  _T_25480; // @[Switch.scala 30:53:@6576.4]
  wire  valid_20_42; // @[Switch.scala 30:36:@6577.4]
  wire  _T_25483; // @[Switch.scala 30:53:@6579.4]
  wire  valid_20_43; // @[Switch.scala 30:36:@6580.4]
  wire  _T_25486; // @[Switch.scala 30:53:@6582.4]
  wire  valid_20_44; // @[Switch.scala 30:36:@6583.4]
  wire  _T_25489; // @[Switch.scala 30:53:@6585.4]
  wire  valid_20_45; // @[Switch.scala 30:36:@6586.4]
  wire  _T_25492; // @[Switch.scala 30:53:@6588.4]
  wire  valid_20_46; // @[Switch.scala 30:36:@6589.4]
  wire  _T_25495; // @[Switch.scala 30:53:@6591.4]
  wire  valid_20_47; // @[Switch.scala 30:36:@6592.4]
  wire  _T_25498; // @[Switch.scala 30:53:@6594.4]
  wire  valid_20_48; // @[Switch.scala 30:36:@6595.4]
  wire  _T_25501; // @[Switch.scala 30:53:@6597.4]
  wire  valid_20_49; // @[Switch.scala 30:36:@6598.4]
  wire  _T_25504; // @[Switch.scala 30:53:@6600.4]
  wire  valid_20_50; // @[Switch.scala 30:36:@6601.4]
  wire  _T_25507; // @[Switch.scala 30:53:@6603.4]
  wire  valid_20_51; // @[Switch.scala 30:36:@6604.4]
  wire  _T_25510; // @[Switch.scala 30:53:@6606.4]
  wire  valid_20_52; // @[Switch.scala 30:36:@6607.4]
  wire  _T_25513; // @[Switch.scala 30:53:@6609.4]
  wire  valid_20_53; // @[Switch.scala 30:36:@6610.4]
  wire  _T_25516; // @[Switch.scala 30:53:@6612.4]
  wire  valid_20_54; // @[Switch.scala 30:36:@6613.4]
  wire  _T_25519; // @[Switch.scala 30:53:@6615.4]
  wire  valid_20_55; // @[Switch.scala 30:36:@6616.4]
  wire  _T_25522; // @[Switch.scala 30:53:@6618.4]
  wire  valid_20_56; // @[Switch.scala 30:36:@6619.4]
  wire  _T_25525; // @[Switch.scala 30:53:@6621.4]
  wire  valid_20_57; // @[Switch.scala 30:36:@6622.4]
  wire  _T_25528; // @[Switch.scala 30:53:@6624.4]
  wire  valid_20_58; // @[Switch.scala 30:36:@6625.4]
  wire  _T_25531; // @[Switch.scala 30:53:@6627.4]
  wire  valid_20_59; // @[Switch.scala 30:36:@6628.4]
  wire  _T_25534; // @[Switch.scala 30:53:@6630.4]
  wire  valid_20_60; // @[Switch.scala 30:36:@6631.4]
  wire  _T_25537; // @[Switch.scala 30:53:@6633.4]
  wire  valid_20_61; // @[Switch.scala 30:36:@6634.4]
  wire  _T_25540; // @[Switch.scala 30:53:@6636.4]
  wire  valid_20_62; // @[Switch.scala 30:36:@6637.4]
  wire  _T_25543; // @[Switch.scala 30:53:@6639.4]
  wire  valid_20_63; // @[Switch.scala 30:36:@6640.4]
  wire [5:0] _T_25609; // @[Mux.scala 31:69:@6642.4]
  wire [5:0] _T_25610; // @[Mux.scala 31:69:@6643.4]
  wire [5:0] _T_25611; // @[Mux.scala 31:69:@6644.4]
  wire [5:0] _T_25612; // @[Mux.scala 31:69:@6645.4]
  wire [5:0] _T_25613; // @[Mux.scala 31:69:@6646.4]
  wire [5:0] _T_25614; // @[Mux.scala 31:69:@6647.4]
  wire [5:0] _T_25615; // @[Mux.scala 31:69:@6648.4]
  wire [5:0] _T_25616; // @[Mux.scala 31:69:@6649.4]
  wire [5:0] _T_25617; // @[Mux.scala 31:69:@6650.4]
  wire [5:0] _T_25618; // @[Mux.scala 31:69:@6651.4]
  wire [5:0] _T_25619; // @[Mux.scala 31:69:@6652.4]
  wire [5:0] _T_25620; // @[Mux.scala 31:69:@6653.4]
  wire [5:0] _T_25621; // @[Mux.scala 31:69:@6654.4]
  wire [5:0] _T_25622; // @[Mux.scala 31:69:@6655.4]
  wire [5:0] _T_25623; // @[Mux.scala 31:69:@6656.4]
  wire [5:0] _T_25624; // @[Mux.scala 31:69:@6657.4]
  wire [5:0] _T_25625; // @[Mux.scala 31:69:@6658.4]
  wire [5:0] _T_25626; // @[Mux.scala 31:69:@6659.4]
  wire [5:0] _T_25627; // @[Mux.scala 31:69:@6660.4]
  wire [5:0] _T_25628; // @[Mux.scala 31:69:@6661.4]
  wire [5:0] _T_25629; // @[Mux.scala 31:69:@6662.4]
  wire [5:0] _T_25630; // @[Mux.scala 31:69:@6663.4]
  wire [5:0] _T_25631; // @[Mux.scala 31:69:@6664.4]
  wire [5:0] _T_25632; // @[Mux.scala 31:69:@6665.4]
  wire [5:0] _T_25633; // @[Mux.scala 31:69:@6666.4]
  wire [5:0] _T_25634; // @[Mux.scala 31:69:@6667.4]
  wire [5:0] _T_25635; // @[Mux.scala 31:69:@6668.4]
  wire [5:0] _T_25636; // @[Mux.scala 31:69:@6669.4]
  wire [5:0] _T_25637; // @[Mux.scala 31:69:@6670.4]
  wire [5:0] _T_25638; // @[Mux.scala 31:69:@6671.4]
  wire [5:0] _T_25639; // @[Mux.scala 31:69:@6672.4]
  wire [5:0] _T_25640; // @[Mux.scala 31:69:@6673.4]
  wire [5:0] _T_25641; // @[Mux.scala 31:69:@6674.4]
  wire [5:0] _T_25642; // @[Mux.scala 31:69:@6675.4]
  wire [5:0] _T_25643; // @[Mux.scala 31:69:@6676.4]
  wire [5:0] _T_25644; // @[Mux.scala 31:69:@6677.4]
  wire [5:0] _T_25645; // @[Mux.scala 31:69:@6678.4]
  wire [5:0] _T_25646; // @[Mux.scala 31:69:@6679.4]
  wire [5:0] _T_25647; // @[Mux.scala 31:69:@6680.4]
  wire [5:0] _T_25648; // @[Mux.scala 31:69:@6681.4]
  wire [5:0] _T_25649; // @[Mux.scala 31:69:@6682.4]
  wire [5:0] _T_25650; // @[Mux.scala 31:69:@6683.4]
  wire [5:0] _T_25651; // @[Mux.scala 31:69:@6684.4]
  wire [5:0] _T_25652; // @[Mux.scala 31:69:@6685.4]
  wire [5:0] _T_25653; // @[Mux.scala 31:69:@6686.4]
  wire [5:0] _T_25654; // @[Mux.scala 31:69:@6687.4]
  wire [5:0] _T_25655; // @[Mux.scala 31:69:@6688.4]
  wire [5:0] _T_25656; // @[Mux.scala 31:69:@6689.4]
  wire [5:0] _T_25657; // @[Mux.scala 31:69:@6690.4]
  wire [5:0] _T_25658; // @[Mux.scala 31:69:@6691.4]
  wire [5:0] _T_25659; // @[Mux.scala 31:69:@6692.4]
  wire [5:0] _T_25660; // @[Mux.scala 31:69:@6693.4]
  wire [5:0] _T_25661; // @[Mux.scala 31:69:@6694.4]
  wire [5:0] _T_25662; // @[Mux.scala 31:69:@6695.4]
  wire [5:0] _T_25663; // @[Mux.scala 31:69:@6696.4]
  wire [5:0] _T_25664; // @[Mux.scala 31:69:@6697.4]
  wire [5:0] _T_25665; // @[Mux.scala 31:69:@6698.4]
  wire [5:0] _T_25666; // @[Mux.scala 31:69:@6699.4]
  wire [5:0] _T_25667; // @[Mux.scala 31:69:@6700.4]
  wire [5:0] _T_25668; // @[Mux.scala 31:69:@6701.4]
  wire [5:0] _T_25669; // @[Mux.scala 31:69:@6702.4]
  wire [5:0] _T_25670; // @[Mux.scala 31:69:@6703.4]
  wire [5:0] select_20; // @[Mux.scala 31:69:@6704.4]
  wire [47:0] _GEN_1281; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1282; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1283; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1284; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1285; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1286; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1287; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1288; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1289; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1290; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1291; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1292; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1293; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1294; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1295; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1296; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1297; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1298; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1299; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1300; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1301; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1302; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1303; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1304; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1305; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1306; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1307; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1308; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1309; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1310; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1311; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1312; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1313; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1314; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1315; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1316; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1317; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1318; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1319; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1320; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1321; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1322; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1323; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1324; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1325; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1326; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1327; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1328; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1329; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1330; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1331; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1332; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1333; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1334; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1335; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1336; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1337; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1338; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1339; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1340; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1341; // @[Switch.scala 33:19:@6706.4]
  wire [47:0] _GEN_1342; // @[Switch.scala 33:19:@6706.4]
  wire [7:0] _T_25679; // @[Switch.scala 34:32:@6713.4]
  wire [15:0] _T_25687; // @[Switch.scala 34:32:@6721.4]
  wire [7:0] _T_25694; // @[Switch.scala 34:32:@6728.4]
  wire [31:0] _T_25703; // @[Switch.scala 34:32:@6737.4]
  wire [7:0] _T_25710; // @[Switch.scala 34:32:@6744.4]
  wire [15:0] _T_25718; // @[Switch.scala 34:32:@6752.4]
  wire [7:0] _T_25725; // @[Switch.scala 34:32:@6759.4]
  wire [31:0] _T_25734; // @[Switch.scala 34:32:@6768.4]
  wire [63:0] _T_25735; // @[Switch.scala 34:32:@6769.4]
  wire  _T_25739; // @[Switch.scala 30:53:@6772.4]
  wire  valid_21_0; // @[Switch.scala 30:36:@6773.4]
  wire  _T_25742; // @[Switch.scala 30:53:@6775.4]
  wire  valid_21_1; // @[Switch.scala 30:36:@6776.4]
  wire  _T_25745; // @[Switch.scala 30:53:@6778.4]
  wire  valid_21_2; // @[Switch.scala 30:36:@6779.4]
  wire  _T_25748; // @[Switch.scala 30:53:@6781.4]
  wire  valid_21_3; // @[Switch.scala 30:36:@6782.4]
  wire  _T_25751; // @[Switch.scala 30:53:@6784.4]
  wire  valid_21_4; // @[Switch.scala 30:36:@6785.4]
  wire  _T_25754; // @[Switch.scala 30:53:@6787.4]
  wire  valid_21_5; // @[Switch.scala 30:36:@6788.4]
  wire  _T_25757; // @[Switch.scala 30:53:@6790.4]
  wire  valid_21_6; // @[Switch.scala 30:36:@6791.4]
  wire  _T_25760; // @[Switch.scala 30:53:@6793.4]
  wire  valid_21_7; // @[Switch.scala 30:36:@6794.4]
  wire  _T_25763; // @[Switch.scala 30:53:@6796.4]
  wire  valid_21_8; // @[Switch.scala 30:36:@6797.4]
  wire  _T_25766; // @[Switch.scala 30:53:@6799.4]
  wire  valid_21_9; // @[Switch.scala 30:36:@6800.4]
  wire  _T_25769; // @[Switch.scala 30:53:@6802.4]
  wire  valid_21_10; // @[Switch.scala 30:36:@6803.4]
  wire  _T_25772; // @[Switch.scala 30:53:@6805.4]
  wire  valid_21_11; // @[Switch.scala 30:36:@6806.4]
  wire  _T_25775; // @[Switch.scala 30:53:@6808.4]
  wire  valid_21_12; // @[Switch.scala 30:36:@6809.4]
  wire  _T_25778; // @[Switch.scala 30:53:@6811.4]
  wire  valid_21_13; // @[Switch.scala 30:36:@6812.4]
  wire  _T_25781; // @[Switch.scala 30:53:@6814.4]
  wire  valid_21_14; // @[Switch.scala 30:36:@6815.4]
  wire  _T_25784; // @[Switch.scala 30:53:@6817.4]
  wire  valid_21_15; // @[Switch.scala 30:36:@6818.4]
  wire  _T_25787; // @[Switch.scala 30:53:@6820.4]
  wire  valid_21_16; // @[Switch.scala 30:36:@6821.4]
  wire  _T_25790; // @[Switch.scala 30:53:@6823.4]
  wire  valid_21_17; // @[Switch.scala 30:36:@6824.4]
  wire  _T_25793; // @[Switch.scala 30:53:@6826.4]
  wire  valid_21_18; // @[Switch.scala 30:36:@6827.4]
  wire  _T_25796; // @[Switch.scala 30:53:@6829.4]
  wire  valid_21_19; // @[Switch.scala 30:36:@6830.4]
  wire  _T_25799; // @[Switch.scala 30:53:@6832.4]
  wire  valid_21_20; // @[Switch.scala 30:36:@6833.4]
  wire  _T_25802; // @[Switch.scala 30:53:@6835.4]
  wire  valid_21_21; // @[Switch.scala 30:36:@6836.4]
  wire  _T_25805; // @[Switch.scala 30:53:@6838.4]
  wire  valid_21_22; // @[Switch.scala 30:36:@6839.4]
  wire  _T_25808; // @[Switch.scala 30:53:@6841.4]
  wire  valid_21_23; // @[Switch.scala 30:36:@6842.4]
  wire  _T_25811; // @[Switch.scala 30:53:@6844.4]
  wire  valid_21_24; // @[Switch.scala 30:36:@6845.4]
  wire  _T_25814; // @[Switch.scala 30:53:@6847.4]
  wire  valid_21_25; // @[Switch.scala 30:36:@6848.4]
  wire  _T_25817; // @[Switch.scala 30:53:@6850.4]
  wire  valid_21_26; // @[Switch.scala 30:36:@6851.4]
  wire  _T_25820; // @[Switch.scala 30:53:@6853.4]
  wire  valid_21_27; // @[Switch.scala 30:36:@6854.4]
  wire  _T_25823; // @[Switch.scala 30:53:@6856.4]
  wire  valid_21_28; // @[Switch.scala 30:36:@6857.4]
  wire  _T_25826; // @[Switch.scala 30:53:@6859.4]
  wire  valid_21_29; // @[Switch.scala 30:36:@6860.4]
  wire  _T_25829; // @[Switch.scala 30:53:@6862.4]
  wire  valid_21_30; // @[Switch.scala 30:36:@6863.4]
  wire  _T_25832; // @[Switch.scala 30:53:@6865.4]
  wire  valid_21_31; // @[Switch.scala 30:36:@6866.4]
  wire  _T_25835; // @[Switch.scala 30:53:@6868.4]
  wire  valid_21_32; // @[Switch.scala 30:36:@6869.4]
  wire  _T_25838; // @[Switch.scala 30:53:@6871.4]
  wire  valid_21_33; // @[Switch.scala 30:36:@6872.4]
  wire  _T_25841; // @[Switch.scala 30:53:@6874.4]
  wire  valid_21_34; // @[Switch.scala 30:36:@6875.4]
  wire  _T_25844; // @[Switch.scala 30:53:@6877.4]
  wire  valid_21_35; // @[Switch.scala 30:36:@6878.4]
  wire  _T_25847; // @[Switch.scala 30:53:@6880.4]
  wire  valid_21_36; // @[Switch.scala 30:36:@6881.4]
  wire  _T_25850; // @[Switch.scala 30:53:@6883.4]
  wire  valid_21_37; // @[Switch.scala 30:36:@6884.4]
  wire  _T_25853; // @[Switch.scala 30:53:@6886.4]
  wire  valid_21_38; // @[Switch.scala 30:36:@6887.4]
  wire  _T_25856; // @[Switch.scala 30:53:@6889.4]
  wire  valid_21_39; // @[Switch.scala 30:36:@6890.4]
  wire  _T_25859; // @[Switch.scala 30:53:@6892.4]
  wire  valid_21_40; // @[Switch.scala 30:36:@6893.4]
  wire  _T_25862; // @[Switch.scala 30:53:@6895.4]
  wire  valid_21_41; // @[Switch.scala 30:36:@6896.4]
  wire  _T_25865; // @[Switch.scala 30:53:@6898.4]
  wire  valid_21_42; // @[Switch.scala 30:36:@6899.4]
  wire  _T_25868; // @[Switch.scala 30:53:@6901.4]
  wire  valid_21_43; // @[Switch.scala 30:36:@6902.4]
  wire  _T_25871; // @[Switch.scala 30:53:@6904.4]
  wire  valid_21_44; // @[Switch.scala 30:36:@6905.4]
  wire  _T_25874; // @[Switch.scala 30:53:@6907.4]
  wire  valid_21_45; // @[Switch.scala 30:36:@6908.4]
  wire  _T_25877; // @[Switch.scala 30:53:@6910.4]
  wire  valid_21_46; // @[Switch.scala 30:36:@6911.4]
  wire  _T_25880; // @[Switch.scala 30:53:@6913.4]
  wire  valid_21_47; // @[Switch.scala 30:36:@6914.4]
  wire  _T_25883; // @[Switch.scala 30:53:@6916.4]
  wire  valid_21_48; // @[Switch.scala 30:36:@6917.4]
  wire  _T_25886; // @[Switch.scala 30:53:@6919.4]
  wire  valid_21_49; // @[Switch.scala 30:36:@6920.4]
  wire  _T_25889; // @[Switch.scala 30:53:@6922.4]
  wire  valid_21_50; // @[Switch.scala 30:36:@6923.4]
  wire  _T_25892; // @[Switch.scala 30:53:@6925.4]
  wire  valid_21_51; // @[Switch.scala 30:36:@6926.4]
  wire  _T_25895; // @[Switch.scala 30:53:@6928.4]
  wire  valid_21_52; // @[Switch.scala 30:36:@6929.4]
  wire  _T_25898; // @[Switch.scala 30:53:@6931.4]
  wire  valid_21_53; // @[Switch.scala 30:36:@6932.4]
  wire  _T_25901; // @[Switch.scala 30:53:@6934.4]
  wire  valid_21_54; // @[Switch.scala 30:36:@6935.4]
  wire  _T_25904; // @[Switch.scala 30:53:@6937.4]
  wire  valid_21_55; // @[Switch.scala 30:36:@6938.4]
  wire  _T_25907; // @[Switch.scala 30:53:@6940.4]
  wire  valid_21_56; // @[Switch.scala 30:36:@6941.4]
  wire  _T_25910; // @[Switch.scala 30:53:@6943.4]
  wire  valid_21_57; // @[Switch.scala 30:36:@6944.4]
  wire  _T_25913; // @[Switch.scala 30:53:@6946.4]
  wire  valid_21_58; // @[Switch.scala 30:36:@6947.4]
  wire  _T_25916; // @[Switch.scala 30:53:@6949.4]
  wire  valid_21_59; // @[Switch.scala 30:36:@6950.4]
  wire  _T_25919; // @[Switch.scala 30:53:@6952.4]
  wire  valid_21_60; // @[Switch.scala 30:36:@6953.4]
  wire  _T_25922; // @[Switch.scala 30:53:@6955.4]
  wire  valid_21_61; // @[Switch.scala 30:36:@6956.4]
  wire  _T_25925; // @[Switch.scala 30:53:@6958.4]
  wire  valid_21_62; // @[Switch.scala 30:36:@6959.4]
  wire  _T_25928; // @[Switch.scala 30:53:@6961.4]
  wire  valid_21_63; // @[Switch.scala 30:36:@6962.4]
  wire [5:0] _T_25994; // @[Mux.scala 31:69:@6964.4]
  wire [5:0] _T_25995; // @[Mux.scala 31:69:@6965.4]
  wire [5:0] _T_25996; // @[Mux.scala 31:69:@6966.4]
  wire [5:0] _T_25997; // @[Mux.scala 31:69:@6967.4]
  wire [5:0] _T_25998; // @[Mux.scala 31:69:@6968.4]
  wire [5:0] _T_25999; // @[Mux.scala 31:69:@6969.4]
  wire [5:0] _T_26000; // @[Mux.scala 31:69:@6970.4]
  wire [5:0] _T_26001; // @[Mux.scala 31:69:@6971.4]
  wire [5:0] _T_26002; // @[Mux.scala 31:69:@6972.4]
  wire [5:0] _T_26003; // @[Mux.scala 31:69:@6973.4]
  wire [5:0] _T_26004; // @[Mux.scala 31:69:@6974.4]
  wire [5:0] _T_26005; // @[Mux.scala 31:69:@6975.4]
  wire [5:0] _T_26006; // @[Mux.scala 31:69:@6976.4]
  wire [5:0] _T_26007; // @[Mux.scala 31:69:@6977.4]
  wire [5:0] _T_26008; // @[Mux.scala 31:69:@6978.4]
  wire [5:0] _T_26009; // @[Mux.scala 31:69:@6979.4]
  wire [5:0] _T_26010; // @[Mux.scala 31:69:@6980.4]
  wire [5:0] _T_26011; // @[Mux.scala 31:69:@6981.4]
  wire [5:0] _T_26012; // @[Mux.scala 31:69:@6982.4]
  wire [5:0] _T_26013; // @[Mux.scala 31:69:@6983.4]
  wire [5:0] _T_26014; // @[Mux.scala 31:69:@6984.4]
  wire [5:0] _T_26015; // @[Mux.scala 31:69:@6985.4]
  wire [5:0] _T_26016; // @[Mux.scala 31:69:@6986.4]
  wire [5:0] _T_26017; // @[Mux.scala 31:69:@6987.4]
  wire [5:0] _T_26018; // @[Mux.scala 31:69:@6988.4]
  wire [5:0] _T_26019; // @[Mux.scala 31:69:@6989.4]
  wire [5:0] _T_26020; // @[Mux.scala 31:69:@6990.4]
  wire [5:0] _T_26021; // @[Mux.scala 31:69:@6991.4]
  wire [5:0] _T_26022; // @[Mux.scala 31:69:@6992.4]
  wire [5:0] _T_26023; // @[Mux.scala 31:69:@6993.4]
  wire [5:0] _T_26024; // @[Mux.scala 31:69:@6994.4]
  wire [5:0] _T_26025; // @[Mux.scala 31:69:@6995.4]
  wire [5:0] _T_26026; // @[Mux.scala 31:69:@6996.4]
  wire [5:0] _T_26027; // @[Mux.scala 31:69:@6997.4]
  wire [5:0] _T_26028; // @[Mux.scala 31:69:@6998.4]
  wire [5:0] _T_26029; // @[Mux.scala 31:69:@6999.4]
  wire [5:0] _T_26030; // @[Mux.scala 31:69:@7000.4]
  wire [5:0] _T_26031; // @[Mux.scala 31:69:@7001.4]
  wire [5:0] _T_26032; // @[Mux.scala 31:69:@7002.4]
  wire [5:0] _T_26033; // @[Mux.scala 31:69:@7003.4]
  wire [5:0] _T_26034; // @[Mux.scala 31:69:@7004.4]
  wire [5:0] _T_26035; // @[Mux.scala 31:69:@7005.4]
  wire [5:0] _T_26036; // @[Mux.scala 31:69:@7006.4]
  wire [5:0] _T_26037; // @[Mux.scala 31:69:@7007.4]
  wire [5:0] _T_26038; // @[Mux.scala 31:69:@7008.4]
  wire [5:0] _T_26039; // @[Mux.scala 31:69:@7009.4]
  wire [5:0] _T_26040; // @[Mux.scala 31:69:@7010.4]
  wire [5:0] _T_26041; // @[Mux.scala 31:69:@7011.4]
  wire [5:0] _T_26042; // @[Mux.scala 31:69:@7012.4]
  wire [5:0] _T_26043; // @[Mux.scala 31:69:@7013.4]
  wire [5:0] _T_26044; // @[Mux.scala 31:69:@7014.4]
  wire [5:0] _T_26045; // @[Mux.scala 31:69:@7015.4]
  wire [5:0] _T_26046; // @[Mux.scala 31:69:@7016.4]
  wire [5:0] _T_26047; // @[Mux.scala 31:69:@7017.4]
  wire [5:0] _T_26048; // @[Mux.scala 31:69:@7018.4]
  wire [5:0] _T_26049; // @[Mux.scala 31:69:@7019.4]
  wire [5:0] _T_26050; // @[Mux.scala 31:69:@7020.4]
  wire [5:0] _T_26051; // @[Mux.scala 31:69:@7021.4]
  wire [5:0] _T_26052; // @[Mux.scala 31:69:@7022.4]
  wire [5:0] _T_26053; // @[Mux.scala 31:69:@7023.4]
  wire [5:0] _T_26054; // @[Mux.scala 31:69:@7024.4]
  wire [5:0] _T_26055; // @[Mux.scala 31:69:@7025.4]
  wire [5:0] select_21; // @[Mux.scala 31:69:@7026.4]
  wire [47:0] _GEN_1345; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1346; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1347; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1348; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1349; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1350; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1351; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1352; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1353; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1354; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1355; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1356; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1357; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1358; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1359; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1360; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1361; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1362; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1363; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1364; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1365; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1366; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1367; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1368; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1369; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1370; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1371; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1372; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1373; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1374; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1375; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1376; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1377; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1378; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1379; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1380; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1381; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1382; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1383; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1384; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1385; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1386; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1387; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1388; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1389; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1390; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1391; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1392; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1393; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1394; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1395; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1396; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1397; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1398; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1399; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1400; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1401; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1402; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1403; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1404; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1405; // @[Switch.scala 33:19:@7028.4]
  wire [47:0] _GEN_1406; // @[Switch.scala 33:19:@7028.4]
  wire [7:0] _T_26064; // @[Switch.scala 34:32:@7035.4]
  wire [15:0] _T_26072; // @[Switch.scala 34:32:@7043.4]
  wire [7:0] _T_26079; // @[Switch.scala 34:32:@7050.4]
  wire [31:0] _T_26088; // @[Switch.scala 34:32:@7059.4]
  wire [7:0] _T_26095; // @[Switch.scala 34:32:@7066.4]
  wire [15:0] _T_26103; // @[Switch.scala 34:32:@7074.4]
  wire [7:0] _T_26110; // @[Switch.scala 34:32:@7081.4]
  wire [31:0] _T_26119; // @[Switch.scala 34:32:@7090.4]
  wire [63:0] _T_26120; // @[Switch.scala 34:32:@7091.4]
  wire  _T_26124; // @[Switch.scala 30:53:@7094.4]
  wire  valid_22_0; // @[Switch.scala 30:36:@7095.4]
  wire  _T_26127; // @[Switch.scala 30:53:@7097.4]
  wire  valid_22_1; // @[Switch.scala 30:36:@7098.4]
  wire  _T_26130; // @[Switch.scala 30:53:@7100.4]
  wire  valid_22_2; // @[Switch.scala 30:36:@7101.4]
  wire  _T_26133; // @[Switch.scala 30:53:@7103.4]
  wire  valid_22_3; // @[Switch.scala 30:36:@7104.4]
  wire  _T_26136; // @[Switch.scala 30:53:@7106.4]
  wire  valid_22_4; // @[Switch.scala 30:36:@7107.4]
  wire  _T_26139; // @[Switch.scala 30:53:@7109.4]
  wire  valid_22_5; // @[Switch.scala 30:36:@7110.4]
  wire  _T_26142; // @[Switch.scala 30:53:@7112.4]
  wire  valid_22_6; // @[Switch.scala 30:36:@7113.4]
  wire  _T_26145; // @[Switch.scala 30:53:@7115.4]
  wire  valid_22_7; // @[Switch.scala 30:36:@7116.4]
  wire  _T_26148; // @[Switch.scala 30:53:@7118.4]
  wire  valid_22_8; // @[Switch.scala 30:36:@7119.4]
  wire  _T_26151; // @[Switch.scala 30:53:@7121.4]
  wire  valid_22_9; // @[Switch.scala 30:36:@7122.4]
  wire  _T_26154; // @[Switch.scala 30:53:@7124.4]
  wire  valid_22_10; // @[Switch.scala 30:36:@7125.4]
  wire  _T_26157; // @[Switch.scala 30:53:@7127.4]
  wire  valid_22_11; // @[Switch.scala 30:36:@7128.4]
  wire  _T_26160; // @[Switch.scala 30:53:@7130.4]
  wire  valid_22_12; // @[Switch.scala 30:36:@7131.4]
  wire  _T_26163; // @[Switch.scala 30:53:@7133.4]
  wire  valid_22_13; // @[Switch.scala 30:36:@7134.4]
  wire  _T_26166; // @[Switch.scala 30:53:@7136.4]
  wire  valid_22_14; // @[Switch.scala 30:36:@7137.4]
  wire  _T_26169; // @[Switch.scala 30:53:@7139.4]
  wire  valid_22_15; // @[Switch.scala 30:36:@7140.4]
  wire  _T_26172; // @[Switch.scala 30:53:@7142.4]
  wire  valid_22_16; // @[Switch.scala 30:36:@7143.4]
  wire  _T_26175; // @[Switch.scala 30:53:@7145.4]
  wire  valid_22_17; // @[Switch.scala 30:36:@7146.4]
  wire  _T_26178; // @[Switch.scala 30:53:@7148.4]
  wire  valid_22_18; // @[Switch.scala 30:36:@7149.4]
  wire  _T_26181; // @[Switch.scala 30:53:@7151.4]
  wire  valid_22_19; // @[Switch.scala 30:36:@7152.4]
  wire  _T_26184; // @[Switch.scala 30:53:@7154.4]
  wire  valid_22_20; // @[Switch.scala 30:36:@7155.4]
  wire  _T_26187; // @[Switch.scala 30:53:@7157.4]
  wire  valid_22_21; // @[Switch.scala 30:36:@7158.4]
  wire  _T_26190; // @[Switch.scala 30:53:@7160.4]
  wire  valid_22_22; // @[Switch.scala 30:36:@7161.4]
  wire  _T_26193; // @[Switch.scala 30:53:@7163.4]
  wire  valid_22_23; // @[Switch.scala 30:36:@7164.4]
  wire  _T_26196; // @[Switch.scala 30:53:@7166.4]
  wire  valid_22_24; // @[Switch.scala 30:36:@7167.4]
  wire  _T_26199; // @[Switch.scala 30:53:@7169.4]
  wire  valid_22_25; // @[Switch.scala 30:36:@7170.4]
  wire  _T_26202; // @[Switch.scala 30:53:@7172.4]
  wire  valid_22_26; // @[Switch.scala 30:36:@7173.4]
  wire  _T_26205; // @[Switch.scala 30:53:@7175.4]
  wire  valid_22_27; // @[Switch.scala 30:36:@7176.4]
  wire  _T_26208; // @[Switch.scala 30:53:@7178.4]
  wire  valid_22_28; // @[Switch.scala 30:36:@7179.4]
  wire  _T_26211; // @[Switch.scala 30:53:@7181.4]
  wire  valid_22_29; // @[Switch.scala 30:36:@7182.4]
  wire  _T_26214; // @[Switch.scala 30:53:@7184.4]
  wire  valid_22_30; // @[Switch.scala 30:36:@7185.4]
  wire  _T_26217; // @[Switch.scala 30:53:@7187.4]
  wire  valid_22_31; // @[Switch.scala 30:36:@7188.4]
  wire  _T_26220; // @[Switch.scala 30:53:@7190.4]
  wire  valid_22_32; // @[Switch.scala 30:36:@7191.4]
  wire  _T_26223; // @[Switch.scala 30:53:@7193.4]
  wire  valid_22_33; // @[Switch.scala 30:36:@7194.4]
  wire  _T_26226; // @[Switch.scala 30:53:@7196.4]
  wire  valid_22_34; // @[Switch.scala 30:36:@7197.4]
  wire  _T_26229; // @[Switch.scala 30:53:@7199.4]
  wire  valid_22_35; // @[Switch.scala 30:36:@7200.4]
  wire  _T_26232; // @[Switch.scala 30:53:@7202.4]
  wire  valid_22_36; // @[Switch.scala 30:36:@7203.4]
  wire  _T_26235; // @[Switch.scala 30:53:@7205.4]
  wire  valid_22_37; // @[Switch.scala 30:36:@7206.4]
  wire  _T_26238; // @[Switch.scala 30:53:@7208.4]
  wire  valid_22_38; // @[Switch.scala 30:36:@7209.4]
  wire  _T_26241; // @[Switch.scala 30:53:@7211.4]
  wire  valid_22_39; // @[Switch.scala 30:36:@7212.4]
  wire  _T_26244; // @[Switch.scala 30:53:@7214.4]
  wire  valid_22_40; // @[Switch.scala 30:36:@7215.4]
  wire  _T_26247; // @[Switch.scala 30:53:@7217.4]
  wire  valid_22_41; // @[Switch.scala 30:36:@7218.4]
  wire  _T_26250; // @[Switch.scala 30:53:@7220.4]
  wire  valid_22_42; // @[Switch.scala 30:36:@7221.4]
  wire  _T_26253; // @[Switch.scala 30:53:@7223.4]
  wire  valid_22_43; // @[Switch.scala 30:36:@7224.4]
  wire  _T_26256; // @[Switch.scala 30:53:@7226.4]
  wire  valid_22_44; // @[Switch.scala 30:36:@7227.4]
  wire  _T_26259; // @[Switch.scala 30:53:@7229.4]
  wire  valid_22_45; // @[Switch.scala 30:36:@7230.4]
  wire  _T_26262; // @[Switch.scala 30:53:@7232.4]
  wire  valid_22_46; // @[Switch.scala 30:36:@7233.4]
  wire  _T_26265; // @[Switch.scala 30:53:@7235.4]
  wire  valid_22_47; // @[Switch.scala 30:36:@7236.4]
  wire  _T_26268; // @[Switch.scala 30:53:@7238.4]
  wire  valid_22_48; // @[Switch.scala 30:36:@7239.4]
  wire  _T_26271; // @[Switch.scala 30:53:@7241.4]
  wire  valid_22_49; // @[Switch.scala 30:36:@7242.4]
  wire  _T_26274; // @[Switch.scala 30:53:@7244.4]
  wire  valid_22_50; // @[Switch.scala 30:36:@7245.4]
  wire  _T_26277; // @[Switch.scala 30:53:@7247.4]
  wire  valid_22_51; // @[Switch.scala 30:36:@7248.4]
  wire  _T_26280; // @[Switch.scala 30:53:@7250.4]
  wire  valid_22_52; // @[Switch.scala 30:36:@7251.4]
  wire  _T_26283; // @[Switch.scala 30:53:@7253.4]
  wire  valid_22_53; // @[Switch.scala 30:36:@7254.4]
  wire  _T_26286; // @[Switch.scala 30:53:@7256.4]
  wire  valid_22_54; // @[Switch.scala 30:36:@7257.4]
  wire  _T_26289; // @[Switch.scala 30:53:@7259.4]
  wire  valid_22_55; // @[Switch.scala 30:36:@7260.4]
  wire  _T_26292; // @[Switch.scala 30:53:@7262.4]
  wire  valid_22_56; // @[Switch.scala 30:36:@7263.4]
  wire  _T_26295; // @[Switch.scala 30:53:@7265.4]
  wire  valid_22_57; // @[Switch.scala 30:36:@7266.4]
  wire  _T_26298; // @[Switch.scala 30:53:@7268.4]
  wire  valid_22_58; // @[Switch.scala 30:36:@7269.4]
  wire  _T_26301; // @[Switch.scala 30:53:@7271.4]
  wire  valid_22_59; // @[Switch.scala 30:36:@7272.4]
  wire  _T_26304; // @[Switch.scala 30:53:@7274.4]
  wire  valid_22_60; // @[Switch.scala 30:36:@7275.4]
  wire  _T_26307; // @[Switch.scala 30:53:@7277.4]
  wire  valid_22_61; // @[Switch.scala 30:36:@7278.4]
  wire  _T_26310; // @[Switch.scala 30:53:@7280.4]
  wire  valid_22_62; // @[Switch.scala 30:36:@7281.4]
  wire  _T_26313; // @[Switch.scala 30:53:@7283.4]
  wire  valid_22_63; // @[Switch.scala 30:36:@7284.4]
  wire [5:0] _T_26379; // @[Mux.scala 31:69:@7286.4]
  wire [5:0] _T_26380; // @[Mux.scala 31:69:@7287.4]
  wire [5:0] _T_26381; // @[Mux.scala 31:69:@7288.4]
  wire [5:0] _T_26382; // @[Mux.scala 31:69:@7289.4]
  wire [5:0] _T_26383; // @[Mux.scala 31:69:@7290.4]
  wire [5:0] _T_26384; // @[Mux.scala 31:69:@7291.4]
  wire [5:0] _T_26385; // @[Mux.scala 31:69:@7292.4]
  wire [5:0] _T_26386; // @[Mux.scala 31:69:@7293.4]
  wire [5:0] _T_26387; // @[Mux.scala 31:69:@7294.4]
  wire [5:0] _T_26388; // @[Mux.scala 31:69:@7295.4]
  wire [5:0] _T_26389; // @[Mux.scala 31:69:@7296.4]
  wire [5:0] _T_26390; // @[Mux.scala 31:69:@7297.4]
  wire [5:0] _T_26391; // @[Mux.scala 31:69:@7298.4]
  wire [5:0] _T_26392; // @[Mux.scala 31:69:@7299.4]
  wire [5:0] _T_26393; // @[Mux.scala 31:69:@7300.4]
  wire [5:0] _T_26394; // @[Mux.scala 31:69:@7301.4]
  wire [5:0] _T_26395; // @[Mux.scala 31:69:@7302.4]
  wire [5:0] _T_26396; // @[Mux.scala 31:69:@7303.4]
  wire [5:0] _T_26397; // @[Mux.scala 31:69:@7304.4]
  wire [5:0] _T_26398; // @[Mux.scala 31:69:@7305.4]
  wire [5:0] _T_26399; // @[Mux.scala 31:69:@7306.4]
  wire [5:0] _T_26400; // @[Mux.scala 31:69:@7307.4]
  wire [5:0] _T_26401; // @[Mux.scala 31:69:@7308.4]
  wire [5:0] _T_26402; // @[Mux.scala 31:69:@7309.4]
  wire [5:0] _T_26403; // @[Mux.scala 31:69:@7310.4]
  wire [5:0] _T_26404; // @[Mux.scala 31:69:@7311.4]
  wire [5:0] _T_26405; // @[Mux.scala 31:69:@7312.4]
  wire [5:0] _T_26406; // @[Mux.scala 31:69:@7313.4]
  wire [5:0] _T_26407; // @[Mux.scala 31:69:@7314.4]
  wire [5:0] _T_26408; // @[Mux.scala 31:69:@7315.4]
  wire [5:0] _T_26409; // @[Mux.scala 31:69:@7316.4]
  wire [5:0] _T_26410; // @[Mux.scala 31:69:@7317.4]
  wire [5:0] _T_26411; // @[Mux.scala 31:69:@7318.4]
  wire [5:0] _T_26412; // @[Mux.scala 31:69:@7319.4]
  wire [5:0] _T_26413; // @[Mux.scala 31:69:@7320.4]
  wire [5:0] _T_26414; // @[Mux.scala 31:69:@7321.4]
  wire [5:0] _T_26415; // @[Mux.scala 31:69:@7322.4]
  wire [5:0] _T_26416; // @[Mux.scala 31:69:@7323.4]
  wire [5:0] _T_26417; // @[Mux.scala 31:69:@7324.4]
  wire [5:0] _T_26418; // @[Mux.scala 31:69:@7325.4]
  wire [5:0] _T_26419; // @[Mux.scala 31:69:@7326.4]
  wire [5:0] _T_26420; // @[Mux.scala 31:69:@7327.4]
  wire [5:0] _T_26421; // @[Mux.scala 31:69:@7328.4]
  wire [5:0] _T_26422; // @[Mux.scala 31:69:@7329.4]
  wire [5:0] _T_26423; // @[Mux.scala 31:69:@7330.4]
  wire [5:0] _T_26424; // @[Mux.scala 31:69:@7331.4]
  wire [5:0] _T_26425; // @[Mux.scala 31:69:@7332.4]
  wire [5:0] _T_26426; // @[Mux.scala 31:69:@7333.4]
  wire [5:0] _T_26427; // @[Mux.scala 31:69:@7334.4]
  wire [5:0] _T_26428; // @[Mux.scala 31:69:@7335.4]
  wire [5:0] _T_26429; // @[Mux.scala 31:69:@7336.4]
  wire [5:0] _T_26430; // @[Mux.scala 31:69:@7337.4]
  wire [5:0] _T_26431; // @[Mux.scala 31:69:@7338.4]
  wire [5:0] _T_26432; // @[Mux.scala 31:69:@7339.4]
  wire [5:0] _T_26433; // @[Mux.scala 31:69:@7340.4]
  wire [5:0] _T_26434; // @[Mux.scala 31:69:@7341.4]
  wire [5:0] _T_26435; // @[Mux.scala 31:69:@7342.4]
  wire [5:0] _T_26436; // @[Mux.scala 31:69:@7343.4]
  wire [5:0] _T_26437; // @[Mux.scala 31:69:@7344.4]
  wire [5:0] _T_26438; // @[Mux.scala 31:69:@7345.4]
  wire [5:0] _T_26439; // @[Mux.scala 31:69:@7346.4]
  wire [5:0] _T_26440; // @[Mux.scala 31:69:@7347.4]
  wire [5:0] select_22; // @[Mux.scala 31:69:@7348.4]
  wire [47:0] _GEN_1409; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1410; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1411; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1412; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1413; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1414; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1415; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1416; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1417; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1418; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1419; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1420; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1421; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1422; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1423; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1424; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1425; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1426; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1427; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1428; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1429; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1430; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1431; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1432; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1433; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1434; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1435; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1436; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1437; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1438; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1439; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1440; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1441; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1442; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1443; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1444; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1445; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1446; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1447; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1448; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1449; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1450; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1451; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1452; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1453; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1454; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1455; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1456; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1457; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1458; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1459; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1460; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1461; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1462; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1463; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1464; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1465; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1466; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1467; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1468; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1469; // @[Switch.scala 33:19:@7350.4]
  wire [47:0] _GEN_1470; // @[Switch.scala 33:19:@7350.4]
  wire [7:0] _T_26449; // @[Switch.scala 34:32:@7357.4]
  wire [15:0] _T_26457; // @[Switch.scala 34:32:@7365.4]
  wire [7:0] _T_26464; // @[Switch.scala 34:32:@7372.4]
  wire [31:0] _T_26473; // @[Switch.scala 34:32:@7381.4]
  wire [7:0] _T_26480; // @[Switch.scala 34:32:@7388.4]
  wire [15:0] _T_26488; // @[Switch.scala 34:32:@7396.4]
  wire [7:0] _T_26495; // @[Switch.scala 34:32:@7403.4]
  wire [31:0] _T_26504; // @[Switch.scala 34:32:@7412.4]
  wire [63:0] _T_26505; // @[Switch.scala 34:32:@7413.4]
  wire  _T_26509; // @[Switch.scala 30:53:@7416.4]
  wire  valid_23_0; // @[Switch.scala 30:36:@7417.4]
  wire  _T_26512; // @[Switch.scala 30:53:@7419.4]
  wire  valid_23_1; // @[Switch.scala 30:36:@7420.4]
  wire  _T_26515; // @[Switch.scala 30:53:@7422.4]
  wire  valid_23_2; // @[Switch.scala 30:36:@7423.4]
  wire  _T_26518; // @[Switch.scala 30:53:@7425.4]
  wire  valid_23_3; // @[Switch.scala 30:36:@7426.4]
  wire  _T_26521; // @[Switch.scala 30:53:@7428.4]
  wire  valid_23_4; // @[Switch.scala 30:36:@7429.4]
  wire  _T_26524; // @[Switch.scala 30:53:@7431.4]
  wire  valid_23_5; // @[Switch.scala 30:36:@7432.4]
  wire  _T_26527; // @[Switch.scala 30:53:@7434.4]
  wire  valid_23_6; // @[Switch.scala 30:36:@7435.4]
  wire  _T_26530; // @[Switch.scala 30:53:@7437.4]
  wire  valid_23_7; // @[Switch.scala 30:36:@7438.4]
  wire  _T_26533; // @[Switch.scala 30:53:@7440.4]
  wire  valid_23_8; // @[Switch.scala 30:36:@7441.4]
  wire  _T_26536; // @[Switch.scala 30:53:@7443.4]
  wire  valid_23_9; // @[Switch.scala 30:36:@7444.4]
  wire  _T_26539; // @[Switch.scala 30:53:@7446.4]
  wire  valid_23_10; // @[Switch.scala 30:36:@7447.4]
  wire  _T_26542; // @[Switch.scala 30:53:@7449.4]
  wire  valid_23_11; // @[Switch.scala 30:36:@7450.4]
  wire  _T_26545; // @[Switch.scala 30:53:@7452.4]
  wire  valid_23_12; // @[Switch.scala 30:36:@7453.4]
  wire  _T_26548; // @[Switch.scala 30:53:@7455.4]
  wire  valid_23_13; // @[Switch.scala 30:36:@7456.4]
  wire  _T_26551; // @[Switch.scala 30:53:@7458.4]
  wire  valid_23_14; // @[Switch.scala 30:36:@7459.4]
  wire  _T_26554; // @[Switch.scala 30:53:@7461.4]
  wire  valid_23_15; // @[Switch.scala 30:36:@7462.4]
  wire  _T_26557; // @[Switch.scala 30:53:@7464.4]
  wire  valid_23_16; // @[Switch.scala 30:36:@7465.4]
  wire  _T_26560; // @[Switch.scala 30:53:@7467.4]
  wire  valid_23_17; // @[Switch.scala 30:36:@7468.4]
  wire  _T_26563; // @[Switch.scala 30:53:@7470.4]
  wire  valid_23_18; // @[Switch.scala 30:36:@7471.4]
  wire  _T_26566; // @[Switch.scala 30:53:@7473.4]
  wire  valid_23_19; // @[Switch.scala 30:36:@7474.4]
  wire  _T_26569; // @[Switch.scala 30:53:@7476.4]
  wire  valid_23_20; // @[Switch.scala 30:36:@7477.4]
  wire  _T_26572; // @[Switch.scala 30:53:@7479.4]
  wire  valid_23_21; // @[Switch.scala 30:36:@7480.4]
  wire  _T_26575; // @[Switch.scala 30:53:@7482.4]
  wire  valid_23_22; // @[Switch.scala 30:36:@7483.4]
  wire  _T_26578; // @[Switch.scala 30:53:@7485.4]
  wire  valid_23_23; // @[Switch.scala 30:36:@7486.4]
  wire  _T_26581; // @[Switch.scala 30:53:@7488.4]
  wire  valid_23_24; // @[Switch.scala 30:36:@7489.4]
  wire  _T_26584; // @[Switch.scala 30:53:@7491.4]
  wire  valid_23_25; // @[Switch.scala 30:36:@7492.4]
  wire  _T_26587; // @[Switch.scala 30:53:@7494.4]
  wire  valid_23_26; // @[Switch.scala 30:36:@7495.4]
  wire  _T_26590; // @[Switch.scala 30:53:@7497.4]
  wire  valid_23_27; // @[Switch.scala 30:36:@7498.4]
  wire  _T_26593; // @[Switch.scala 30:53:@7500.4]
  wire  valid_23_28; // @[Switch.scala 30:36:@7501.4]
  wire  _T_26596; // @[Switch.scala 30:53:@7503.4]
  wire  valid_23_29; // @[Switch.scala 30:36:@7504.4]
  wire  _T_26599; // @[Switch.scala 30:53:@7506.4]
  wire  valid_23_30; // @[Switch.scala 30:36:@7507.4]
  wire  _T_26602; // @[Switch.scala 30:53:@7509.4]
  wire  valid_23_31; // @[Switch.scala 30:36:@7510.4]
  wire  _T_26605; // @[Switch.scala 30:53:@7512.4]
  wire  valid_23_32; // @[Switch.scala 30:36:@7513.4]
  wire  _T_26608; // @[Switch.scala 30:53:@7515.4]
  wire  valid_23_33; // @[Switch.scala 30:36:@7516.4]
  wire  _T_26611; // @[Switch.scala 30:53:@7518.4]
  wire  valid_23_34; // @[Switch.scala 30:36:@7519.4]
  wire  _T_26614; // @[Switch.scala 30:53:@7521.4]
  wire  valid_23_35; // @[Switch.scala 30:36:@7522.4]
  wire  _T_26617; // @[Switch.scala 30:53:@7524.4]
  wire  valid_23_36; // @[Switch.scala 30:36:@7525.4]
  wire  _T_26620; // @[Switch.scala 30:53:@7527.4]
  wire  valid_23_37; // @[Switch.scala 30:36:@7528.4]
  wire  _T_26623; // @[Switch.scala 30:53:@7530.4]
  wire  valid_23_38; // @[Switch.scala 30:36:@7531.4]
  wire  _T_26626; // @[Switch.scala 30:53:@7533.4]
  wire  valid_23_39; // @[Switch.scala 30:36:@7534.4]
  wire  _T_26629; // @[Switch.scala 30:53:@7536.4]
  wire  valid_23_40; // @[Switch.scala 30:36:@7537.4]
  wire  _T_26632; // @[Switch.scala 30:53:@7539.4]
  wire  valid_23_41; // @[Switch.scala 30:36:@7540.4]
  wire  _T_26635; // @[Switch.scala 30:53:@7542.4]
  wire  valid_23_42; // @[Switch.scala 30:36:@7543.4]
  wire  _T_26638; // @[Switch.scala 30:53:@7545.4]
  wire  valid_23_43; // @[Switch.scala 30:36:@7546.4]
  wire  _T_26641; // @[Switch.scala 30:53:@7548.4]
  wire  valid_23_44; // @[Switch.scala 30:36:@7549.4]
  wire  _T_26644; // @[Switch.scala 30:53:@7551.4]
  wire  valid_23_45; // @[Switch.scala 30:36:@7552.4]
  wire  _T_26647; // @[Switch.scala 30:53:@7554.4]
  wire  valid_23_46; // @[Switch.scala 30:36:@7555.4]
  wire  _T_26650; // @[Switch.scala 30:53:@7557.4]
  wire  valid_23_47; // @[Switch.scala 30:36:@7558.4]
  wire  _T_26653; // @[Switch.scala 30:53:@7560.4]
  wire  valid_23_48; // @[Switch.scala 30:36:@7561.4]
  wire  _T_26656; // @[Switch.scala 30:53:@7563.4]
  wire  valid_23_49; // @[Switch.scala 30:36:@7564.4]
  wire  _T_26659; // @[Switch.scala 30:53:@7566.4]
  wire  valid_23_50; // @[Switch.scala 30:36:@7567.4]
  wire  _T_26662; // @[Switch.scala 30:53:@7569.4]
  wire  valid_23_51; // @[Switch.scala 30:36:@7570.4]
  wire  _T_26665; // @[Switch.scala 30:53:@7572.4]
  wire  valid_23_52; // @[Switch.scala 30:36:@7573.4]
  wire  _T_26668; // @[Switch.scala 30:53:@7575.4]
  wire  valid_23_53; // @[Switch.scala 30:36:@7576.4]
  wire  _T_26671; // @[Switch.scala 30:53:@7578.4]
  wire  valid_23_54; // @[Switch.scala 30:36:@7579.4]
  wire  _T_26674; // @[Switch.scala 30:53:@7581.4]
  wire  valid_23_55; // @[Switch.scala 30:36:@7582.4]
  wire  _T_26677; // @[Switch.scala 30:53:@7584.4]
  wire  valid_23_56; // @[Switch.scala 30:36:@7585.4]
  wire  _T_26680; // @[Switch.scala 30:53:@7587.4]
  wire  valid_23_57; // @[Switch.scala 30:36:@7588.4]
  wire  _T_26683; // @[Switch.scala 30:53:@7590.4]
  wire  valid_23_58; // @[Switch.scala 30:36:@7591.4]
  wire  _T_26686; // @[Switch.scala 30:53:@7593.4]
  wire  valid_23_59; // @[Switch.scala 30:36:@7594.4]
  wire  _T_26689; // @[Switch.scala 30:53:@7596.4]
  wire  valid_23_60; // @[Switch.scala 30:36:@7597.4]
  wire  _T_26692; // @[Switch.scala 30:53:@7599.4]
  wire  valid_23_61; // @[Switch.scala 30:36:@7600.4]
  wire  _T_26695; // @[Switch.scala 30:53:@7602.4]
  wire  valid_23_62; // @[Switch.scala 30:36:@7603.4]
  wire  _T_26698; // @[Switch.scala 30:53:@7605.4]
  wire  valid_23_63; // @[Switch.scala 30:36:@7606.4]
  wire [5:0] _T_26764; // @[Mux.scala 31:69:@7608.4]
  wire [5:0] _T_26765; // @[Mux.scala 31:69:@7609.4]
  wire [5:0] _T_26766; // @[Mux.scala 31:69:@7610.4]
  wire [5:0] _T_26767; // @[Mux.scala 31:69:@7611.4]
  wire [5:0] _T_26768; // @[Mux.scala 31:69:@7612.4]
  wire [5:0] _T_26769; // @[Mux.scala 31:69:@7613.4]
  wire [5:0] _T_26770; // @[Mux.scala 31:69:@7614.4]
  wire [5:0] _T_26771; // @[Mux.scala 31:69:@7615.4]
  wire [5:0] _T_26772; // @[Mux.scala 31:69:@7616.4]
  wire [5:0] _T_26773; // @[Mux.scala 31:69:@7617.4]
  wire [5:0] _T_26774; // @[Mux.scala 31:69:@7618.4]
  wire [5:0] _T_26775; // @[Mux.scala 31:69:@7619.4]
  wire [5:0] _T_26776; // @[Mux.scala 31:69:@7620.4]
  wire [5:0] _T_26777; // @[Mux.scala 31:69:@7621.4]
  wire [5:0] _T_26778; // @[Mux.scala 31:69:@7622.4]
  wire [5:0] _T_26779; // @[Mux.scala 31:69:@7623.4]
  wire [5:0] _T_26780; // @[Mux.scala 31:69:@7624.4]
  wire [5:0] _T_26781; // @[Mux.scala 31:69:@7625.4]
  wire [5:0] _T_26782; // @[Mux.scala 31:69:@7626.4]
  wire [5:0] _T_26783; // @[Mux.scala 31:69:@7627.4]
  wire [5:0] _T_26784; // @[Mux.scala 31:69:@7628.4]
  wire [5:0] _T_26785; // @[Mux.scala 31:69:@7629.4]
  wire [5:0] _T_26786; // @[Mux.scala 31:69:@7630.4]
  wire [5:0] _T_26787; // @[Mux.scala 31:69:@7631.4]
  wire [5:0] _T_26788; // @[Mux.scala 31:69:@7632.4]
  wire [5:0] _T_26789; // @[Mux.scala 31:69:@7633.4]
  wire [5:0] _T_26790; // @[Mux.scala 31:69:@7634.4]
  wire [5:0] _T_26791; // @[Mux.scala 31:69:@7635.4]
  wire [5:0] _T_26792; // @[Mux.scala 31:69:@7636.4]
  wire [5:0] _T_26793; // @[Mux.scala 31:69:@7637.4]
  wire [5:0] _T_26794; // @[Mux.scala 31:69:@7638.4]
  wire [5:0] _T_26795; // @[Mux.scala 31:69:@7639.4]
  wire [5:0] _T_26796; // @[Mux.scala 31:69:@7640.4]
  wire [5:0] _T_26797; // @[Mux.scala 31:69:@7641.4]
  wire [5:0] _T_26798; // @[Mux.scala 31:69:@7642.4]
  wire [5:0] _T_26799; // @[Mux.scala 31:69:@7643.4]
  wire [5:0] _T_26800; // @[Mux.scala 31:69:@7644.4]
  wire [5:0] _T_26801; // @[Mux.scala 31:69:@7645.4]
  wire [5:0] _T_26802; // @[Mux.scala 31:69:@7646.4]
  wire [5:0] _T_26803; // @[Mux.scala 31:69:@7647.4]
  wire [5:0] _T_26804; // @[Mux.scala 31:69:@7648.4]
  wire [5:0] _T_26805; // @[Mux.scala 31:69:@7649.4]
  wire [5:0] _T_26806; // @[Mux.scala 31:69:@7650.4]
  wire [5:0] _T_26807; // @[Mux.scala 31:69:@7651.4]
  wire [5:0] _T_26808; // @[Mux.scala 31:69:@7652.4]
  wire [5:0] _T_26809; // @[Mux.scala 31:69:@7653.4]
  wire [5:0] _T_26810; // @[Mux.scala 31:69:@7654.4]
  wire [5:0] _T_26811; // @[Mux.scala 31:69:@7655.4]
  wire [5:0] _T_26812; // @[Mux.scala 31:69:@7656.4]
  wire [5:0] _T_26813; // @[Mux.scala 31:69:@7657.4]
  wire [5:0] _T_26814; // @[Mux.scala 31:69:@7658.4]
  wire [5:0] _T_26815; // @[Mux.scala 31:69:@7659.4]
  wire [5:0] _T_26816; // @[Mux.scala 31:69:@7660.4]
  wire [5:0] _T_26817; // @[Mux.scala 31:69:@7661.4]
  wire [5:0] _T_26818; // @[Mux.scala 31:69:@7662.4]
  wire [5:0] _T_26819; // @[Mux.scala 31:69:@7663.4]
  wire [5:0] _T_26820; // @[Mux.scala 31:69:@7664.4]
  wire [5:0] _T_26821; // @[Mux.scala 31:69:@7665.4]
  wire [5:0] _T_26822; // @[Mux.scala 31:69:@7666.4]
  wire [5:0] _T_26823; // @[Mux.scala 31:69:@7667.4]
  wire [5:0] _T_26824; // @[Mux.scala 31:69:@7668.4]
  wire [5:0] _T_26825; // @[Mux.scala 31:69:@7669.4]
  wire [5:0] select_23; // @[Mux.scala 31:69:@7670.4]
  wire [47:0] _GEN_1473; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1474; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1475; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1476; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1477; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1478; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1479; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1480; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1481; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1482; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1483; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1484; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1485; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1486; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1487; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1488; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1489; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1490; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1491; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1492; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1493; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1494; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1495; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1496; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1497; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1498; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1499; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1500; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1501; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1502; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1503; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1504; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1505; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1506; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1507; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1508; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1509; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1510; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1511; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1512; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1513; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1514; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1515; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1516; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1517; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1518; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1519; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1520; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1521; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1522; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1523; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1524; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1525; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1526; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1527; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1528; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1529; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1530; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1531; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1532; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1533; // @[Switch.scala 33:19:@7672.4]
  wire [47:0] _GEN_1534; // @[Switch.scala 33:19:@7672.4]
  wire [7:0] _T_26834; // @[Switch.scala 34:32:@7679.4]
  wire [15:0] _T_26842; // @[Switch.scala 34:32:@7687.4]
  wire [7:0] _T_26849; // @[Switch.scala 34:32:@7694.4]
  wire [31:0] _T_26858; // @[Switch.scala 34:32:@7703.4]
  wire [7:0] _T_26865; // @[Switch.scala 34:32:@7710.4]
  wire [15:0] _T_26873; // @[Switch.scala 34:32:@7718.4]
  wire [7:0] _T_26880; // @[Switch.scala 34:32:@7725.4]
  wire [31:0] _T_26889; // @[Switch.scala 34:32:@7734.4]
  wire [63:0] _T_26890; // @[Switch.scala 34:32:@7735.4]
  wire  _T_26894; // @[Switch.scala 30:53:@7738.4]
  wire  valid_24_0; // @[Switch.scala 30:36:@7739.4]
  wire  _T_26897; // @[Switch.scala 30:53:@7741.4]
  wire  valid_24_1; // @[Switch.scala 30:36:@7742.4]
  wire  _T_26900; // @[Switch.scala 30:53:@7744.4]
  wire  valid_24_2; // @[Switch.scala 30:36:@7745.4]
  wire  _T_26903; // @[Switch.scala 30:53:@7747.4]
  wire  valid_24_3; // @[Switch.scala 30:36:@7748.4]
  wire  _T_26906; // @[Switch.scala 30:53:@7750.4]
  wire  valid_24_4; // @[Switch.scala 30:36:@7751.4]
  wire  _T_26909; // @[Switch.scala 30:53:@7753.4]
  wire  valid_24_5; // @[Switch.scala 30:36:@7754.4]
  wire  _T_26912; // @[Switch.scala 30:53:@7756.4]
  wire  valid_24_6; // @[Switch.scala 30:36:@7757.4]
  wire  _T_26915; // @[Switch.scala 30:53:@7759.4]
  wire  valid_24_7; // @[Switch.scala 30:36:@7760.4]
  wire  _T_26918; // @[Switch.scala 30:53:@7762.4]
  wire  valid_24_8; // @[Switch.scala 30:36:@7763.4]
  wire  _T_26921; // @[Switch.scala 30:53:@7765.4]
  wire  valid_24_9; // @[Switch.scala 30:36:@7766.4]
  wire  _T_26924; // @[Switch.scala 30:53:@7768.4]
  wire  valid_24_10; // @[Switch.scala 30:36:@7769.4]
  wire  _T_26927; // @[Switch.scala 30:53:@7771.4]
  wire  valid_24_11; // @[Switch.scala 30:36:@7772.4]
  wire  _T_26930; // @[Switch.scala 30:53:@7774.4]
  wire  valid_24_12; // @[Switch.scala 30:36:@7775.4]
  wire  _T_26933; // @[Switch.scala 30:53:@7777.4]
  wire  valid_24_13; // @[Switch.scala 30:36:@7778.4]
  wire  _T_26936; // @[Switch.scala 30:53:@7780.4]
  wire  valid_24_14; // @[Switch.scala 30:36:@7781.4]
  wire  _T_26939; // @[Switch.scala 30:53:@7783.4]
  wire  valid_24_15; // @[Switch.scala 30:36:@7784.4]
  wire  _T_26942; // @[Switch.scala 30:53:@7786.4]
  wire  valid_24_16; // @[Switch.scala 30:36:@7787.4]
  wire  _T_26945; // @[Switch.scala 30:53:@7789.4]
  wire  valid_24_17; // @[Switch.scala 30:36:@7790.4]
  wire  _T_26948; // @[Switch.scala 30:53:@7792.4]
  wire  valid_24_18; // @[Switch.scala 30:36:@7793.4]
  wire  _T_26951; // @[Switch.scala 30:53:@7795.4]
  wire  valid_24_19; // @[Switch.scala 30:36:@7796.4]
  wire  _T_26954; // @[Switch.scala 30:53:@7798.4]
  wire  valid_24_20; // @[Switch.scala 30:36:@7799.4]
  wire  _T_26957; // @[Switch.scala 30:53:@7801.4]
  wire  valid_24_21; // @[Switch.scala 30:36:@7802.4]
  wire  _T_26960; // @[Switch.scala 30:53:@7804.4]
  wire  valid_24_22; // @[Switch.scala 30:36:@7805.4]
  wire  _T_26963; // @[Switch.scala 30:53:@7807.4]
  wire  valid_24_23; // @[Switch.scala 30:36:@7808.4]
  wire  _T_26966; // @[Switch.scala 30:53:@7810.4]
  wire  valid_24_24; // @[Switch.scala 30:36:@7811.4]
  wire  _T_26969; // @[Switch.scala 30:53:@7813.4]
  wire  valid_24_25; // @[Switch.scala 30:36:@7814.4]
  wire  _T_26972; // @[Switch.scala 30:53:@7816.4]
  wire  valid_24_26; // @[Switch.scala 30:36:@7817.4]
  wire  _T_26975; // @[Switch.scala 30:53:@7819.4]
  wire  valid_24_27; // @[Switch.scala 30:36:@7820.4]
  wire  _T_26978; // @[Switch.scala 30:53:@7822.4]
  wire  valid_24_28; // @[Switch.scala 30:36:@7823.4]
  wire  _T_26981; // @[Switch.scala 30:53:@7825.4]
  wire  valid_24_29; // @[Switch.scala 30:36:@7826.4]
  wire  _T_26984; // @[Switch.scala 30:53:@7828.4]
  wire  valid_24_30; // @[Switch.scala 30:36:@7829.4]
  wire  _T_26987; // @[Switch.scala 30:53:@7831.4]
  wire  valid_24_31; // @[Switch.scala 30:36:@7832.4]
  wire  _T_26990; // @[Switch.scala 30:53:@7834.4]
  wire  valid_24_32; // @[Switch.scala 30:36:@7835.4]
  wire  _T_26993; // @[Switch.scala 30:53:@7837.4]
  wire  valid_24_33; // @[Switch.scala 30:36:@7838.4]
  wire  _T_26996; // @[Switch.scala 30:53:@7840.4]
  wire  valid_24_34; // @[Switch.scala 30:36:@7841.4]
  wire  _T_26999; // @[Switch.scala 30:53:@7843.4]
  wire  valid_24_35; // @[Switch.scala 30:36:@7844.4]
  wire  _T_27002; // @[Switch.scala 30:53:@7846.4]
  wire  valid_24_36; // @[Switch.scala 30:36:@7847.4]
  wire  _T_27005; // @[Switch.scala 30:53:@7849.4]
  wire  valid_24_37; // @[Switch.scala 30:36:@7850.4]
  wire  _T_27008; // @[Switch.scala 30:53:@7852.4]
  wire  valid_24_38; // @[Switch.scala 30:36:@7853.4]
  wire  _T_27011; // @[Switch.scala 30:53:@7855.4]
  wire  valid_24_39; // @[Switch.scala 30:36:@7856.4]
  wire  _T_27014; // @[Switch.scala 30:53:@7858.4]
  wire  valid_24_40; // @[Switch.scala 30:36:@7859.4]
  wire  _T_27017; // @[Switch.scala 30:53:@7861.4]
  wire  valid_24_41; // @[Switch.scala 30:36:@7862.4]
  wire  _T_27020; // @[Switch.scala 30:53:@7864.4]
  wire  valid_24_42; // @[Switch.scala 30:36:@7865.4]
  wire  _T_27023; // @[Switch.scala 30:53:@7867.4]
  wire  valid_24_43; // @[Switch.scala 30:36:@7868.4]
  wire  _T_27026; // @[Switch.scala 30:53:@7870.4]
  wire  valid_24_44; // @[Switch.scala 30:36:@7871.4]
  wire  _T_27029; // @[Switch.scala 30:53:@7873.4]
  wire  valid_24_45; // @[Switch.scala 30:36:@7874.4]
  wire  _T_27032; // @[Switch.scala 30:53:@7876.4]
  wire  valid_24_46; // @[Switch.scala 30:36:@7877.4]
  wire  _T_27035; // @[Switch.scala 30:53:@7879.4]
  wire  valid_24_47; // @[Switch.scala 30:36:@7880.4]
  wire  _T_27038; // @[Switch.scala 30:53:@7882.4]
  wire  valid_24_48; // @[Switch.scala 30:36:@7883.4]
  wire  _T_27041; // @[Switch.scala 30:53:@7885.4]
  wire  valid_24_49; // @[Switch.scala 30:36:@7886.4]
  wire  _T_27044; // @[Switch.scala 30:53:@7888.4]
  wire  valid_24_50; // @[Switch.scala 30:36:@7889.4]
  wire  _T_27047; // @[Switch.scala 30:53:@7891.4]
  wire  valid_24_51; // @[Switch.scala 30:36:@7892.4]
  wire  _T_27050; // @[Switch.scala 30:53:@7894.4]
  wire  valid_24_52; // @[Switch.scala 30:36:@7895.4]
  wire  _T_27053; // @[Switch.scala 30:53:@7897.4]
  wire  valid_24_53; // @[Switch.scala 30:36:@7898.4]
  wire  _T_27056; // @[Switch.scala 30:53:@7900.4]
  wire  valid_24_54; // @[Switch.scala 30:36:@7901.4]
  wire  _T_27059; // @[Switch.scala 30:53:@7903.4]
  wire  valid_24_55; // @[Switch.scala 30:36:@7904.4]
  wire  _T_27062; // @[Switch.scala 30:53:@7906.4]
  wire  valid_24_56; // @[Switch.scala 30:36:@7907.4]
  wire  _T_27065; // @[Switch.scala 30:53:@7909.4]
  wire  valid_24_57; // @[Switch.scala 30:36:@7910.4]
  wire  _T_27068; // @[Switch.scala 30:53:@7912.4]
  wire  valid_24_58; // @[Switch.scala 30:36:@7913.4]
  wire  _T_27071; // @[Switch.scala 30:53:@7915.4]
  wire  valid_24_59; // @[Switch.scala 30:36:@7916.4]
  wire  _T_27074; // @[Switch.scala 30:53:@7918.4]
  wire  valid_24_60; // @[Switch.scala 30:36:@7919.4]
  wire  _T_27077; // @[Switch.scala 30:53:@7921.4]
  wire  valid_24_61; // @[Switch.scala 30:36:@7922.4]
  wire  _T_27080; // @[Switch.scala 30:53:@7924.4]
  wire  valid_24_62; // @[Switch.scala 30:36:@7925.4]
  wire  _T_27083; // @[Switch.scala 30:53:@7927.4]
  wire  valid_24_63; // @[Switch.scala 30:36:@7928.4]
  wire [5:0] _T_27149; // @[Mux.scala 31:69:@7930.4]
  wire [5:0] _T_27150; // @[Mux.scala 31:69:@7931.4]
  wire [5:0] _T_27151; // @[Mux.scala 31:69:@7932.4]
  wire [5:0] _T_27152; // @[Mux.scala 31:69:@7933.4]
  wire [5:0] _T_27153; // @[Mux.scala 31:69:@7934.4]
  wire [5:0] _T_27154; // @[Mux.scala 31:69:@7935.4]
  wire [5:0] _T_27155; // @[Mux.scala 31:69:@7936.4]
  wire [5:0] _T_27156; // @[Mux.scala 31:69:@7937.4]
  wire [5:0] _T_27157; // @[Mux.scala 31:69:@7938.4]
  wire [5:0] _T_27158; // @[Mux.scala 31:69:@7939.4]
  wire [5:0] _T_27159; // @[Mux.scala 31:69:@7940.4]
  wire [5:0] _T_27160; // @[Mux.scala 31:69:@7941.4]
  wire [5:0] _T_27161; // @[Mux.scala 31:69:@7942.4]
  wire [5:0] _T_27162; // @[Mux.scala 31:69:@7943.4]
  wire [5:0] _T_27163; // @[Mux.scala 31:69:@7944.4]
  wire [5:0] _T_27164; // @[Mux.scala 31:69:@7945.4]
  wire [5:0] _T_27165; // @[Mux.scala 31:69:@7946.4]
  wire [5:0] _T_27166; // @[Mux.scala 31:69:@7947.4]
  wire [5:0] _T_27167; // @[Mux.scala 31:69:@7948.4]
  wire [5:0] _T_27168; // @[Mux.scala 31:69:@7949.4]
  wire [5:0] _T_27169; // @[Mux.scala 31:69:@7950.4]
  wire [5:0] _T_27170; // @[Mux.scala 31:69:@7951.4]
  wire [5:0] _T_27171; // @[Mux.scala 31:69:@7952.4]
  wire [5:0] _T_27172; // @[Mux.scala 31:69:@7953.4]
  wire [5:0] _T_27173; // @[Mux.scala 31:69:@7954.4]
  wire [5:0] _T_27174; // @[Mux.scala 31:69:@7955.4]
  wire [5:0] _T_27175; // @[Mux.scala 31:69:@7956.4]
  wire [5:0] _T_27176; // @[Mux.scala 31:69:@7957.4]
  wire [5:0] _T_27177; // @[Mux.scala 31:69:@7958.4]
  wire [5:0] _T_27178; // @[Mux.scala 31:69:@7959.4]
  wire [5:0] _T_27179; // @[Mux.scala 31:69:@7960.4]
  wire [5:0] _T_27180; // @[Mux.scala 31:69:@7961.4]
  wire [5:0] _T_27181; // @[Mux.scala 31:69:@7962.4]
  wire [5:0] _T_27182; // @[Mux.scala 31:69:@7963.4]
  wire [5:0] _T_27183; // @[Mux.scala 31:69:@7964.4]
  wire [5:0] _T_27184; // @[Mux.scala 31:69:@7965.4]
  wire [5:0] _T_27185; // @[Mux.scala 31:69:@7966.4]
  wire [5:0] _T_27186; // @[Mux.scala 31:69:@7967.4]
  wire [5:0] _T_27187; // @[Mux.scala 31:69:@7968.4]
  wire [5:0] _T_27188; // @[Mux.scala 31:69:@7969.4]
  wire [5:0] _T_27189; // @[Mux.scala 31:69:@7970.4]
  wire [5:0] _T_27190; // @[Mux.scala 31:69:@7971.4]
  wire [5:0] _T_27191; // @[Mux.scala 31:69:@7972.4]
  wire [5:0] _T_27192; // @[Mux.scala 31:69:@7973.4]
  wire [5:0] _T_27193; // @[Mux.scala 31:69:@7974.4]
  wire [5:0] _T_27194; // @[Mux.scala 31:69:@7975.4]
  wire [5:0] _T_27195; // @[Mux.scala 31:69:@7976.4]
  wire [5:0] _T_27196; // @[Mux.scala 31:69:@7977.4]
  wire [5:0] _T_27197; // @[Mux.scala 31:69:@7978.4]
  wire [5:0] _T_27198; // @[Mux.scala 31:69:@7979.4]
  wire [5:0] _T_27199; // @[Mux.scala 31:69:@7980.4]
  wire [5:0] _T_27200; // @[Mux.scala 31:69:@7981.4]
  wire [5:0] _T_27201; // @[Mux.scala 31:69:@7982.4]
  wire [5:0] _T_27202; // @[Mux.scala 31:69:@7983.4]
  wire [5:0] _T_27203; // @[Mux.scala 31:69:@7984.4]
  wire [5:0] _T_27204; // @[Mux.scala 31:69:@7985.4]
  wire [5:0] _T_27205; // @[Mux.scala 31:69:@7986.4]
  wire [5:0] _T_27206; // @[Mux.scala 31:69:@7987.4]
  wire [5:0] _T_27207; // @[Mux.scala 31:69:@7988.4]
  wire [5:0] _T_27208; // @[Mux.scala 31:69:@7989.4]
  wire [5:0] _T_27209; // @[Mux.scala 31:69:@7990.4]
  wire [5:0] _T_27210; // @[Mux.scala 31:69:@7991.4]
  wire [5:0] select_24; // @[Mux.scala 31:69:@7992.4]
  wire [47:0] _GEN_1537; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1538; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1539; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1540; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1541; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1542; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1543; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1544; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1545; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1546; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1547; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1548; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1549; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1550; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1551; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1552; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1553; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1554; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1555; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1556; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1557; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1558; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1559; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1560; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1561; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1562; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1563; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1564; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1565; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1566; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1567; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1568; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1569; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1570; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1571; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1572; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1573; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1574; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1575; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1576; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1577; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1578; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1579; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1580; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1581; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1582; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1583; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1584; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1585; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1586; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1587; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1588; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1589; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1590; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1591; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1592; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1593; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1594; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1595; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1596; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1597; // @[Switch.scala 33:19:@7994.4]
  wire [47:0] _GEN_1598; // @[Switch.scala 33:19:@7994.4]
  wire [7:0] _T_27219; // @[Switch.scala 34:32:@8001.4]
  wire [15:0] _T_27227; // @[Switch.scala 34:32:@8009.4]
  wire [7:0] _T_27234; // @[Switch.scala 34:32:@8016.4]
  wire [31:0] _T_27243; // @[Switch.scala 34:32:@8025.4]
  wire [7:0] _T_27250; // @[Switch.scala 34:32:@8032.4]
  wire [15:0] _T_27258; // @[Switch.scala 34:32:@8040.4]
  wire [7:0] _T_27265; // @[Switch.scala 34:32:@8047.4]
  wire [31:0] _T_27274; // @[Switch.scala 34:32:@8056.4]
  wire [63:0] _T_27275; // @[Switch.scala 34:32:@8057.4]
  wire  _T_27279; // @[Switch.scala 30:53:@8060.4]
  wire  valid_25_0; // @[Switch.scala 30:36:@8061.4]
  wire  _T_27282; // @[Switch.scala 30:53:@8063.4]
  wire  valid_25_1; // @[Switch.scala 30:36:@8064.4]
  wire  _T_27285; // @[Switch.scala 30:53:@8066.4]
  wire  valid_25_2; // @[Switch.scala 30:36:@8067.4]
  wire  _T_27288; // @[Switch.scala 30:53:@8069.4]
  wire  valid_25_3; // @[Switch.scala 30:36:@8070.4]
  wire  _T_27291; // @[Switch.scala 30:53:@8072.4]
  wire  valid_25_4; // @[Switch.scala 30:36:@8073.4]
  wire  _T_27294; // @[Switch.scala 30:53:@8075.4]
  wire  valid_25_5; // @[Switch.scala 30:36:@8076.4]
  wire  _T_27297; // @[Switch.scala 30:53:@8078.4]
  wire  valid_25_6; // @[Switch.scala 30:36:@8079.4]
  wire  _T_27300; // @[Switch.scala 30:53:@8081.4]
  wire  valid_25_7; // @[Switch.scala 30:36:@8082.4]
  wire  _T_27303; // @[Switch.scala 30:53:@8084.4]
  wire  valid_25_8; // @[Switch.scala 30:36:@8085.4]
  wire  _T_27306; // @[Switch.scala 30:53:@8087.4]
  wire  valid_25_9; // @[Switch.scala 30:36:@8088.4]
  wire  _T_27309; // @[Switch.scala 30:53:@8090.4]
  wire  valid_25_10; // @[Switch.scala 30:36:@8091.4]
  wire  _T_27312; // @[Switch.scala 30:53:@8093.4]
  wire  valid_25_11; // @[Switch.scala 30:36:@8094.4]
  wire  _T_27315; // @[Switch.scala 30:53:@8096.4]
  wire  valid_25_12; // @[Switch.scala 30:36:@8097.4]
  wire  _T_27318; // @[Switch.scala 30:53:@8099.4]
  wire  valid_25_13; // @[Switch.scala 30:36:@8100.4]
  wire  _T_27321; // @[Switch.scala 30:53:@8102.4]
  wire  valid_25_14; // @[Switch.scala 30:36:@8103.4]
  wire  _T_27324; // @[Switch.scala 30:53:@8105.4]
  wire  valid_25_15; // @[Switch.scala 30:36:@8106.4]
  wire  _T_27327; // @[Switch.scala 30:53:@8108.4]
  wire  valid_25_16; // @[Switch.scala 30:36:@8109.4]
  wire  _T_27330; // @[Switch.scala 30:53:@8111.4]
  wire  valid_25_17; // @[Switch.scala 30:36:@8112.4]
  wire  _T_27333; // @[Switch.scala 30:53:@8114.4]
  wire  valid_25_18; // @[Switch.scala 30:36:@8115.4]
  wire  _T_27336; // @[Switch.scala 30:53:@8117.4]
  wire  valid_25_19; // @[Switch.scala 30:36:@8118.4]
  wire  _T_27339; // @[Switch.scala 30:53:@8120.4]
  wire  valid_25_20; // @[Switch.scala 30:36:@8121.4]
  wire  _T_27342; // @[Switch.scala 30:53:@8123.4]
  wire  valid_25_21; // @[Switch.scala 30:36:@8124.4]
  wire  _T_27345; // @[Switch.scala 30:53:@8126.4]
  wire  valid_25_22; // @[Switch.scala 30:36:@8127.4]
  wire  _T_27348; // @[Switch.scala 30:53:@8129.4]
  wire  valid_25_23; // @[Switch.scala 30:36:@8130.4]
  wire  _T_27351; // @[Switch.scala 30:53:@8132.4]
  wire  valid_25_24; // @[Switch.scala 30:36:@8133.4]
  wire  _T_27354; // @[Switch.scala 30:53:@8135.4]
  wire  valid_25_25; // @[Switch.scala 30:36:@8136.4]
  wire  _T_27357; // @[Switch.scala 30:53:@8138.4]
  wire  valid_25_26; // @[Switch.scala 30:36:@8139.4]
  wire  _T_27360; // @[Switch.scala 30:53:@8141.4]
  wire  valid_25_27; // @[Switch.scala 30:36:@8142.4]
  wire  _T_27363; // @[Switch.scala 30:53:@8144.4]
  wire  valid_25_28; // @[Switch.scala 30:36:@8145.4]
  wire  _T_27366; // @[Switch.scala 30:53:@8147.4]
  wire  valid_25_29; // @[Switch.scala 30:36:@8148.4]
  wire  _T_27369; // @[Switch.scala 30:53:@8150.4]
  wire  valid_25_30; // @[Switch.scala 30:36:@8151.4]
  wire  _T_27372; // @[Switch.scala 30:53:@8153.4]
  wire  valid_25_31; // @[Switch.scala 30:36:@8154.4]
  wire  _T_27375; // @[Switch.scala 30:53:@8156.4]
  wire  valid_25_32; // @[Switch.scala 30:36:@8157.4]
  wire  _T_27378; // @[Switch.scala 30:53:@8159.4]
  wire  valid_25_33; // @[Switch.scala 30:36:@8160.4]
  wire  _T_27381; // @[Switch.scala 30:53:@8162.4]
  wire  valid_25_34; // @[Switch.scala 30:36:@8163.4]
  wire  _T_27384; // @[Switch.scala 30:53:@8165.4]
  wire  valid_25_35; // @[Switch.scala 30:36:@8166.4]
  wire  _T_27387; // @[Switch.scala 30:53:@8168.4]
  wire  valid_25_36; // @[Switch.scala 30:36:@8169.4]
  wire  _T_27390; // @[Switch.scala 30:53:@8171.4]
  wire  valid_25_37; // @[Switch.scala 30:36:@8172.4]
  wire  _T_27393; // @[Switch.scala 30:53:@8174.4]
  wire  valid_25_38; // @[Switch.scala 30:36:@8175.4]
  wire  _T_27396; // @[Switch.scala 30:53:@8177.4]
  wire  valid_25_39; // @[Switch.scala 30:36:@8178.4]
  wire  _T_27399; // @[Switch.scala 30:53:@8180.4]
  wire  valid_25_40; // @[Switch.scala 30:36:@8181.4]
  wire  _T_27402; // @[Switch.scala 30:53:@8183.4]
  wire  valid_25_41; // @[Switch.scala 30:36:@8184.4]
  wire  _T_27405; // @[Switch.scala 30:53:@8186.4]
  wire  valid_25_42; // @[Switch.scala 30:36:@8187.4]
  wire  _T_27408; // @[Switch.scala 30:53:@8189.4]
  wire  valid_25_43; // @[Switch.scala 30:36:@8190.4]
  wire  _T_27411; // @[Switch.scala 30:53:@8192.4]
  wire  valid_25_44; // @[Switch.scala 30:36:@8193.4]
  wire  _T_27414; // @[Switch.scala 30:53:@8195.4]
  wire  valid_25_45; // @[Switch.scala 30:36:@8196.4]
  wire  _T_27417; // @[Switch.scala 30:53:@8198.4]
  wire  valid_25_46; // @[Switch.scala 30:36:@8199.4]
  wire  _T_27420; // @[Switch.scala 30:53:@8201.4]
  wire  valid_25_47; // @[Switch.scala 30:36:@8202.4]
  wire  _T_27423; // @[Switch.scala 30:53:@8204.4]
  wire  valid_25_48; // @[Switch.scala 30:36:@8205.4]
  wire  _T_27426; // @[Switch.scala 30:53:@8207.4]
  wire  valid_25_49; // @[Switch.scala 30:36:@8208.4]
  wire  _T_27429; // @[Switch.scala 30:53:@8210.4]
  wire  valid_25_50; // @[Switch.scala 30:36:@8211.4]
  wire  _T_27432; // @[Switch.scala 30:53:@8213.4]
  wire  valid_25_51; // @[Switch.scala 30:36:@8214.4]
  wire  _T_27435; // @[Switch.scala 30:53:@8216.4]
  wire  valid_25_52; // @[Switch.scala 30:36:@8217.4]
  wire  _T_27438; // @[Switch.scala 30:53:@8219.4]
  wire  valid_25_53; // @[Switch.scala 30:36:@8220.4]
  wire  _T_27441; // @[Switch.scala 30:53:@8222.4]
  wire  valid_25_54; // @[Switch.scala 30:36:@8223.4]
  wire  _T_27444; // @[Switch.scala 30:53:@8225.4]
  wire  valid_25_55; // @[Switch.scala 30:36:@8226.4]
  wire  _T_27447; // @[Switch.scala 30:53:@8228.4]
  wire  valid_25_56; // @[Switch.scala 30:36:@8229.4]
  wire  _T_27450; // @[Switch.scala 30:53:@8231.4]
  wire  valid_25_57; // @[Switch.scala 30:36:@8232.4]
  wire  _T_27453; // @[Switch.scala 30:53:@8234.4]
  wire  valid_25_58; // @[Switch.scala 30:36:@8235.4]
  wire  _T_27456; // @[Switch.scala 30:53:@8237.4]
  wire  valid_25_59; // @[Switch.scala 30:36:@8238.4]
  wire  _T_27459; // @[Switch.scala 30:53:@8240.4]
  wire  valid_25_60; // @[Switch.scala 30:36:@8241.4]
  wire  _T_27462; // @[Switch.scala 30:53:@8243.4]
  wire  valid_25_61; // @[Switch.scala 30:36:@8244.4]
  wire  _T_27465; // @[Switch.scala 30:53:@8246.4]
  wire  valid_25_62; // @[Switch.scala 30:36:@8247.4]
  wire  _T_27468; // @[Switch.scala 30:53:@8249.4]
  wire  valid_25_63; // @[Switch.scala 30:36:@8250.4]
  wire [5:0] _T_27534; // @[Mux.scala 31:69:@8252.4]
  wire [5:0] _T_27535; // @[Mux.scala 31:69:@8253.4]
  wire [5:0] _T_27536; // @[Mux.scala 31:69:@8254.4]
  wire [5:0] _T_27537; // @[Mux.scala 31:69:@8255.4]
  wire [5:0] _T_27538; // @[Mux.scala 31:69:@8256.4]
  wire [5:0] _T_27539; // @[Mux.scala 31:69:@8257.4]
  wire [5:0] _T_27540; // @[Mux.scala 31:69:@8258.4]
  wire [5:0] _T_27541; // @[Mux.scala 31:69:@8259.4]
  wire [5:0] _T_27542; // @[Mux.scala 31:69:@8260.4]
  wire [5:0] _T_27543; // @[Mux.scala 31:69:@8261.4]
  wire [5:0] _T_27544; // @[Mux.scala 31:69:@8262.4]
  wire [5:0] _T_27545; // @[Mux.scala 31:69:@8263.4]
  wire [5:0] _T_27546; // @[Mux.scala 31:69:@8264.4]
  wire [5:0] _T_27547; // @[Mux.scala 31:69:@8265.4]
  wire [5:0] _T_27548; // @[Mux.scala 31:69:@8266.4]
  wire [5:0] _T_27549; // @[Mux.scala 31:69:@8267.4]
  wire [5:0] _T_27550; // @[Mux.scala 31:69:@8268.4]
  wire [5:0] _T_27551; // @[Mux.scala 31:69:@8269.4]
  wire [5:0] _T_27552; // @[Mux.scala 31:69:@8270.4]
  wire [5:0] _T_27553; // @[Mux.scala 31:69:@8271.4]
  wire [5:0] _T_27554; // @[Mux.scala 31:69:@8272.4]
  wire [5:0] _T_27555; // @[Mux.scala 31:69:@8273.4]
  wire [5:0] _T_27556; // @[Mux.scala 31:69:@8274.4]
  wire [5:0] _T_27557; // @[Mux.scala 31:69:@8275.4]
  wire [5:0] _T_27558; // @[Mux.scala 31:69:@8276.4]
  wire [5:0] _T_27559; // @[Mux.scala 31:69:@8277.4]
  wire [5:0] _T_27560; // @[Mux.scala 31:69:@8278.4]
  wire [5:0] _T_27561; // @[Mux.scala 31:69:@8279.4]
  wire [5:0] _T_27562; // @[Mux.scala 31:69:@8280.4]
  wire [5:0] _T_27563; // @[Mux.scala 31:69:@8281.4]
  wire [5:0] _T_27564; // @[Mux.scala 31:69:@8282.4]
  wire [5:0] _T_27565; // @[Mux.scala 31:69:@8283.4]
  wire [5:0] _T_27566; // @[Mux.scala 31:69:@8284.4]
  wire [5:0] _T_27567; // @[Mux.scala 31:69:@8285.4]
  wire [5:0] _T_27568; // @[Mux.scala 31:69:@8286.4]
  wire [5:0] _T_27569; // @[Mux.scala 31:69:@8287.4]
  wire [5:0] _T_27570; // @[Mux.scala 31:69:@8288.4]
  wire [5:0] _T_27571; // @[Mux.scala 31:69:@8289.4]
  wire [5:0] _T_27572; // @[Mux.scala 31:69:@8290.4]
  wire [5:0] _T_27573; // @[Mux.scala 31:69:@8291.4]
  wire [5:0] _T_27574; // @[Mux.scala 31:69:@8292.4]
  wire [5:0] _T_27575; // @[Mux.scala 31:69:@8293.4]
  wire [5:0] _T_27576; // @[Mux.scala 31:69:@8294.4]
  wire [5:0] _T_27577; // @[Mux.scala 31:69:@8295.4]
  wire [5:0] _T_27578; // @[Mux.scala 31:69:@8296.4]
  wire [5:0] _T_27579; // @[Mux.scala 31:69:@8297.4]
  wire [5:0] _T_27580; // @[Mux.scala 31:69:@8298.4]
  wire [5:0] _T_27581; // @[Mux.scala 31:69:@8299.4]
  wire [5:0] _T_27582; // @[Mux.scala 31:69:@8300.4]
  wire [5:0] _T_27583; // @[Mux.scala 31:69:@8301.4]
  wire [5:0] _T_27584; // @[Mux.scala 31:69:@8302.4]
  wire [5:0] _T_27585; // @[Mux.scala 31:69:@8303.4]
  wire [5:0] _T_27586; // @[Mux.scala 31:69:@8304.4]
  wire [5:0] _T_27587; // @[Mux.scala 31:69:@8305.4]
  wire [5:0] _T_27588; // @[Mux.scala 31:69:@8306.4]
  wire [5:0] _T_27589; // @[Mux.scala 31:69:@8307.4]
  wire [5:0] _T_27590; // @[Mux.scala 31:69:@8308.4]
  wire [5:0] _T_27591; // @[Mux.scala 31:69:@8309.4]
  wire [5:0] _T_27592; // @[Mux.scala 31:69:@8310.4]
  wire [5:0] _T_27593; // @[Mux.scala 31:69:@8311.4]
  wire [5:0] _T_27594; // @[Mux.scala 31:69:@8312.4]
  wire [5:0] _T_27595; // @[Mux.scala 31:69:@8313.4]
  wire [5:0] select_25; // @[Mux.scala 31:69:@8314.4]
  wire [47:0] _GEN_1601; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1602; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1603; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1604; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1605; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1606; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1607; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1608; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1609; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1610; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1611; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1612; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1613; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1614; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1615; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1616; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1617; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1618; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1619; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1620; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1621; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1622; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1623; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1624; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1625; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1626; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1627; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1628; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1629; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1630; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1631; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1632; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1633; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1634; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1635; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1636; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1637; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1638; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1639; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1640; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1641; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1642; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1643; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1644; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1645; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1646; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1647; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1648; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1649; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1650; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1651; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1652; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1653; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1654; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1655; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1656; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1657; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1658; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1659; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1660; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1661; // @[Switch.scala 33:19:@8316.4]
  wire [47:0] _GEN_1662; // @[Switch.scala 33:19:@8316.4]
  wire [7:0] _T_27604; // @[Switch.scala 34:32:@8323.4]
  wire [15:0] _T_27612; // @[Switch.scala 34:32:@8331.4]
  wire [7:0] _T_27619; // @[Switch.scala 34:32:@8338.4]
  wire [31:0] _T_27628; // @[Switch.scala 34:32:@8347.4]
  wire [7:0] _T_27635; // @[Switch.scala 34:32:@8354.4]
  wire [15:0] _T_27643; // @[Switch.scala 34:32:@8362.4]
  wire [7:0] _T_27650; // @[Switch.scala 34:32:@8369.4]
  wire [31:0] _T_27659; // @[Switch.scala 34:32:@8378.4]
  wire [63:0] _T_27660; // @[Switch.scala 34:32:@8379.4]
  wire  _T_27664; // @[Switch.scala 30:53:@8382.4]
  wire  valid_26_0; // @[Switch.scala 30:36:@8383.4]
  wire  _T_27667; // @[Switch.scala 30:53:@8385.4]
  wire  valid_26_1; // @[Switch.scala 30:36:@8386.4]
  wire  _T_27670; // @[Switch.scala 30:53:@8388.4]
  wire  valid_26_2; // @[Switch.scala 30:36:@8389.4]
  wire  _T_27673; // @[Switch.scala 30:53:@8391.4]
  wire  valid_26_3; // @[Switch.scala 30:36:@8392.4]
  wire  _T_27676; // @[Switch.scala 30:53:@8394.4]
  wire  valid_26_4; // @[Switch.scala 30:36:@8395.4]
  wire  _T_27679; // @[Switch.scala 30:53:@8397.4]
  wire  valid_26_5; // @[Switch.scala 30:36:@8398.4]
  wire  _T_27682; // @[Switch.scala 30:53:@8400.4]
  wire  valid_26_6; // @[Switch.scala 30:36:@8401.4]
  wire  _T_27685; // @[Switch.scala 30:53:@8403.4]
  wire  valid_26_7; // @[Switch.scala 30:36:@8404.4]
  wire  _T_27688; // @[Switch.scala 30:53:@8406.4]
  wire  valid_26_8; // @[Switch.scala 30:36:@8407.4]
  wire  _T_27691; // @[Switch.scala 30:53:@8409.4]
  wire  valid_26_9; // @[Switch.scala 30:36:@8410.4]
  wire  _T_27694; // @[Switch.scala 30:53:@8412.4]
  wire  valid_26_10; // @[Switch.scala 30:36:@8413.4]
  wire  _T_27697; // @[Switch.scala 30:53:@8415.4]
  wire  valid_26_11; // @[Switch.scala 30:36:@8416.4]
  wire  _T_27700; // @[Switch.scala 30:53:@8418.4]
  wire  valid_26_12; // @[Switch.scala 30:36:@8419.4]
  wire  _T_27703; // @[Switch.scala 30:53:@8421.4]
  wire  valid_26_13; // @[Switch.scala 30:36:@8422.4]
  wire  _T_27706; // @[Switch.scala 30:53:@8424.4]
  wire  valid_26_14; // @[Switch.scala 30:36:@8425.4]
  wire  _T_27709; // @[Switch.scala 30:53:@8427.4]
  wire  valid_26_15; // @[Switch.scala 30:36:@8428.4]
  wire  _T_27712; // @[Switch.scala 30:53:@8430.4]
  wire  valid_26_16; // @[Switch.scala 30:36:@8431.4]
  wire  _T_27715; // @[Switch.scala 30:53:@8433.4]
  wire  valid_26_17; // @[Switch.scala 30:36:@8434.4]
  wire  _T_27718; // @[Switch.scala 30:53:@8436.4]
  wire  valid_26_18; // @[Switch.scala 30:36:@8437.4]
  wire  _T_27721; // @[Switch.scala 30:53:@8439.4]
  wire  valid_26_19; // @[Switch.scala 30:36:@8440.4]
  wire  _T_27724; // @[Switch.scala 30:53:@8442.4]
  wire  valid_26_20; // @[Switch.scala 30:36:@8443.4]
  wire  _T_27727; // @[Switch.scala 30:53:@8445.4]
  wire  valid_26_21; // @[Switch.scala 30:36:@8446.4]
  wire  _T_27730; // @[Switch.scala 30:53:@8448.4]
  wire  valid_26_22; // @[Switch.scala 30:36:@8449.4]
  wire  _T_27733; // @[Switch.scala 30:53:@8451.4]
  wire  valid_26_23; // @[Switch.scala 30:36:@8452.4]
  wire  _T_27736; // @[Switch.scala 30:53:@8454.4]
  wire  valid_26_24; // @[Switch.scala 30:36:@8455.4]
  wire  _T_27739; // @[Switch.scala 30:53:@8457.4]
  wire  valid_26_25; // @[Switch.scala 30:36:@8458.4]
  wire  _T_27742; // @[Switch.scala 30:53:@8460.4]
  wire  valid_26_26; // @[Switch.scala 30:36:@8461.4]
  wire  _T_27745; // @[Switch.scala 30:53:@8463.4]
  wire  valid_26_27; // @[Switch.scala 30:36:@8464.4]
  wire  _T_27748; // @[Switch.scala 30:53:@8466.4]
  wire  valid_26_28; // @[Switch.scala 30:36:@8467.4]
  wire  _T_27751; // @[Switch.scala 30:53:@8469.4]
  wire  valid_26_29; // @[Switch.scala 30:36:@8470.4]
  wire  _T_27754; // @[Switch.scala 30:53:@8472.4]
  wire  valid_26_30; // @[Switch.scala 30:36:@8473.4]
  wire  _T_27757; // @[Switch.scala 30:53:@8475.4]
  wire  valid_26_31; // @[Switch.scala 30:36:@8476.4]
  wire  _T_27760; // @[Switch.scala 30:53:@8478.4]
  wire  valid_26_32; // @[Switch.scala 30:36:@8479.4]
  wire  _T_27763; // @[Switch.scala 30:53:@8481.4]
  wire  valid_26_33; // @[Switch.scala 30:36:@8482.4]
  wire  _T_27766; // @[Switch.scala 30:53:@8484.4]
  wire  valid_26_34; // @[Switch.scala 30:36:@8485.4]
  wire  _T_27769; // @[Switch.scala 30:53:@8487.4]
  wire  valid_26_35; // @[Switch.scala 30:36:@8488.4]
  wire  _T_27772; // @[Switch.scala 30:53:@8490.4]
  wire  valid_26_36; // @[Switch.scala 30:36:@8491.4]
  wire  _T_27775; // @[Switch.scala 30:53:@8493.4]
  wire  valid_26_37; // @[Switch.scala 30:36:@8494.4]
  wire  _T_27778; // @[Switch.scala 30:53:@8496.4]
  wire  valid_26_38; // @[Switch.scala 30:36:@8497.4]
  wire  _T_27781; // @[Switch.scala 30:53:@8499.4]
  wire  valid_26_39; // @[Switch.scala 30:36:@8500.4]
  wire  _T_27784; // @[Switch.scala 30:53:@8502.4]
  wire  valid_26_40; // @[Switch.scala 30:36:@8503.4]
  wire  _T_27787; // @[Switch.scala 30:53:@8505.4]
  wire  valid_26_41; // @[Switch.scala 30:36:@8506.4]
  wire  _T_27790; // @[Switch.scala 30:53:@8508.4]
  wire  valid_26_42; // @[Switch.scala 30:36:@8509.4]
  wire  _T_27793; // @[Switch.scala 30:53:@8511.4]
  wire  valid_26_43; // @[Switch.scala 30:36:@8512.4]
  wire  _T_27796; // @[Switch.scala 30:53:@8514.4]
  wire  valid_26_44; // @[Switch.scala 30:36:@8515.4]
  wire  _T_27799; // @[Switch.scala 30:53:@8517.4]
  wire  valid_26_45; // @[Switch.scala 30:36:@8518.4]
  wire  _T_27802; // @[Switch.scala 30:53:@8520.4]
  wire  valid_26_46; // @[Switch.scala 30:36:@8521.4]
  wire  _T_27805; // @[Switch.scala 30:53:@8523.4]
  wire  valid_26_47; // @[Switch.scala 30:36:@8524.4]
  wire  _T_27808; // @[Switch.scala 30:53:@8526.4]
  wire  valid_26_48; // @[Switch.scala 30:36:@8527.4]
  wire  _T_27811; // @[Switch.scala 30:53:@8529.4]
  wire  valid_26_49; // @[Switch.scala 30:36:@8530.4]
  wire  _T_27814; // @[Switch.scala 30:53:@8532.4]
  wire  valid_26_50; // @[Switch.scala 30:36:@8533.4]
  wire  _T_27817; // @[Switch.scala 30:53:@8535.4]
  wire  valid_26_51; // @[Switch.scala 30:36:@8536.4]
  wire  _T_27820; // @[Switch.scala 30:53:@8538.4]
  wire  valid_26_52; // @[Switch.scala 30:36:@8539.4]
  wire  _T_27823; // @[Switch.scala 30:53:@8541.4]
  wire  valid_26_53; // @[Switch.scala 30:36:@8542.4]
  wire  _T_27826; // @[Switch.scala 30:53:@8544.4]
  wire  valid_26_54; // @[Switch.scala 30:36:@8545.4]
  wire  _T_27829; // @[Switch.scala 30:53:@8547.4]
  wire  valid_26_55; // @[Switch.scala 30:36:@8548.4]
  wire  _T_27832; // @[Switch.scala 30:53:@8550.4]
  wire  valid_26_56; // @[Switch.scala 30:36:@8551.4]
  wire  _T_27835; // @[Switch.scala 30:53:@8553.4]
  wire  valid_26_57; // @[Switch.scala 30:36:@8554.4]
  wire  _T_27838; // @[Switch.scala 30:53:@8556.4]
  wire  valid_26_58; // @[Switch.scala 30:36:@8557.4]
  wire  _T_27841; // @[Switch.scala 30:53:@8559.4]
  wire  valid_26_59; // @[Switch.scala 30:36:@8560.4]
  wire  _T_27844; // @[Switch.scala 30:53:@8562.4]
  wire  valid_26_60; // @[Switch.scala 30:36:@8563.4]
  wire  _T_27847; // @[Switch.scala 30:53:@8565.4]
  wire  valid_26_61; // @[Switch.scala 30:36:@8566.4]
  wire  _T_27850; // @[Switch.scala 30:53:@8568.4]
  wire  valid_26_62; // @[Switch.scala 30:36:@8569.4]
  wire  _T_27853; // @[Switch.scala 30:53:@8571.4]
  wire  valid_26_63; // @[Switch.scala 30:36:@8572.4]
  wire [5:0] _T_27919; // @[Mux.scala 31:69:@8574.4]
  wire [5:0] _T_27920; // @[Mux.scala 31:69:@8575.4]
  wire [5:0] _T_27921; // @[Mux.scala 31:69:@8576.4]
  wire [5:0] _T_27922; // @[Mux.scala 31:69:@8577.4]
  wire [5:0] _T_27923; // @[Mux.scala 31:69:@8578.4]
  wire [5:0] _T_27924; // @[Mux.scala 31:69:@8579.4]
  wire [5:0] _T_27925; // @[Mux.scala 31:69:@8580.4]
  wire [5:0] _T_27926; // @[Mux.scala 31:69:@8581.4]
  wire [5:0] _T_27927; // @[Mux.scala 31:69:@8582.4]
  wire [5:0] _T_27928; // @[Mux.scala 31:69:@8583.4]
  wire [5:0] _T_27929; // @[Mux.scala 31:69:@8584.4]
  wire [5:0] _T_27930; // @[Mux.scala 31:69:@8585.4]
  wire [5:0] _T_27931; // @[Mux.scala 31:69:@8586.4]
  wire [5:0] _T_27932; // @[Mux.scala 31:69:@8587.4]
  wire [5:0] _T_27933; // @[Mux.scala 31:69:@8588.4]
  wire [5:0] _T_27934; // @[Mux.scala 31:69:@8589.4]
  wire [5:0] _T_27935; // @[Mux.scala 31:69:@8590.4]
  wire [5:0] _T_27936; // @[Mux.scala 31:69:@8591.4]
  wire [5:0] _T_27937; // @[Mux.scala 31:69:@8592.4]
  wire [5:0] _T_27938; // @[Mux.scala 31:69:@8593.4]
  wire [5:0] _T_27939; // @[Mux.scala 31:69:@8594.4]
  wire [5:0] _T_27940; // @[Mux.scala 31:69:@8595.4]
  wire [5:0] _T_27941; // @[Mux.scala 31:69:@8596.4]
  wire [5:0] _T_27942; // @[Mux.scala 31:69:@8597.4]
  wire [5:0] _T_27943; // @[Mux.scala 31:69:@8598.4]
  wire [5:0] _T_27944; // @[Mux.scala 31:69:@8599.4]
  wire [5:0] _T_27945; // @[Mux.scala 31:69:@8600.4]
  wire [5:0] _T_27946; // @[Mux.scala 31:69:@8601.4]
  wire [5:0] _T_27947; // @[Mux.scala 31:69:@8602.4]
  wire [5:0] _T_27948; // @[Mux.scala 31:69:@8603.4]
  wire [5:0] _T_27949; // @[Mux.scala 31:69:@8604.4]
  wire [5:0] _T_27950; // @[Mux.scala 31:69:@8605.4]
  wire [5:0] _T_27951; // @[Mux.scala 31:69:@8606.4]
  wire [5:0] _T_27952; // @[Mux.scala 31:69:@8607.4]
  wire [5:0] _T_27953; // @[Mux.scala 31:69:@8608.4]
  wire [5:0] _T_27954; // @[Mux.scala 31:69:@8609.4]
  wire [5:0] _T_27955; // @[Mux.scala 31:69:@8610.4]
  wire [5:0] _T_27956; // @[Mux.scala 31:69:@8611.4]
  wire [5:0] _T_27957; // @[Mux.scala 31:69:@8612.4]
  wire [5:0] _T_27958; // @[Mux.scala 31:69:@8613.4]
  wire [5:0] _T_27959; // @[Mux.scala 31:69:@8614.4]
  wire [5:0] _T_27960; // @[Mux.scala 31:69:@8615.4]
  wire [5:0] _T_27961; // @[Mux.scala 31:69:@8616.4]
  wire [5:0] _T_27962; // @[Mux.scala 31:69:@8617.4]
  wire [5:0] _T_27963; // @[Mux.scala 31:69:@8618.4]
  wire [5:0] _T_27964; // @[Mux.scala 31:69:@8619.4]
  wire [5:0] _T_27965; // @[Mux.scala 31:69:@8620.4]
  wire [5:0] _T_27966; // @[Mux.scala 31:69:@8621.4]
  wire [5:0] _T_27967; // @[Mux.scala 31:69:@8622.4]
  wire [5:0] _T_27968; // @[Mux.scala 31:69:@8623.4]
  wire [5:0] _T_27969; // @[Mux.scala 31:69:@8624.4]
  wire [5:0] _T_27970; // @[Mux.scala 31:69:@8625.4]
  wire [5:0] _T_27971; // @[Mux.scala 31:69:@8626.4]
  wire [5:0] _T_27972; // @[Mux.scala 31:69:@8627.4]
  wire [5:0] _T_27973; // @[Mux.scala 31:69:@8628.4]
  wire [5:0] _T_27974; // @[Mux.scala 31:69:@8629.4]
  wire [5:0] _T_27975; // @[Mux.scala 31:69:@8630.4]
  wire [5:0] _T_27976; // @[Mux.scala 31:69:@8631.4]
  wire [5:0] _T_27977; // @[Mux.scala 31:69:@8632.4]
  wire [5:0] _T_27978; // @[Mux.scala 31:69:@8633.4]
  wire [5:0] _T_27979; // @[Mux.scala 31:69:@8634.4]
  wire [5:0] _T_27980; // @[Mux.scala 31:69:@8635.4]
  wire [5:0] select_26; // @[Mux.scala 31:69:@8636.4]
  wire [47:0] _GEN_1665; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1666; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1667; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1668; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1669; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1670; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1671; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1672; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1673; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1674; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1675; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1676; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1677; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1678; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1679; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1680; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1681; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1682; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1683; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1684; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1685; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1686; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1687; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1688; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1689; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1690; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1691; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1692; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1693; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1694; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1695; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1696; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1697; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1698; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1699; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1700; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1701; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1702; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1703; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1704; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1705; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1706; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1707; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1708; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1709; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1710; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1711; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1712; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1713; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1714; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1715; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1716; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1717; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1718; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1719; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1720; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1721; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1722; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1723; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1724; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1725; // @[Switch.scala 33:19:@8638.4]
  wire [47:0] _GEN_1726; // @[Switch.scala 33:19:@8638.4]
  wire [7:0] _T_27989; // @[Switch.scala 34:32:@8645.4]
  wire [15:0] _T_27997; // @[Switch.scala 34:32:@8653.4]
  wire [7:0] _T_28004; // @[Switch.scala 34:32:@8660.4]
  wire [31:0] _T_28013; // @[Switch.scala 34:32:@8669.4]
  wire [7:0] _T_28020; // @[Switch.scala 34:32:@8676.4]
  wire [15:0] _T_28028; // @[Switch.scala 34:32:@8684.4]
  wire [7:0] _T_28035; // @[Switch.scala 34:32:@8691.4]
  wire [31:0] _T_28044; // @[Switch.scala 34:32:@8700.4]
  wire [63:0] _T_28045; // @[Switch.scala 34:32:@8701.4]
  wire  _T_28049; // @[Switch.scala 30:53:@8704.4]
  wire  valid_27_0; // @[Switch.scala 30:36:@8705.4]
  wire  _T_28052; // @[Switch.scala 30:53:@8707.4]
  wire  valid_27_1; // @[Switch.scala 30:36:@8708.4]
  wire  _T_28055; // @[Switch.scala 30:53:@8710.4]
  wire  valid_27_2; // @[Switch.scala 30:36:@8711.4]
  wire  _T_28058; // @[Switch.scala 30:53:@8713.4]
  wire  valid_27_3; // @[Switch.scala 30:36:@8714.4]
  wire  _T_28061; // @[Switch.scala 30:53:@8716.4]
  wire  valid_27_4; // @[Switch.scala 30:36:@8717.4]
  wire  _T_28064; // @[Switch.scala 30:53:@8719.4]
  wire  valid_27_5; // @[Switch.scala 30:36:@8720.4]
  wire  _T_28067; // @[Switch.scala 30:53:@8722.4]
  wire  valid_27_6; // @[Switch.scala 30:36:@8723.4]
  wire  _T_28070; // @[Switch.scala 30:53:@8725.4]
  wire  valid_27_7; // @[Switch.scala 30:36:@8726.4]
  wire  _T_28073; // @[Switch.scala 30:53:@8728.4]
  wire  valid_27_8; // @[Switch.scala 30:36:@8729.4]
  wire  _T_28076; // @[Switch.scala 30:53:@8731.4]
  wire  valid_27_9; // @[Switch.scala 30:36:@8732.4]
  wire  _T_28079; // @[Switch.scala 30:53:@8734.4]
  wire  valid_27_10; // @[Switch.scala 30:36:@8735.4]
  wire  _T_28082; // @[Switch.scala 30:53:@8737.4]
  wire  valid_27_11; // @[Switch.scala 30:36:@8738.4]
  wire  _T_28085; // @[Switch.scala 30:53:@8740.4]
  wire  valid_27_12; // @[Switch.scala 30:36:@8741.4]
  wire  _T_28088; // @[Switch.scala 30:53:@8743.4]
  wire  valid_27_13; // @[Switch.scala 30:36:@8744.4]
  wire  _T_28091; // @[Switch.scala 30:53:@8746.4]
  wire  valid_27_14; // @[Switch.scala 30:36:@8747.4]
  wire  _T_28094; // @[Switch.scala 30:53:@8749.4]
  wire  valid_27_15; // @[Switch.scala 30:36:@8750.4]
  wire  _T_28097; // @[Switch.scala 30:53:@8752.4]
  wire  valid_27_16; // @[Switch.scala 30:36:@8753.4]
  wire  _T_28100; // @[Switch.scala 30:53:@8755.4]
  wire  valid_27_17; // @[Switch.scala 30:36:@8756.4]
  wire  _T_28103; // @[Switch.scala 30:53:@8758.4]
  wire  valid_27_18; // @[Switch.scala 30:36:@8759.4]
  wire  _T_28106; // @[Switch.scala 30:53:@8761.4]
  wire  valid_27_19; // @[Switch.scala 30:36:@8762.4]
  wire  _T_28109; // @[Switch.scala 30:53:@8764.4]
  wire  valid_27_20; // @[Switch.scala 30:36:@8765.4]
  wire  _T_28112; // @[Switch.scala 30:53:@8767.4]
  wire  valid_27_21; // @[Switch.scala 30:36:@8768.4]
  wire  _T_28115; // @[Switch.scala 30:53:@8770.4]
  wire  valid_27_22; // @[Switch.scala 30:36:@8771.4]
  wire  _T_28118; // @[Switch.scala 30:53:@8773.4]
  wire  valid_27_23; // @[Switch.scala 30:36:@8774.4]
  wire  _T_28121; // @[Switch.scala 30:53:@8776.4]
  wire  valid_27_24; // @[Switch.scala 30:36:@8777.4]
  wire  _T_28124; // @[Switch.scala 30:53:@8779.4]
  wire  valid_27_25; // @[Switch.scala 30:36:@8780.4]
  wire  _T_28127; // @[Switch.scala 30:53:@8782.4]
  wire  valid_27_26; // @[Switch.scala 30:36:@8783.4]
  wire  _T_28130; // @[Switch.scala 30:53:@8785.4]
  wire  valid_27_27; // @[Switch.scala 30:36:@8786.4]
  wire  _T_28133; // @[Switch.scala 30:53:@8788.4]
  wire  valid_27_28; // @[Switch.scala 30:36:@8789.4]
  wire  _T_28136; // @[Switch.scala 30:53:@8791.4]
  wire  valid_27_29; // @[Switch.scala 30:36:@8792.4]
  wire  _T_28139; // @[Switch.scala 30:53:@8794.4]
  wire  valid_27_30; // @[Switch.scala 30:36:@8795.4]
  wire  _T_28142; // @[Switch.scala 30:53:@8797.4]
  wire  valid_27_31; // @[Switch.scala 30:36:@8798.4]
  wire  _T_28145; // @[Switch.scala 30:53:@8800.4]
  wire  valid_27_32; // @[Switch.scala 30:36:@8801.4]
  wire  _T_28148; // @[Switch.scala 30:53:@8803.4]
  wire  valid_27_33; // @[Switch.scala 30:36:@8804.4]
  wire  _T_28151; // @[Switch.scala 30:53:@8806.4]
  wire  valid_27_34; // @[Switch.scala 30:36:@8807.4]
  wire  _T_28154; // @[Switch.scala 30:53:@8809.4]
  wire  valid_27_35; // @[Switch.scala 30:36:@8810.4]
  wire  _T_28157; // @[Switch.scala 30:53:@8812.4]
  wire  valid_27_36; // @[Switch.scala 30:36:@8813.4]
  wire  _T_28160; // @[Switch.scala 30:53:@8815.4]
  wire  valid_27_37; // @[Switch.scala 30:36:@8816.4]
  wire  _T_28163; // @[Switch.scala 30:53:@8818.4]
  wire  valid_27_38; // @[Switch.scala 30:36:@8819.4]
  wire  _T_28166; // @[Switch.scala 30:53:@8821.4]
  wire  valid_27_39; // @[Switch.scala 30:36:@8822.4]
  wire  _T_28169; // @[Switch.scala 30:53:@8824.4]
  wire  valid_27_40; // @[Switch.scala 30:36:@8825.4]
  wire  _T_28172; // @[Switch.scala 30:53:@8827.4]
  wire  valid_27_41; // @[Switch.scala 30:36:@8828.4]
  wire  _T_28175; // @[Switch.scala 30:53:@8830.4]
  wire  valid_27_42; // @[Switch.scala 30:36:@8831.4]
  wire  _T_28178; // @[Switch.scala 30:53:@8833.4]
  wire  valid_27_43; // @[Switch.scala 30:36:@8834.4]
  wire  _T_28181; // @[Switch.scala 30:53:@8836.4]
  wire  valid_27_44; // @[Switch.scala 30:36:@8837.4]
  wire  _T_28184; // @[Switch.scala 30:53:@8839.4]
  wire  valid_27_45; // @[Switch.scala 30:36:@8840.4]
  wire  _T_28187; // @[Switch.scala 30:53:@8842.4]
  wire  valid_27_46; // @[Switch.scala 30:36:@8843.4]
  wire  _T_28190; // @[Switch.scala 30:53:@8845.4]
  wire  valid_27_47; // @[Switch.scala 30:36:@8846.4]
  wire  _T_28193; // @[Switch.scala 30:53:@8848.4]
  wire  valid_27_48; // @[Switch.scala 30:36:@8849.4]
  wire  _T_28196; // @[Switch.scala 30:53:@8851.4]
  wire  valid_27_49; // @[Switch.scala 30:36:@8852.4]
  wire  _T_28199; // @[Switch.scala 30:53:@8854.4]
  wire  valid_27_50; // @[Switch.scala 30:36:@8855.4]
  wire  _T_28202; // @[Switch.scala 30:53:@8857.4]
  wire  valid_27_51; // @[Switch.scala 30:36:@8858.4]
  wire  _T_28205; // @[Switch.scala 30:53:@8860.4]
  wire  valid_27_52; // @[Switch.scala 30:36:@8861.4]
  wire  _T_28208; // @[Switch.scala 30:53:@8863.4]
  wire  valid_27_53; // @[Switch.scala 30:36:@8864.4]
  wire  _T_28211; // @[Switch.scala 30:53:@8866.4]
  wire  valid_27_54; // @[Switch.scala 30:36:@8867.4]
  wire  _T_28214; // @[Switch.scala 30:53:@8869.4]
  wire  valid_27_55; // @[Switch.scala 30:36:@8870.4]
  wire  _T_28217; // @[Switch.scala 30:53:@8872.4]
  wire  valid_27_56; // @[Switch.scala 30:36:@8873.4]
  wire  _T_28220; // @[Switch.scala 30:53:@8875.4]
  wire  valid_27_57; // @[Switch.scala 30:36:@8876.4]
  wire  _T_28223; // @[Switch.scala 30:53:@8878.4]
  wire  valid_27_58; // @[Switch.scala 30:36:@8879.4]
  wire  _T_28226; // @[Switch.scala 30:53:@8881.4]
  wire  valid_27_59; // @[Switch.scala 30:36:@8882.4]
  wire  _T_28229; // @[Switch.scala 30:53:@8884.4]
  wire  valid_27_60; // @[Switch.scala 30:36:@8885.4]
  wire  _T_28232; // @[Switch.scala 30:53:@8887.4]
  wire  valid_27_61; // @[Switch.scala 30:36:@8888.4]
  wire  _T_28235; // @[Switch.scala 30:53:@8890.4]
  wire  valid_27_62; // @[Switch.scala 30:36:@8891.4]
  wire  _T_28238; // @[Switch.scala 30:53:@8893.4]
  wire  valid_27_63; // @[Switch.scala 30:36:@8894.4]
  wire [5:0] _T_28304; // @[Mux.scala 31:69:@8896.4]
  wire [5:0] _T_28305; // @[Mux.scala 31:69:@8897.4]
  wire [5:0] _T_28306; // @[Mux.scala 31:69:@8898.4]
  wire [5:0] _T_28307; // @[Mux.scala 31:69:@8899.4]
  wire [5:0] _T_28308; // @[Mux.scala 31:69:@8900.4]
  wire [5:0] _T_28309; // @[Mux.scala 31:69:@8901.4]
  wire [5:0] _T_28310; // @[Mux.scala 31:69:@8902.4]
  wire [5:0] _T_28311; // @[Mux.scala 31:69:@8903.4]
  wire [5:0] _T_28312; // @[Mux.scala 31:69:@8904.4]
  wire [5:0] _T_28313; // @[Mux.scala 31:69:@8905.4]
  wire [5:0] _T_28314; // @[Mux.scala 31:69:@8906.4]
  wire [5:0] _T_28315; // @[Mux.scala 31:69:@8907.4]
  wire [5:0] _T_28316; // @[Mux.scala 31:69:@8908.4]
  wire [5:0] _T_28317; // @[Mux.scala 31:69:@8909.4]
  wire [5:0] _T_28318; // @[Mux.scala 31:69:@8910.4]
  wire [5:0] _T_28319; // @[Mux.scala 31:69:@8911.4]
  wire [5:0] _T_28320; // @[Mux.scala 31:69:@8912.4]
  wire [5:0] _T_28321; // @[Mux.scala 31:69:@8913.4]
  wire [5:0] _T_28322; // @[Mux.scala 31:69:@8914.4]
  wire [5:0] _T_28323; // @[Mux.scala 31:69:@8915.4]
  wire [5:0] _T_28324; // @[Mux.scala 31:69:@8916.4]
  wire [5:0] _T_28325; // @[Mux.scala 31:69:@8917.4]
  wire [5:0] _T_28326; // @[Mux.scala 31:69:@8918.4]
  wire [5:0] _T_28327; // @[Mux.scala 31:69:@8919.4]
  wire [5:0] _T_28328; // @[Mux.scala 31:69:@8920.4]
  wire [5:0] _T_28329; // @[Mux.scala 31:69:@8921.4]
  wire [5:0] _T_28330; // @[Mux.scala 31:69:@8922.4]
  wire [5:0] _T_28331; // @[Mux.scala 31:69:@8923.4]
  wire [5:0] _T_28332; // @[Mux.scala 31:69:@8924.4]
  wire [5:0] _T_28333; // @[Mux.scala 31:69:@8925.4]
  wire [5:0] _T_28334; // @[Mux.scala 31:69:@8926.4]
  wire [5:0] _T_28335; // @[Mux.scala 31:69:@8927.4]
  wire [5:0] _T_28336; // @[Mux.scala 31:69:@8928.4]
  wire [5:0] _T_28337; // @[Mux.scala 31:69:@8929.4]
  wire [5:0] _T_28338; // @[Mux.scala 31:69:@8930.4]
  wire [5:0] _T_28339; // @[Mux.scala 31:69:@8931.4]
  wire [5:0] _T_28340; // @[Mux.scala 31:69:@8932.4]
  wire [5:0] _T_28341; // @[Mux.scala 31:69:@8933.4]
  wire [5:0] _T_28342; // @[Mux.scala 31:69:@8934.4]
  wire [5:0] _T_28343; // @[Mux.scala 31:69:@8935.4]
  wire [5:0] _T_28344; // @[Mux.scala 31:69:@8936.4]
  wire [5:0] _T_28345; // @[Mux.scala 31:69:@8937.4]
  wire [5:0] _T_28346; // @[Mux.scala 31:69:@8938.4]
  wire [5:0] _T_28347; // @[Mux.scala 31:69:@8939.4]
  wire [5:0] _T_28348; // @[Mux.scala 31:69:@8940.4]
  wire [5:0] _T_28349; // @[Mux.scala 31:69:@8941.4]
  wire [5:0] _T_28350; // @[Mux.scala 31:69:@8942.4]
  wire [5:0] _T_28351; // @[Mux.scala 31:69:@8943.4]
  wire [5:0] _T_28352; // @[Mux.scala 31:69:@8944.4]
  wire [5:0] _T_28353; // @[Mux.scala 31:69:@8945.4]
  wire [5:0] _T_28354; // @[Mux.scala 31:69:@8946.4]
  wire [5:0] _T_28355; // @[Mux.scala 31:69:@8947.4]
  wire [5:0] _T_28356; // @[Mux.scala 31:69:@8948.4]
  wire [5:0] _T_28357; // @[Mux.scala 31:69:@8949.4]
  wire [5:0] _T_28358; // @[Mux.scala 31:69:@8950.4]
  wire [5:0] _T_28359; // @[Mux.scala 31:69:@8951.4]
  wire [5:0] _T_28360; // @[Mux.scala 31:69:@8952.4]
  wire [5:0] _T_28361; // @[Mux.scala 31:69:@8953.4]
  wire [5:0] _T_28362; // @[Mux.scala 31:69:@8954.4]
  wire [5:0] _T_28363; // @[Mux.scala 31:69:@8955.4]
  wire [5:0] _T_28364; // @[Mux.scala 31:69:@8956.4]
  wire [5:0] _T_28365; // @[Mux.scala 31:69:@8957.4]
  wire [5:0] select_27; // @[Mux.scala 31:69:@8958.4]
  wire [47:0] _GEN_1729; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1730; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1731; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1732; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1733; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1734; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1735; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1736; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1737; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1738; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1739; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1740; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1741; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1742; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1743; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1744; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1745; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1746; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1747; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1748; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1749; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1750; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1751; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1752; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1753; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1754; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1755; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1756; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1757; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1758; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1759; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1760; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1761; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1762; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1763; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1764; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1765; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1766; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1767; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1768; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1769; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1770; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1771; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1772; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1773; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1774; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1775; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1776; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1777; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1778; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1779; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1780; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1781; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1782; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1783; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1784; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1785; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1786; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1787; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1788; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1789; // @[Switch.scala 33:19:@8960.4]
  wire [47:0] _GEN_1790; // @[Switch.scala 33:19:@8960.4]
  wire [7:0] _T_28374; // @[Switch.scala 34:32:@8967.4]
  wire [15:0] _T_28382; // @[Switch.scala 34:32:@8975.4]
  wire [7:0] _T_28389; // @[Switch.scala 34:32:@8982.4]
  wire [31:0] _T_28398; // @[Switch.scala 34:32:@8991.4]
  wire [7:0] _T_28405; // @[Switch.scala 34:32:@8998.4]
  wire [15:0] _T_28413; // @[Switch.scala 34:32:@9006.4]
  wire [7:0] _T_28420; // @[Switch.scala 34:32:@9013.4]
  wire [31:0] _T_28429; // @[Switch.scala 34:32:@9022.4]
  wire [63:0] _T_28430; // @[Switch.scala 34:32:@9023.4]
  wire  _T_28434; // @[Switch.scala 30:53:@9026.4]
  wire  valid_28_0; // @[Switch.scala 30:36:@9027.4]
  wire  _T_28437; // @[Switch.scala 30:53:@9029.4]
  wire  valid_28_1; // @[Switch.scala 30:36:@9030.4]
  wire  _T_28440; // @[Switch.scala 30:53:@9032.4]
  wire  valid_28_2; // @[Switch.scala 30:36:@9033.4]
  wire  _T_28443; // @[Switch.scala 30:53:@9035.4]
  wire  valid_28_3; // @[Switch.scala 30:36:@9036.4]
  wire  _T_28446; // @[Switch.scala 30:53:@9038.4]
  wire  valid_28_4; // @[Switch.scala 30:36:@9039.4]
  wire  _T_28449; // @[Switch.scala 30:53:@9041.4]
  wire  valid_28_5; // @[Switch.scala 30:36:@9042.4]
  wire  _T_28452; // @[Switch.scala 30:53:@9044.4]
  wire  valid_28_6; // @[Switch.scala 30:36:@9045.4]
  wire  _T_28455; // @[Switch.scala 30:53:@9047.4]
  wire  valid_28_7; // @[Switch.scala 30:36:@9048.4]
  wire  _T_28458; // @[Switch.scala 30:53:@9050.4]
  wire  valid_28_8; // @[Switch.scala 30:36:@9051.4]
  wire  _T_28461; // @[Switch.scala 30:53:@9053.4]
  wire  valid_28_9; // @[Switch.scala 30:36:@9054.4]
  wire  _T_28464; // @[Switch.scala 30:53:@9056.4]
  wire  valid_28_10; // @[Switch.scala 30:36:@9057.4]
  wire  _T_28467; // @[Switch.scala 30:53:@9059.4]
  wire  valid_28_11; // @[Switch.scala 30:36:@9060.4]
  wire  _T_28470; // @[Switch.scala 30:53:@9062.4]
  wire  valid_28_12; // @[Switch.scala 30:36:@9063.4]
  wire  _T_28473; // @[Switch.scala 30:53:@9065.4]
  wire  valid_28_13; // @[Switch.scala 30:36:@9066.4]
  wire  _T_28476; // @[Switch.scala 30:53:@9068.4]
  wire  valid_28_14; // @[Switch.scala 30:36:@9069.4]
  wire  _T_28479; // @[Switch.scala 30:53:@9071.4]
  wire  valid_28_15; // @[Switch.scala 30:36:@9072.4]
  wire  _T_28482; // @[Switch.scala 30:53:@9074.4]
  wire  valid_28_16; // @[Switch.scala 30:36:@9075.4]
  wire  _T_28485; // @[Switch.scala 30:53:@9077.4]
  wire  valid_28_17; // @[Switch.scala 30:36:@9078.4]
  wire  _T_28488; // @[Switch.scala 30:53:@9080.4]
  wire  valid_28_18; // @[Switch.scala 30:36:@9081.4]
  wire  _T_28491; // @[Switch.scala 30:53:@9083.4]
  wire  valid_28_19; // @[Switch.scala 30:36:@9084.4]
  wire  _T_28494; // @[Switch.scala 30:53:@9086.4]
  wire  valid_28_20; // @[Switch.scala 30:36:@9087.4]
  wire  _T_28497; // @[Switch.scala 30:53:@9089.4]
  wire  valid_28_21; // @[Switch.scala 30:36:@9090.4]
  wire  _T_28500; // @[Switch.scala 30:53:@9092.4]
  wire  valid_28_22; // @[Switch.scala 30:36:@9093.4]
  wire  _T_28503; // @[Switch.scala 30:53:@9095.4]
  wire  valid_28_23; // @[Switch.scala 30:36:@9096.4]
  wire  _T_28506; // @[Switch.scala 30:53:@9098.4]
  wire  valid_28_24; // @[Switch.scala 30:36:@9099.4]
  wire  _T_28509; // @[Switch.scala 30:53:@9101.4]
  wire  valid_28_25; // @[Switch.scala 30:36:@9102.4]
  wire  _T_28512; // @[Switch.scala 30:53:@9104.4]
  wire  valid_28_26; // @[Switch.scala 30:36:@9105.4]
  wire  _T_28515; // @[Switch.scala 30:53:@9107.4]
  wire  valid_28_27; // @[Switch.scala 30:36:@9108.4]
  wire  _T_28518; // @[Switch.scala 30:53:@9110.4]
  wire  valid_28_28; // @[Switch.scala 30:36:@9111.4]
  wire  _T_28521; // @[Switch.scala 30:53:@9113.4]
  wire  valid_28_29; // @[Switch.scala 30:36:@9114.4]
  wire  _T_28524; // @[Switch.scala 30:53:@9116.4]
  wire  valid_28_30; // @[Switch.scala 30:36:@9117.4]
  wire  _T_28527; // @[Switch.scala 30:53:@9119.4]
  wire  valid_28_31; // @[Switch.scala 30:36:@9120.4]
  wire  _T_28530; // @[Switch.scala 30:53:@9122.4]
  wire  valid_28_32; // @[Switch.scala 30:36:@9123.4]
  wire  _T_28533; // @[Switch.scala 30:53:@9125.4]
  wire  valid_28_33; // @[Switch.scala 30:36:@9126.4]
  wire  _T_28536; // @[Switch.scala 30:53:@9128.4]
  wire  valid_28_34; // @[Switch.scala 30:36:@9129.4]
  wire  _T_28539; // @[Switch.scala 30:53:@9131.4]
  wire  valid_28_35; // @[Switch.scala 30:36:@9132.4]
  wire  _T_28542; // @[Switch.scala 30:53:@9134.4]
  wire  valid_28_36; // @[Switch.scala 30:36:@9135.4]
  wire  _T_28545; // @[Switch.scala 30:53:@9137.4]
  wire  valid_28_37; // @[Switch.scala 30:36:@9138.4]
  wire  _T_28548; // @[Switch.scala 30:53:@9140.4]
  wire  valid_28_38; // @[Switch.scala 30:36:@9141.4]
  wire  _T_28551; // @[Switch.scala 30:53:@9143.4]
  wire  valid_28_39; // @[Switch.scala 30:36:@9144.4]
  wire  _T_28554; // @[Switch.scala 30:53:@9146.4]
  wire  valid_28_40; // @[Switch.scala 30:36:@9147.4]
  wire  _T_28557; // @[Switch.scala 30:53:@9149.4]
  wire  valid_28_41; // @[Switch.scala 30:36:@9150.4]
  wire  _T_28560; // @[Switch.scala 30:53:@9152.4]
  wire  valid_28_42; // @[Switch.scala 30:36:@9153.4]
  wire  _T_28563; // @[Switch.scala 30:53:@9155.4]
  wire  valid_28_43; // @[Switch.scala 30:36:@9156.4]
  wire  _T_28566; // @[Switch.scala 30:53:@9158.4]
  wire  valid_28_44; // @[Switch.scala 30:36:@9159.4]
  wire  _T_28569; // @[Switch.scala 30:53:@9161.4]
  wire  valid_28_45; // @[Switch.scala 30:36:@9162.4]
  wire  _T_28572; // @[Switch.scala 30:53:@9164.4]
  wire  valid_28_46; // @[Switch.scala 30:36:@9165.4]
  wire  _T_28575; // @[Switch.scala 30:53:@9167.4]
  wire  valid_28_47; // @[Switch.scala 30:36:@9168.4]
  wire  _T_28578; // @[Switch.scala 30:53:@9170.4]
  wire  valid_28_48; // @[Switch.scala 30:36:@9171.4]
  wire  _T_28581; // @[Switch.scala 30:53:@9173.4]
  wire  valid_28_49; // @[Switch.scala 30:36:@9174.4]
  wire  _T_28584; // @[Switch.scala 30:53:@9176.4]
  wire  valid_28_50; // @[Switch.scala 30:36:@9177.4]
  wire  _T_28587; // @[Switch.scala 30:53:@9179.4]
  wire  valid_28_51; // @[Switch.scala 30:36:@9180.4]
  wire  _T_28590; // @[Switch.scala 30:53:@9182.4]
  wire  valid_28_52; // @[Switch.scala 30:36:@9183.4]
  wire  _T_28593; // @[Switch.scala 30:53:@9185.4]
  wire  valid_28_53; // @[Switch.scala 30:36:@9186.4]
  wire  _T_28596; // @[Switch.scala 30:53:@9188.4]
  wire  valid_28_54; // @[Switch.scala 30:36:@9189.4]
  wire  _T_28599; // @[Switch.scala 30:53:@9191.4]
  wire  valid_28_55; // @[Switch.scala 30:36:@9192.4]
  wire  _T_28602; // @[Switch.scala 30:53:@9194.4]
  wire  valid_28_56; // @[Switch.scala 30:36:@9195.4]
  wire  _T_28605; // @[Switch.scala 30:53:@9197.4]
  wire  valid_28_57; // @[Switch.scala 30:36:@9198.4]
  wire  _T_28608; // @[Switch.scala 30:53:@9200.4]
  wire  valid_28_58; // @[Switch.scala 30:36:@9201.4]
  wire  _T_28611; // @[Switch.scala 30:53:@9203.4]
  wire  valid_28_59; // @[Switch.scala 30:36:@9204.4]
  wire  _T_28614; // @[Switch.scala 30:53:@9206.4]
  wire  valid_28_60; // @[Switch.scala 30:36:@9207.4]
  wire  _T_28617; // @[Switch.scala 30:53:@9209.4]
  wire  valid_28_61; // @[Switch.scala 30:36:@9210.4]
  wire  _T_28620; // @[Switch.scala 30:53:@9212.4]
  wire  valid_28_62; // @[Switch.scala 30:36:@9213.4]
  wire  _T_28623; // @[Switch.scala 30:53:@9215.4]
  wire  valid_28_63; // @[Switch.scala 30:36:@9216.4]
  wire [5:0] _T_28689; // @[Mux.scala 31:69:@9218.4]
  wire [5:0] _T_28690; // @[Mux.scala 31:69:@9219.4]
  wire [5:0] _T_28691; // @[Mux.scala 31:69:@9220.4]
  wire [5:0] _T_28692; // @[Mux.scala 31:69:@9221.4]
  wire [5:0] _T_28693; // @[Mux.scala 31:69:@9222.4]
  wire [5:0] _T_28694; // @[Mux.scala 31:69:@9223.4]
  wire [5:0] _T_28695; // @[Mux.scala 31:69:@9224.4]
  wire [5:0] _T_28696; // @[Mux.scala 31:69:@9225.4]
  wire [5:0] _T_28697; // @[Mux.scala 31:69:@9226.4]
  wire [5:0] _T_28698; // @[Mux.scala 31:69:@9227.4]
  wire [5:0] _T_28699; // @[Mux.scala 31:69:@9228.4]
  wire [5:0] _T_28700; // @[Mux.scala 31:69:@9229.4]
  wire [5:0] _T_28701; // @[Mux.scala 31:69:@9230.4]
  wire [5:0] _T_28702; // @[Mux.scala 31:69:@9231.4]
  wire [5:0] _T_28703; // @[Mux.scala 31:69:@9232.4]
  wire [5:0] _T_28704; // @[Mux.scala 31:69:@9233.4]
  wire [5:0] _T_28705; // @[Mux.scala 31:69:@9234.4]
  wire [5:0] _T_28706; // @[Mux.scala 31:69:@9235.4]
  wire [5:0] _T_28707; // @[Mux.scala 31:69:@9236.4]
  wire [5:0] _T_28708; // @[Mux.scala 31:69:@9237.4]
  wire [5:0] _T_28709; // @[Mux.scala 31:69:@9238.4]
  wire [5:0] _T_28710; // @[Mux.scala 31:69:@9239.4]
  wire [5:0] _T_28711; // @[Mux.scala 31:69:@9240.4]
  wire [5:0] _T_28712; // @[Mux.scala 31:69:@9241.4]
  wire [5:0] _T_28713; // @[Mux.scala 31:69:@9242.4]
  wire [5:0] _T_28714; // @[Mux.scala 31:69:@9243.4]
  wire [5:0] _T_28715; // @[Mux.scala 31:69:@9244.4]
  wire [5:0] _T_28716; // @[Mux.scala 31:69:@9245.4]
  wire [5:0] _T_28717; // @[Mux.scala 31:69:@9246.4]
  wire [5:0] _T_28718; // @[Mux.scala 31:69:@9247.4]
  wire [5:0] _T_28719; // @[Mux.scala 31:69:@9248.4]
  wire [5:0] _T_28720; // @[Mux.scala 31:69:@9249.4]
  wire [5:0] _T_28721; // @[Mux.scala 31:69:@9250.4]
  wire [5:0] _T_28722; // @[Mux.scala 31:69:@9251.4]
  wire [5:0] _T_28723; // @[Mux.scala 31:69:@9252.4]
  wire [5:0] _T_28724; // @[Mux.scala 31:69:@9253.4]
  wire [5:0] _T_28725; // @[Mux.scala 31:69:@9254.4]
  wire [5:0] _T_28726; // @[Mux.scala 31:69:@9255.4]
  wire [5:0] _T_28727; // @[Mux.scala 31:69:@9256.4]
  wire [5:0] _T_28728; // @[Mux.scala 31:69:@9257.4]
  wire [5:0] _T_28729; // @[Mux.scala 31:69:@9258.4]
  wire [5:0] _T_28730; // @[Mux.scala 31:69:@9259.4]
  wire [5:0] _T_28731; // @[Mux.scala 31:69:@9260.4]
  wire [5:0] _T_28732; // @[Mux.scala 31:69:@9261.4]
  wire [5:0] _T_28733; // @[Mux.scala 31:69:@9262.4]
  wire [5:0] _T_28734; // @[Mux.scala 31:69:@9263.4]
  wire [5:0] _T_28735; // @[Mux.scala 31:69:@9264.4]
  wire [5:0] _T_28736; // @[Mux.scala 31:69:@9265.4]
  wire [5:0] _T_28737; // @[Mux.scala 31:69:@9266.4]
  wire [5:0] _T_28738; // @[Mux.scala 31:69:@9267.4]
  wire [5:0] _T_28739; // @[Mux.scala 31:69:@9268.4]
  wire [5:0] _T_28740; // @[Mux.scala 31:69:@9269.4]
  wire [5:0] _T_28741; // @[Mux.scala 31:69:@9270.4]
  wire [5:0] _T_28742; // @[Mux.scala 31:69:@9271.4]
  wire [5:0] _T_28743; // @[Mux.scala 31:69:@9272.4]
  wire [5:0] _T_28744; // @[Mux.scala 31:69:@9273.4]
  wire [5:0] _T_28745; // @[Mux.scala 31:69:@9274.4]
  wire [5:0] _T_28746; // @[Mux.scala 31:69:@9275.4]
  wire [5:0] _T_28747; // @[Mux.scala 31:69:@9276.4]
  wire [5:0] _T_28748; // @[Mux.scala 31:69:@9277.4]
  wire [5:0] _T_28749; // @[Mux.scala 31:69:@9278.4]
  wire [5:0] _T_28750; // @[Mux.scala 31:69:@9279.4]
  wire [5:0] select_28; // @[Mux.scala 31:69:@9280.4]
  wire [47:0] _GEN_1793; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1794; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1795; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1796; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1797; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1798; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1799; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1800; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1801; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1802; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1803; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1804; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1805; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1806; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1807; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1808; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1809; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1810; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1811; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1812; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1813; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1814; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1815; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1816; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1817; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1818; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1819; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1820; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1821; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1822; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1823; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1824; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1825; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1826; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1827; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1828; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1829; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1830; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1831; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1832; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1833; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1834; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1835; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1836; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1837; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1838; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1839; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1840; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1841; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1842; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1843; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1844; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1845; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1846; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1847; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1848; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1849; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1850; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1851; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1852; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1853; // @[Switch.scala 33:19:@9282.4]
  wire [47:0] _GEN_1854; // @[Switch.scala 33:19:@9282.4]
  wire [7:0] _T_28759; // @[Switch.scala 34:32:@9289.4]
  wire [15:0] _T_28767; // @[Switch.scala 34:32:@9297.4]
  wire [7:0] _T_28774; // @[Switch.scala 34:32:@9304.4]
  wire [31:0] _T_28783; // @[Switch.scala 34:32:@9313.4]
  wire [7:0] _T_28790; // @[Switch.scala 34:32:@9320.4]
  wire [15:0] _T_28798; // @[Switch.scala 34:32:@9328.4]
  wire [7:0] _T_28805; // @[Switch.scala 34:32:@9335.4]
  wire [31:0] _T_28814; // @[Switch.scala 34:32:@9344.4]
  wire [63:0] _T_28815; // @[Switch.scala 34:32:@9345.4]
  wire  _T_28819; // @[Switch.scala 30:53:@9348.4]
  wire  valid_29_0; // @[Switch.scala 30:36:@9349.4]
  wire  _T_28822; // @[Switch.scala 30:53:@9351.4]
  wire  valid_29_1; // @[Switch.scala 30:36:@9352.4]
  wire  _T_28825; // @[Switch.scala 30:53:@9354.4]
  wire  valid_29_2; // @[Switch.scala 30:36:@9355.4]
  wire  _T_28828; // @[Switch.scala 30:53:@9357.4]
  wire  valid_29_3; // @[Switch.scala 30:36:@9358.4]
  wire  _T_28831; // @[Switch.scala 30:53:@9360.4]
  wire  valid_29_4; // @[Switch.scala 30:36:@9361.4]
  wire  _T_28834; // @[Switch.scala 30:53:@9363.4]
  wire  valid_29_5; // @[Switch.scala 30:36:@9364.4]
  wire  _T_28837; // @[Switch.scala 30:53:@9366.4]
  wire  valid_29_6; // @[Switch.scala 30:36:@9367.4]
  wire  _T_28840; // @[Switch.scala 30:53:@9369.4]
  wire  valid_29_7; // @[Switch.scala 30:36:@9370.4]
  wire  _T_28843; // @[Switch.scala 30:53:@9372.4]
  wire  valid_29_8; // @[Switch.scala 30:36:@9373.4]
  wire  _T_28846; // @[Switch.scala 30:53:@9375.4]
  wire  valid_29_9; // @[Switch.scala 30:36:@9376.4]
  wire  _T_28849; // @[Switch.scala 30:53:@9378.4]
  wire  valid_29_10; // @[Switch.scala 30:36:@9379.4]
  wire  _T_28852; // @[Switch.scala 30:53:@9381.4]
  wire  valid_29_11; // @[Switch.scala 30:36:@9382.4]
  wire  _T_28855; // @[Switch.scala 30:53:@9384.4]
  wire  valid_29_12; // @[Switch.scala 30:36:@9385.4]
  wire  _T_28858; // @[Switch.scala 30:53:@9387.4]
  wire  valid_29_13; // @[Switch.scala 30:36:@9388.4]
  wire  _T_28861; // @[Switch.scala 30:53:@9390.4]
  wire  valid_29_14; // @[Switch.scala 30:36:@9391.4]
  wire  _T_28864; // @[Switch.scala 30:53:@9393.4]
  wire  valid_29_15; // @[Switch.scala 30:36:@9394.4]
  wire  _T_28867; // @[Switch.scala 30:53:@9396.4]
  wire  valid_29_16; // @[Switch.scala 30:36:@9397.4]
  wire  _T_28870; // @[Switch.scala 30:53:@9399.4]
  wire  valid_29_17; // @[Switch.scala 30:36:@9400.4]
  wire  _T_28873; // @[Switch.scala 30:53:@9402.4]
  wire  valid_29_18; // @[Switch.scala 30:36:@9403.4]
  wire  _T_28876; // @[Switch.scala 30:53:@9405.4]
  wire  valid_29_19; // @[Switch.scala 30:36:@9406.4]
  wire  _T_28879; // @[Switch.scala 30:53:@9408.4]
  wire  valid_29_20; // @[Switch.scala 30:36:@9409.4]
  wire  _T_28882; // @[Switch.scala 30:53:@9411.4]
  wire  valid_29_21; // @[Switch.scala 30:36:@9412.4]
  wire  _T_28885; // @[Switch.scala 30:53:@9414.4]
  wire  valid_29_22; // @[Switch.scala 30:36:@9415.4]
  wire  _T_28888; // @[Switch.scala 30:53:@9417.4]
  wire  valid_29_23; // @[Switch.scala 30:36:@9418.4]
  wire  _T_28891; // @[Switch.scala 30:53:@9420.4]
  wire  valid_29_24; // @[Switch.scala 30:36:@9421.4]
  wire  _T_28894; // @[Switch.scala 30:53:@9423.4]
  wire  valid_29_25; // @[Switch.scala 30:36:@9424.4]
  wire  _T_28897; // @[Switch.scala 30:53:@9426.4]
  wire  valid_29_26; // @[Switch.scala 30:36:@9427.4]
  wire  _T_28900; // @[Switch.scala 30:53:@9429.4]
  wire  valid_29_27; // @[Switch.scala 30:36:@9430.4]
  wire  _T_28903; // @[Switch.scala 30:53:@9432.4]
  wire  valid_29_28; // @[Switch.scala 30:36:@9433.4]
  wire  _T_28906; // @[Switch.scala 30:53:@9435.4]
  wire  valid_29_29; // @[Switch.scala 30:36:@9436.4]
  wire  _T_28909; // @[Switch.scala 30:53:@9438.4]
  wire  valid_29_30; // @[Switch.scala 30:36:@9439.4]
  wire  _T_28912; // @[Switch.scala 30:53:@9441.4]
  wire  valid_29_31; // @[Switch.scala 30:36:@9442.4]
  wire  _T_28915; // @[Switch.scala 30:53:@9444.4]
  wire  valid_29_32; // @[Switch.scala 30:36:@9445.4]
  wire  _T_28918; // @[Switch.scala 30:53:@9447.4]
  wire  valid_29_33; // @[Switch.scala 30:36:@9448.4]
  wire  _T_28921; // @[Switch.scala 30:53:@9450.4]
  wire  valid_29_34; // @[Switch.scala 30:36:@9451.4]
  wire  _T_28924; // @[Switch.scala 30:53:@9453.4]
  wire  valid_29_35; // @[Switch.scala 30:36:@9454.4]
  wire  _T_28927; // @[Switch.scala 30:53:@9456.4]
  wire  valid_29_36; // @[Switch.scala 30:36:@9457.4]
  wire  _T_28930; // @[Switch.scala 30:53:@9459.4]
  wire  valid_29_37; // @[Switch.scala 30:36:@9460.4]
  wire  _T_28933; // @[Switch.scala 30:53:@9462.4]
  wire  valid_29_38; // @[Switch.scala 30:36:@9463.4]
  wire  _T_28936; // @[Switch.scala 30:53:@9465.4]
  wire  valid_29_39; // @[Switch.scala 30:36:@9466.4]
  wire  _T_28939; // @[Switch.scala 30:53:@9468.4]
  wire  valid_29_40; // @[Switch.scala 30:36:@9469.4]
  wire  _T_28942; // @[Switch.scala 30:53:@9471.4]
  wire  valid_29_41; // @[Switch.scala 30:36:@9472.4]
  wire  _T_28945; // @[Switch.scala 30:53:@9474.4]
  wire  valid_29_42; // @[Switch.scala 30:36:@9475.4]
  wire  _T_28948; // @[Switch.scala 30:53:@9477.4]
  wire  valid_29_43; // @[Switch.scala 30:36:@9478.4]
  wire  _T_28951; // @[Switch.scala 30:53:@9480.4]
  wire  valid_29_44; // @[Switch.scala 30:36:@9481.4]
  wire  _T_28954; // @[Switch.scala 30:53:@9483.4]
  wire  valid_29_45; // @[Switch.scala 30:36:@9484.4]
  wire  _T_28957; // @[Switch.scala 30:53:@9486.4]
  wire  valid_29_46; // @[Switch.scala 30:36:@9487.4]
  wire  _T_28960; // @[Switch.scala 30:53:@9489.4]
  wire  valid_29_47; // @[Switch.scala 30:36:@9490.4]
  wire  _T_28963; // @[Switch.scala 30:53:@9492.4]
  wire  valid_29_48; // @[Switch.scala 30:36:@9493.4]
  wire  _T_28966; // @[Switch.scala 30:53:@9495.4]
  wire  valid_29_49; // @[Switch.scala 30:36:@9496.4]
  wire  _T_28969; // @[Switch.scala 30:53:@9498.4]
  wire  valid_29_50; // @[Switch.scala 30:36:@9499.4]
  wire  _T_28972; // @[Switch.scala 30:53:@9501.4]
  wire  valid_29_51; // @[Switch.scala 30:36:@9502.4]
  wire  _T_28975; // @[Switch.scala 30:53:@9504.4]
  wire  valid_29_52; // @[Switch.scala 30:36:@9505.4]
  wire  _T_28978; // @[Switch.scala 30:53:@9507.4]
  wire  valid_29_53; // @[Switch.scala 30:36:@9508.4]
  wire  _T_28981; // @[Switch.scala 30:53:@9510.4]
  wire  valid_29_54; // @[Switch.scala 30:36:@9511.4]
  wire  _T_28984; // @[Switch.scala 30:53:@9513.4]
  wire  valid_29_55; // @[Switch.scala 30:36:@9514.4]
  wire  _T_28987; // @[Switch.scala 30:53:@9516.4]
  wire  valid_29_56; // @[Switch.scala 30:36:@9517.4]
  wire  _T_28990; // @[Switch.scala 30:53:@9519.4]
  wire  valid_29_57; // @[Switch.scala 30:36:@9520.4]
  wire  _T_28993; // @[Switch.scala 30:53:@9522.4]
  wire  valid_29_58; // @[Switch.scala 30:36:@9523.4]
  wire  _T_28996; // @[Switch.scala 30:53:@9525.4]
  wire  valid_29_59; // @[Switch.scala 30:36:@9526.4]
  wire  _T_28999; // @[Switch.scala 30:53:@9528.4]
  wire  valid_29_60; // @[Switch.scala 30:36:@9529.4]
  wire  _T_29002; // @[Switch.scala 30:53:@9531.4]
  wire  valid_29_61; // @[Switch.scala 30:36:@9532.4]
  wire  _T_29005; // @[Switch.scala 30:53:@9534.4]
  wire  valid_29_62; // @[Switch.scala 30:36:@9535.4]
  wire  _T_29008; // @[Switch.scala 30:53:@9537.4]
  wire  valid_29_63; // @[Switch.scala 30:36:@9538.4]
  wire [5:0] _T_29074; // @[Mux.scala 31:69:@9540.4]
  wire [5:0] _T_29075; // @[Mux.scala 31:69:@9541.4]
  wire [5:0] _T_29076; // @[Mux.scala 31:69:@9542.4]
  wire [5:0] _T_29077; // @[Mux.scala 31:69:@9543.4]
  wire [5:0] _T_29078; // @[Mux.scala 31:69:@9544.4]
  wire [5:0] _T_29079; // @[Mux.scala 31:69:@9545.4]
  wire [5:0] _T_29080; // @[Mux.scala 31:69:@9546.4]
  wire [5:0] _T_29081; // @[Mux.scala 31:69:@9547.4]
  wire [5:0] _T_29082; // @[Mux.scala 31:69:@9548.4]
  wire [5:0] _T_29083; // @[Mux.scala 31:69:@9549.4]
  wire [5:0] _T_29084; // @[Mux.scala 31:69:@9550.4]
  wire [5:0] _T_29085; // @[Mux.scala 31:69:@9551.4]
  wire [5:0] _T_29086; // @[Mux.scala 31:69:@9552.4]
  wire [5:0] _T_29087; // @[Mux.scala 31:69:@9553.4]
  wire [5:0] _T_29088; // @[Mux.scala 31:69:@9554.4]
  wire [5:0] _T_29089; // @[Mux.scala 31:69:@9555.4]
  wire [5:0] _T_29090; // @[Mux.scala 31:69:@9556.4]
  wire [5:0] _T_29091; // @[Mux.scala 31:69:@9557.4]
  wire [5:0] _T_29092; // @[Mux.scala 31:69:@9558.4]
  wire [5:0] _T_29093; // @[Mux.scala 31:69:@9559.4]
  wire [5:0] _T_29094; // @[Mux.scala 31:69:@9560.4]
  wire [5:0] _T_29095; // @[Mux.scala 31:69:@9561.4]
  wire [5:0] _T_29096; // @[Mux.scala 31:69:@9562.4]
  wire [5:0] _T_29097; // @[Mux.scala 31:69:@9563.4]
  wire [5:0] _T_29098; // @[Mux.scala 31:69:@9564.4]
  wire [5:0] _T_29099; // @[Mux.scala 31:69:@9565.4]
  wire [5:0] _T_29100; // @[Mux.scala 31:69:@9566.4]
  wire [5:0] _T_29101; // @[Mux.scala 31:69:@9567.4]
  wire [5:0] _T_29102; // @[Mux.scala 31:69:@9568.4]
  wire [5:0] _T_29103; // @[Mux.scala 31:69:@9569.4]
  wire [5:0] _T_29104; // @[Mux.scala 31:69:@9570.4]
  wire [5:0] _T_29105; // @[Mux.scala 31:69:@9571.4]
  wire [5:0] _T_29106; // @[Mux.scala 31:69:@9572.4]
  wire [5:0] _T_29107; // @[Mux.scala 31:69:@9573.4]
  wire [5:0] _T_29108; // @[Mux.scala 31:69:@9574.4]
  wire [5:0] _T_29109; // @[Mux.scala 31:69:@9575.4]
  wire [5:0] _T_29110; // @[Mux.scala 31:69:@9576.4]
  wire [5:0] _T_29111; // @[Mux.scala 31:69:@9577.4]
  wire [5:0] _T_29112; // @[Mux.scala 31:69:@9578.4]
  wire [5:0] _T_29113; // @[Mux.scala 31:69:@9579.4]
  wire [5:0] _T_29114; // @[Mux.scala 31:69:@9580.4]
  wire [5:0] _T_29115; // @[Mux.scala 31:69:@9581.4]
  wire [5:0] _T_29116; // @[Mux.scala 31:69:@9582.4]
  wire [5:0] _T_29117; // @[Mux.scala 31:69:@9583.4]
  wire [5:0] _T_29118; // @[Mux.scala 31:69:@9584.4]
  wire [5:0] _T_29119; // @[Mux.scala 31:69:@9585.4]
  wire [5:0] _T_29120; // @[Mux.scala 31:69:@9586.4]
  wire [5:0] _T_29121; // @[Mux.scala 31:69:@9587.4]
  wire [5:0] _T_29122; // @[Mux.scala 31:69:@9588.4]
  wire [5:0] _T_29123; // @[Mux.scala 31:69:@9589.4]
  wire [5:0] _T_29124; // @[Mux.scala 31:69:@9590.4]
  wire [5:0] _T_29125; // @[Mux.scala 31:69:@9591.4]
  wire [5:0] _T_29126; // @[Mux.scala 31:69:@9592.4]
  wire [5:0] _T_29127; // @[Mux.scala 31:69:@9593.4]
  wire [5:0] _T_29128; // @[Mux.scala 31:69:@9594.4]
  wire [5:0] _T_29129; // @[Mux.scala 31:69:@9595.4]
  wire [5:0] _T_29130; // @[Mux.scala 31:69:@9596.4]
  wire [5:0] _T_29131; // @[Mux.scala 31:69:@9597.4]
  wire [5:0] _T_29132; // @[Mux.scala 31:69:@9598.4]
  wire [5:0] _T_29133; // @[Mux.scala 31:69:@9599.4]
  wire [5:0] _T_29134; // @[Mux.scala 31:69:@9600.4]
  wire [5:0] _T_29135; // @[Mux.scala 31:69:@9601.4]
  wire [5:0] select_29; // @[Mux.scala 31:69:@9602.4]
  wire [47:0] _GEN_1857; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1858; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1859; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1860; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1861; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1862; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1863; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1864; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1865; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1866; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1867; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1868; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1869; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1870; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1871; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1872; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1873; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1874; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1875; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1876; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1877; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1878; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1879; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1880; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1881; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1882; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1883; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1884; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1885; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1886; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1887; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1888; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1889; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1890; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1891; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1892; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1893; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1894; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1895; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1896; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1897; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1898; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1899; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1900; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1901; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1902; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1903; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1904; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1905; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1906; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1907; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1908; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1909; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1910; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1911; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1912; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1913; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1914; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1915; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1916; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1917; // @[Switch.scala 33:19:@9604.4]
  wire [47:0] _GEN_1918; // @[Switch.scala 33:19:@9604.4]
  wire [7:0] _T_29144; // @[Switch.scala 34:32:@9611.4]
  wire [15:0] _T_29152; // @[Switch.scala 34:32:@9619.4]
  wire [7:0] _T_29159; // @[Switch.scala 34:32:@9626.4]
  wire [31:0] _T_29168; // @[Switch.scala 34:32:@9635.4]
  wire [7:0] _T_29175; // @[Switch.scala 34:32:@9642.4]
  wire [15:0] _T_29183; // @[Switch.scala 34:32:@9650.4]
  wire [7:0] _T_29190; // @[Switch.scala 34:32:@9657.4]
  wire [31:0] _T_29199; // @[Switch.scala 34:32:@9666.4]
  wire [63:0] _T_29200; // @[Switch.scala 34:32:@9667.4]
  wire  _T_29204; // @[Switch.scala 30:53:@9670.4]
  wire  valid_30_0; // @[Switch.scala 30:36:@9671.4]
  wire  _T_29207; // @[Switch.scala 30:53:@9673.4]
  wire  valid_30_1; // @[Switch.scala 30:36:@9674.4]
  wire  _T_29210; // @[Switch.scala 30:53:@9676.4]
  wire  valid_30_2; // @[Switch.scala 30:36:@9677.4]
  wire  _T_29213; // @[Switch.scala 30:53:@9679.4]
  wire  valid_30_3; // @[Switch.scala 30:36:@9680.4]
  wire  _T_29216; // @[Switch.scala 30:53:@9682.4]
  wire  valid_30_4; // @[Switch.scala 30:36:@9683.4]
  wire  _T_29219; // @[Switch.scala 30:53:@9685.4]
  wire  valid_30_5; // @[Switch.scala 30:36:@9686.4]
  wire  _T_29222; // @[Switch.scala 30:53:@9688.4]
  wire  valid_30_6; // @[Switch.scala 30:36:@9689.4]
  wire  _T_29225; // @[Switch.scala 30:53:@9691.4]
  wire  valid_30_7; // @[Switch.scala 30:36:@9692.4]
  wire  _T_29228; // @[Switch.scala 30:53:@9694.4]
  wire  valid_30_8; // @[Switch.scala 30:36:@9695.4]
  wire  _T_29231; // @[Switch.scala 30:53:@9697.4]
  wire  valid_30_9; // @[Switch.scala 30:36:@9698.4]
  wire  _T_29234; // @[Switch.scala 30:53:@9700.4]
  wire  valid_30_10; // @[Switch.scala 30:36:@9701.4]
  wire  _T_29237; // @[Switch.scala 30:53:@9703.4]
  wire  valid_30_11; // @[Switch.scala 30:36:@9704.4]
  wire  _T_29240; // @[Switch.scala 30:53:@9706.4]
  wire  valid_30_12; // @[Switch.scala 30:36:@9707.4]
  wire  _T_29243; // @[Switch.scala 30:53:@9709.4]
  wire  valid_30_13; // @[Switch.scala 30:36:@9710.4]
  wire  _T_29246; // @[Switch.scala 30:53:@9712.4]
  wire  valid_30_14; // @[Switch.scala 30:36:@9713.4]
  wire  _T_29249; // @[Switch.scala 30:53:@9715.4]
  wire  valid_30_15; // @[Switch.scala 30:36:@9716.4]
  wire  _T_29252; // @[Switch.scala 30:53:@9718.4]
  wire  valid_30_16; // @[Switch.scala 30:36:@9719.4]
  wire  _T_29255; // @[Switch.scala 30:53:@9721.4]
  wire  valid_30_17; // @[Switch.scala 30:36:@9722.4]
  wire  _T_29258; // @[Switch.scala 30:53:@9724.4]
  wire  valid_30_18; // @[Switch.scala 30:36:@9725.4]
  wire  _T_29261; // @[Switch.scala 30:53:@9727.4]
  wire  valid_30_19; // @[Switch.scala 30:36:@9728.4]
  wire  _T_29264; // @[Switch.scala 30:53:@9730.4]
  wire  valid_30_20; // @[Switch.scala 30:36:@9731.4]
  wire  _T_29267; // @[Switch.scala 30:53:@9733.4]
  wire  valid_30_21; // @[Switch.scala 30:36:@9734.4]
  wire  _T_29270; // @[Switch.scala 30:53:@9736.4]
  wire  valid_30_22; // @[Switch.scala 30:36:@9737.4]
  wire  _T_29273; // @[Switch.scala 30:53:@9739.4]
  wire  valid_30_23; // @[Switch.scala 30:36:@9740.4]
  wire  _T_29276; // @[Switch.scala 30:53:@9742.4]
  wire  valid_30_24; // @[Switch.scala 30:36:@9743.4]
  wire  _T_29279; // @[Switch.scala 30:53:@9745.4]
  wire  valid_30_25; // @[Switch.scala 30:36:@9746.4]
  wire  _T_29282; // @[Switch.scala 30:53:@9748.4]
  wire  valid_30_26; // @[Switch.scala 30:36:@9749.4]
  wire  _T_29285; // @[Switch.scala 30:53:@9751.4]
  wire  valid_30_27; // @[Switch.scala 30:36:@9752.4]
  wire  _T_29288; // @[Switch.scala 30:53:@9754.4]
  wire  valid_30_28; // @[Switch.scala 30:36:@9755.4]
  wire  _T_29291; // @[Switch.scala 30:53:@9757.4]
  wire  valid_30_29; // @[Switch.scala 30:36:@9758.4]
  wire  _T_29294; // @[Switch.scala 30:53:@9760.4]
  wire  valid_30_30; // @[Switch.scala 30:36:@9761.4]
  wire  _T_29297; // @[Switch.scala 30:53:@9763.4]
  wire  valid_30_31; // @[Switch.scala 30:36:@9764.4]
  wire  _T_29300; // @[Switch.scala 30:53:@9766.4]
  wire  valid_30_32; // @[Switch.scala 30:36:@9767.4]
  wire  _T_29303; // @[Switch.scala 30:53:@9769.4]
  wire  valid_30_33; // @[Switch.scala 30:36:@9770.4]
  wire  _T_29306; // @[Switch.scala 30:53:@9772.4]
  wire  valid_30_34; // @[Switch.scala 30:36:@9773.4]
  wire  _T_29309; // @[Switch.scala 30:53:@9775.4]
  wire  valid_30_35; // @[Switch.scala 30:36:@9776.4]
  wire  _T_29312; // @[Switch.scala 30:53:@9778.4]
  wire  valid_30_36; // @[Switch.scala 30:36:@9779.4]
  wire  _T_29315; // @[Switch.scala 30:53:@9781.4]
  wire  valid_30_37; // @[Switch.scala 30:36:@9782.4]
  wire  _T_29318; // @[Switch.scala 30:53:@9784.4]
  wire  valid_30_38; // @[Switch.scala 30:36:@9785.4]
  wire  _T_29321; // @[Switch.scala 30:53:@9787.4]
  wire  valid_30_39; // @[Switch.scala 30:36:@9788.4]
  wire  _T_29324; // @[Switch.scala 30:53:@9790.4]
  wire  valid_30_40; // @[Switch.scala 30:36:@9791.4]
  wire  _T_29327; // @[Switch.scala 30:53:@9793.4]
  wire  valid_30_41; // @[Switch.scala 30:36:@9794.4]
  wire  _T_29330; // @[Switch.scala 30:53:@9796.4]
  wire  valid_30_42; // @[Switch.scala 30:36:@9797.4]
  wire  _T_29333; // @[Switch.scala 30:53:@9799.4]
  wire  valid_30_43; // @[Switch.scala 30:36:@9800.4]
  wire  _T_29336; // @[Switch.scala 30:53:@9802.4]
  wire  valid_30_44; // @[Switch.scala 30:36:@9803.4]
  wire  _T_29339; // @[Switch.scala 30:53:@9805.4]
  wire  valid_30_45; // @[Switch.scala 30:36:@9806.4]
  wire  _T_29342; // @[Switch.scala 30:53:@9808.4]
  wire  valid_30_46; // @[Switch.scala 30:36:@9809.4]
  wire  _T_29345; // @[Switch.scala 30:53:@9811.4]
  wire  valid_30_47; // @[Switch.scala 30:36:@9812.4]
  wire  _T_29348; // @[Switch.scala 30:53:@9814.4]
  wire  valid_30_48; // @[Switch.scala 30:36:@9815.4]
  wire  _T_29351; // @[Switch.scala 30:53:@9817.4]
  wire  valid_30_49; // @[Switch.scala 30:36:@9818.4]
  wire  _T_29354; // @[Switch.scala 30:53:@9820.4]
  wire  valid_30_50; // @[Switch.scala 30:36:@9821.4]
  wire  _T_29357; // @[Switch.scala 30:53:@9823.4]
  wire  valid_30_51; // @[Switch.scala 30:36:@9824.4]
  wire  _T_29360; // @[Switch.scala 30:53:@9826.4]
  wire  valid_30_52; // @[Switch.scala 30:36:@9827.4]
  wire  _T_29363; // @[Switch.scala 30:53:@9829.4]
  wire  valid_30_53; // @[Switch.scala 30:36:@9830.4]
  wire  _T_29366; // @[Switch.scala 30:53:@9832.4]
  wire  valid_30_54; // @[Switch.scala 30:36:@9833.4]
  wire  _T_29369; // @[Switch.scala 30:53:@9835.4]
  wire  valid_30_55; // @[Switch.scala 30:36:@9836.4]
  wire  _T_29372; // @[Switch.scala 30:53:@9838.4]
  wire  valid_30_56; // @[Switch.scala 30:36:@9839.4]
  wire  _T_29375; // @[Switch.scala 30:53:@9841.4]
  wire  valid_30_57; // @[Switch.scala 30:36:@9842.4]
  wire  _T_29378; // @[Switch.scala 30:53:@9844.4]
  wire  valid_30_58; // @[Switch.scala 30:36:@9845.4]
  wire  _T_29381; // @[Switch.scala 30:53:@9847.4]
  wire  valid_30_59; // @[Switch.scala 30:36:@9848.4]
  wire  _T_29384; // @[Switch.scala 30:53:@9850.4]
  wire  valid_30_60; // @[Switch.scala 30:36:@9851.4]
  wire  _T_29387; // @[Switch.scala 30:53:@9853.4]
  wire  valid_30_61; // @[Switch.scala 30:36:@9854.4]
  wire  _T_29390; // @[Switch.scala 30:53:@9856.4]
  wire  valid_30_62; // @[Switch.scala 30:36:@9857.4]
  wire  _T_29393; // @[Switch.scala 30:53:@9859.4]
  wire  valid_30_63; // @[Switch.scala 30:36:@9860.4]
  wire [5:0] _T_29459; // @[Mux.scala 31:69:@9862.4]
  wire [5:0] _T_29460; // @[Mux.scala 31:69:@9863.4]
  wire [5:0] _T_29461; // @[Mux.scala 31:69:@9864.4]
  wire [5:0] _T_29462; // @[Mux.scala 31:69:@9865.4]
  wire [5:0] _T_29463; // @[Mux.scala 31:69:@9866.4]
  wire [5:0] _T_29464; // @[Mux.scala 31:69:@9867.4]
  wire [5:0] _T_29465; // @[Mux.scala 31:69:@9868.4]
  wire [5:0] _T_29466; // @[Mux.scala 31:69:@9869.4]
  wire [5:0] _T_29467; // @[Mux.scala 31:69:@9870.4]
  wire [5:0] _T_29468; // @[Mux.scala 31:69:@9871.4]
  wire [5:0] _T_29469; // @[Mux.scala 31:69:@9872.4]
  wire [5:0] _T_29470; // @[Mux.scala 31:69:@9873.4]
  wire [5:0] _T_29471; // @[Mux.scala 31:69:@9874.4]
  wire [5:0] _T_29472; // @[Mux.scala 31:69:@9875.4]
  wire [5:0] _T_29473; // @[Mux.scala 31:69:@9876.4]
  wire [5:0] _T_29474; // @[Mux.scala 31:69:@9877.4]
  wire [5:0] _T_29475; // @[Mux.scala 31:69:@9878.4]
  wire [5:0] _T_29476; // @[Mux.scala 31:69:@9879.4]
  wire [5:0] _T_29477; // @[Mux.scala 31:69:@9880.4]
  wire [5:0] _T_29478; // @[Mux.scala 31:69:@9881.4]
  wire [5:0] _T_29479; // @[Mux.scala 31:69:@9882.4]
  wire [5:0] _T_29480; // @[Mux.scala 31:69:@9883.4]
  wire [5:0] _T_29481; // @[Mux.scala 31:69:@9884.4]
  wire [5:0] _T_29482; // @[Mux.scala 31:69:@9885.4]
  wire [5:0] _T_29483; // @[Mux.scala 31:69:@9886.4]
  wire [5:0] _T_29484; // @[Mux.scala 31:69:@9887.4]
  wire [5:0] _T_29485; // @[Mux.scala 31:69:@9888.4]
  wire [5:0] _T_29486; // @[Mux.scala 31:69:@9889.4]
  wire [5:0] _T_29487; // @[Mux.scala 31:69:@9890.4]
  wire [5:0] _T_29488; // @[Mux.scala 31:69:@9891.4]
  wire [5:0] _T_29489; // @[Mux.scala 31:69:@9892.4]
  wire [5:0] _T_29490; // @[Mux.scala 31:69:@9893.4]
  wire [5:0] _T_29491; // @[Mux.scala 31:69:@9894.4]
  wire [5:0] _T_29492; // @[Mux.scala 31:69:@9895.4]
  wire [5:0] _T_29493; // @[Mux.scala 31:69:@9896.4]
  wire [5:0] _T_29494; // @[Mux.scala 31:69:@9897.4]
  wire [5:0] _T_29495; // @[Mux.scala 31:69:@9898.4]
  wire [5:0] _T_29496; // @[Mux.scala 31:69:@9899.4]
  wire [5:0] _T_29497; // @[Mux.scala 31:69:@9900.4]
  wire [5:0] _T_29498; // @[Mux.scala 31:69:@9901.4]
  wire [5:0] _T_29499; // @[Mux.scala 31:69:@9902.4]
  wire [5:0] _T_29500; // @[Mux.scala 31:69:@9903.4]
  wire [5:0] _T_29501; // @[Mux.scala 31:69:@9904.4]
  wire [5:0] _T_29502; // @[Mux.scala 31:69:@9905.4]
  wire [5:0] _T_29503; // @[Mux.scala 31:69:@9906.4]
  wire [5:0] _T_29504; // @[Mux.scala 31:69:@9907.4]
  wire [5:0] _T_29505; // @[Mux.scala 31:69:@9908.4]
  wire [5:0] _T_29506; // @[Mux.scala 31:69:@9909.4]
  wire [5:0] _T_29507; // @[Mux.scala 31:69:@9910.4]
  wire [5:0] _T_29508; // @[Mux.scala 31:69:@9911.4]
  wire [5:0] _T_29509; // @[Mux.scala 31:69:@9912.4]
  wire [5:0] _T_29510; // @[Mux.scala 31:69:@9913.4]
  wire [5:0] _T_29511; // @[Mux.scala 31:69:@9914.4]
  wire [5:0] _T_29512; // @[Mux.scala 31:69:@9915.4]
  wire [5:0] _T_29513; // @[Mux.scala 31:69:@9916.4]
  wire [5:0] _T_29514; // @[Mux.scala 31:69:@9917.4]
  wire [5:0] _T_29515; // @[Mux.scala 31:69:@9918.4]
  wire [5:0] _T_29516; // @[Mux.scala 31:69:@9919.4]
  wire [5:0] _T_29517; // @[Mux.scala 31:69:@9920.4]
  wire [5:0] _T_29518; // @[Mux.scala 31:69:@9921.4]
  wire [5:0] _T_29519; // @[Mux.scala 31:69:@9922.4]
  wire [5:0] _T_29520; // @[Mux.scala 31:69:@9923.4]
  wire [5:0] select_30; // @[Mux.scala 31:69:@9924.4]
  wire [47:0] _GEN_1921; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1922; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1923; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1924; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1925; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1926; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1927; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1928; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1929; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1930; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1931; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1932; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1933; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1934; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1935; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1936; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1937; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1938; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1939; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1940; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1941; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1942; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1943; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1944; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1945; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1946; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1947; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1948; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1949; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1950; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1951; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1952; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1953; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1954; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1955; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1956; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1957; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1958; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1959; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1960; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1961; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1962; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1963; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1964; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1965; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1966; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1967; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1968; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1969; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1970; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1971; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1972; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1973; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1974; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1975; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1976; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1977; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1978; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1979; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1980; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1981; // @[Switch.scala 33:19:@9926.4]
  wire [47:0] _GEN_1982; // @[Switch.scala 33:19:@9926.4]
  wire [7:0] _T_29529; // @[Switch.scala 34:32:@9933.4]
  wire [15:0] _T_29537; // @[Switch.scala 34:32:@9941.4]
  wire [7:0] _T_29544; // @[Switch.scala 34:32:@9948.4]
  wire [31:0] _T_29553; // @[Switch.scala 34:32:@9957.4]
  wire [7:0] _T_29560; // @[Switch.scala 34:32:@9964.4]
  wire [15:0] _T_29568; // @[Switch.scala 34:32:@9972.4]
  wire [7:0] _T_29575; // @[Switch.scala 34:32:@9979.4]
  wire [31:0] _T_29584; // @[Switch.scala 34:32:@9988.4]
  wire [63:0] _T_29585; // @[Switch.scala 34:32:@9989.4]
  wire  _T_29589; // @[Switch.scala 30:53:@9992.4]
  wire  valid_31_0; // @[Switch.scala 30:36:@9993.4]
  wire  _T_29592; // @[Switch.scala 30:53:@9995.4]
  wire  valid_31_1; // @[Switch.scala 30:36:@9996.4]
  wire  _T_29595; // @[Switch.scala 30:53:@9998.4]
  wire  valid_31_2; // @[Switch.scala 30:36:@9999.4]
  wire  _T_29598; // @[Switch.scala 30:53:@10001.4]
  wire  valid_31_3; // @[Switch.scala 30:36:@10002.4]
  wire  _T_29601; // @[Switch.scala 30:53:@10004.4]
  wire  valid_31_4; // @[Switch.scala 30:36:@10005.4]
  wire  _T_29604; // @[Switch.scala 30:53:@10007.4]
  wire  valid_31_5; // @[Switch.scala 30:36:@10008.4]
  wire  _T_29607; // @[Switch.scala 30:53:@10010.4]
  wire  valid_31_6; // @[Switch.scala 30:36:@10011.4]
  wire  _T_29610; // @[Switch.scala 30:53:@10013.4]
  wire  valid_31_7; // @[Switch.scala 30:36:@10014.4]
  wire  _T_29613; // @[Switch.scala 30:53:@10016.4]
  wire  valid_31_8; // @[Switch.scala 30:36:@10017.4]
  wire  _T_29616; // @[Switch.scala 30:53:@10019.4]
  wire  valid_31_9; // @[Switch.scala 30:36:@10020.4]
  wire  _T_29619; // @[Switch.scala 30:53:@10022.4]
  wire  valid_31_10; // @[Switch.scala 30:36:@10023.4]
  wire  _T_29622; // @[Switch.scala 30:53:@10025.4]
  wire  valid_31_11; // @[Switch.scala 30:36:@10026.4]
  wire  _T_29625; // @[Switch.scala 30:53:@10028.4]
  wire  valid_31_12; // @[Switch.scala 30:36:@10029.4]
  wire  _T_29628; // @[Switch.scala 30:53:@10031.4]
  wire  valid_31_13; // @[Switch.scala 30:36:@10032.4]
  wire  _T_29631; // @[Switch.scala 30:53:@10034.4]
  wire  valid_31_14; // @[Switch.scala 30:36:@10035.4]
  wire  _T_29634; // @[Switch.scala 30:53:@10037.4]
  wire  valid_31_15; // @[Switch.scala 30:36:@10038.4]
  wire  _T_29637; // @[Switch.scala 30:53:@10040.4]
  wire  valid_31_16; // @[Switch.scala 30:36:@10041.4]
  wire  _T_29640; // @[Switch.scala 30:53:@10043.4]
  wire  valid_31_17; // @[Switch.scala 30:36:@10044.4]
  wire  _T_29643; // @[Switch.scala 30:53:@10046.4]
  wire  valid_31_18; // @[Switch.scala 30:36:@10047.4]
  wire  _T_29646; // @[Switch.scala 30:53:@10049.4]
  wire  valid_31_19; // @[Switch.scala 30:36:@10050.4]
  wire  _T_29649; // @[Switch.scala 30:53:@10052.4]
  wire  valid_31_20; // @[Switch.scala 30:36:@10053.4]
  wire  _T_29652; // @[Switch.scala 30:53:@10055.4]
  wire  valid_31_21; // @[Switch.scala 30:36:@10056.4]
  wire  _T_29655; // @[Switch.scala 30:53:@10058.4]
  wire  valid_31_22; // @[Switch.scala 30:36:@10059.4]
  wire  _T_29658; // @[Switch.scala 30:53:@10061.4]
  wire  valid_31_23; // @[Switch.scala 30:36:@10062.4]
  wire  _T_29661; // @[Switch.scala 30:53:@10064.4]
  wire  valid_31_24; // @[Switch.scala 30:36:@10065.4]
  wire  _T_29664; // @[Switch.scala 30:53:@10067.4]
  wire  valid_31_25; // @[Switch.scala 30:36:@10068.4]
  wire  _T_29667; // @[Switch.scala 30:53:@10070.4]
  wire  valid_31_26; // @[Switch.scala 30:36:@10071.4]
  wire  _T_29670; // @[Switch.scala 30:53:@10073.4]
  wire  valid_31_27; // @[Switch.scala 30:36:@10074.4]
  wire  _T_29673; // @[Switch.scala 30:53:@10076.4]
  wire  valid_31_28; // @[Switch.scala 30:36:@10077.4]
  wire  _T_29676; // @[Switch.scala 30:53:@10079.4]
  wire  valid_31_29; // @[Switch.scala 30:36:@10080.4]
  wire  _T_29679; // @[Switch.scala 30:53:@10082.4]
  wire  valid_31_30; // @[Switch.scala 30:36:@10083.4]
  wire  _T_29682; // @[Switch.scala 30:53:@10085.4]
  wire  valid_31_31; // @[Switch.scala 30:36:@10086.4]
  wire  _T_29685; // @[Switch.scala 30:53:@10088.4]
  wire  valid_31_32; // @[Switch.scala 30:36:@10089.4]
  wire  _T_29688; // @[Switch.scala 30:53:@10091.4]
  wire  valid_31_33; // @[Switch.scala 30:36:@10092.4]
  wire  _T_29691; // @[Switch.scala 30:53:@10094.4]
  wire  valid_31_34; // @[Switch.scala 30:36:@10095.4]
  wire  _T_29694; // @[Switch.scala 30:53:@10097.4]
  wire  valid_31_35; // @[Switch.scala 30:36:@10098.4]
  wire  _T_29697; // @[Switch.scala 30:53:@10100.4]
  wire  valid_31_36; // @[Switch.scala 30:36:@10101.4]
  wire  _T_29700; // @[Switch.scala 30:53:@10103.4]
  wire  valid_31_37; // @[Switch.scala 30:36:@10104.4]
  wire  _T_29703; // @[Switch.scala 30:53:@10106.4]
  wire  valid_31_38; // @[Switch.scala 30:36:@10107.4]
  wire  _T_29706; // @[Switch.scala 30:53:@10109.4]
  wire  valid_31_39; // @[Switch.scala 30:36:@10110.4]
  wire  _T_29709; // @[Switch.scala 30:53:@10112.4]
  wire  valid_31_40; // @[Switch.scala 30:36:@10113.4]
  wire  _T_29712; // @[Switch.scala 30:53:@10115.4]
  wire  valid_31_41; // @[Switch.scala 30:36:@10116.4]
  wire  _T_29715; // @[Switch.scala 30:53:@10118.4]
  wire  valid_31_42; // @[Switch.scala 30:36:@10119.4]
  wire  _T_29718; // @[Switch.scala 30:53:@10121.4]
  wire  valid_31_43; // @[Switch.scala 30:36:@10122.4]
  wire  _T_29721; // @[Switch.scala 30:53:@10124.4]
  wire  valid_31_44; // @[Switch.scala 30:36:@10125.4]
  wire  _T_29724; // @[Switch.scala 30:53:@10127.4]
  wire  valid_31_45; // @[Switch.scala 30:36:@10128.4]
  wire  _T_29727; // @[Switch.scala 30:53:@10130.4]
  wire  valid_31_46; // @[Switch.scala 30:36:@10131.4]
  wire  _T_29730; // @[Switch.scala 30:53:@10133.4]
  wire  valid_31_47; // @[Switch.scala 30:36:@10134.4]
  wire  _T_29733; // @[Switch.scala 30:53:@10136.4]
  wire  valid_31_48; // @[Switch.scala 30:36:@10137.4]
  wire  _T_29736; // @[Switch.scala 30:53:@10139.4]
  wire  valid_31_49; // @[Switch.scala 30:36:@10140.4]
  wire  _T_29739; // @[Switch.scala 30:53:@10142.4]
  wire  valid_31_50; // @[Switch.scala 30:36:@10143.4]
  wire  _T_29742; // @[Switch.scala 30:53:@10145.4]
  wire  valid_31_51; // @[Switch.scala 30:36:@10146.4]
  wire  _T_29745; // @[Switch.scala 30:53:@10148.4]
  wire  valid_31_52; // @[Switch.scala 30:36:@10149.4]
  wire  _T_29748; // @[Switch.scala 30:53:@10151.4]
  wire  valid_31_53; // @[Switch.scala 30:36:@10152.4]
  wire  _T_29751; // @[Switch.scala 30:53:@10154.4]
  wire  valid_31_54; // @[Switch.scala 30:36:@10155.4]
  wire  _T_29754; // @[Switch.scala 30:53:@10157.4]
  wire  valid_31_55; // @[Switch.scala 30:36:@10158.4]
  wire  _T_29757; // @[Switch.scala 30:53:@10160.4]
  wire  valid_31_56; // @[Switch.scala 30:36:@10161.4]
  wire  _T_29760; // @[Switch.scala 30:53:@10163.4]
  wire  valid_31_57; // @[Switch.scala 30:36:@10164.4]
  wire  _T_29763; // @[Switch.scala 30:53:@10166.4]
  wire  valid_31_58; // @[Switch.scala 30:36:@10167.4]
  wire  _T_29766; // @[Switch.scala 30:53:@10169.4]
  wire  valid_31_59; // @[Switch.scala 30:36:@10170.4]
  wire  _T_29769; // @[Switch.scala 30:53:@10172.4]
  wire  valid_31_60; // @[Switch.scala 30:36:@10173.4]
  wire  _T_29772; // @[Switch.scala 30:53:@10175.4]
  wire  valid_31_61; // @[Switch.scala 30:36:@10176.4]
  wire  _T_29775; // @[Switch.scala 30:53:@10178.4]
  wire  valid_31_62; // @[Switch.scala 30:36:@10179.4]
  wire  _T_29778; // @[Switch.scala 30:53:@10181.4]
  wire  valid_31_63; // @[Switch.scala 30:36:@10182.4]
  wire [5:0] _T_29844; // @[Mux.scala 31:69:@10184.4]
  wire [5:0] _T_29845; // @[Mux.scala 31:69:@10185.4]
  wire [5:0] _T_29846; // @[Mux.scala 31:69:@10186.4]
  wire [5:0] _T_29847; // @[Mux.scala 31:69:@10187.4]
  wire [5:0] _T_29848; // @[Mux.scala 31:69:@10188.4]
  wire [5:0] _T_29849; // @[Mux.scala 31:69:@10189.4]
  wire [5:0] _T_29850; // @[Mux.scala 31:69:@10190.4]
  wire [5:0] _T_29851; // @[Mux.scala 31:69:@10191.4]
  wire [5:0] _T_29852; // @[Mux.scala 31:69:@10192.4]
  wire [5:0] _T_29853; // @[Mux.scala 31:69:@10193.4]
  wire [5:0] _T_29854; // @[Mux.scala 31:69:@10194.4]
  wire [5:0] _T_29855; // @[Mux.scala 31:69:@10195.4]
  wire [5:0] _T_29856; // @[Mux.scala 31:69:@10196.4]
  wire [5:0] _T_29857; // @[Mux.scala 31:69:@10197.4]
  wire [5:0] _T_29858; // @[Mux.scala 31:69:@10198.4]
  wire [5:0] _T_29859; // @[Mux.scala 31:69:@10199.4]
  wire [5:0] _T_29860; // @[Mux.scala 31:69:@10200.4]
  wire [5:0] _T_29861; // @[Mux.scala 31:69:@10201.4]
  wire [5:0] _T_29862; // @[Mux.scala 31:69:@10202.4]
  wire [5:0] _T_29863; // @[Mux.scala 31:69:@10203.4]
  wire [5:0] _T_29864; // @[Mux.scala 31:69:@10204.4]
  wire [5:0] _T_29865; // @[Mux.scala 31:69:@10205.4]
  wire [5:0] _T_29866; // @[Mux.scala 31:69:@10206.4]
  wire [5:0] _T_29867; // @[Mux.scala 31:69:@10207.4]
  wire [5:0] _T_29868; // @[Mux.scala 31:69:@10208.4]
  wire [5:0] _T_29869; // @[Mux.scala 31:69:@10209.4]
  wire [5:0] _T_29870; // @[Mux.scala 31:69:@10210.4]
  wire [5:0] _T_29871; // @[Mux.scala 31:69:@10211.4]
  wire [5:0] _T_29872; // @[Mux.scala 31:69:@10212.4]
  wire [5:0] _T_29873; // @[Mux.scala 31:69:@10213.4]
  wire [5:0] _T_29874; // @[Mux.scala 31:69:@10214.4]
  wire [5:0] _T_29875; // @[Mux.scala 31:69:@10215.4]
  wire [5:0] _T_29876; // @[Mux.scala 31:69:@10216.4]
  wire [5:0] _T_29877; // @[Mux.scala 31:69:@10217.4]
  wire [5:0] _T_29878; // @[Mux.scala 31:69:@10218.4]
  wire [5:0] _T_29879; // @[Mux.scala 31:69:@10219.4]
  wire [5:0] _T_29880; // @[Mux.scala 31:69:@10220.4]
  wire [5:0] _T_29881; // @[Mux.scala 31:69:@10221.4]
  wire [5:0] _T_29882; // @[Mux.scala 31:69:@10222.4]
  wire [5:0] _T_29883; // @[Mux.scala 31:69:@10223.4]
  wire [5:0] _T_29884; // @[Mux.scala 31:69:@10224.4]
  wire [5:0] _T_29885; // @[Mux.scala 31:69:@10225.4]
  wire [5:0] _T_29886; // @[Mux.scala 31:69:@10226.4]
  wire [5:0] _T_29887; // @[Mux.scala 31:69:@10227.4]
  wire [5:0] _T_29888; // @[Mux.scala 31:69:@10228.4]
  wire [5:0] _T_29889; // @[Mux.scala 31:69:@10229.4]
  wire [5:0] _T_29890; // @[Mux.scala 31:69:@10230.4]
  wire [5:0] _T_29891; // @[Mux.scala 31:69:@10231.4]
  wire [5:0] _T_29892; // @[Mux.scala 31:69:@10232.4]
  wire [5:0] _T_29893; // @[Mux.scala 31:69:@10233.4]
  wire [5:0] _T_29894; // @[Mux.scala 31:69:@10234.4]
  wire [5:0] _T_29895; // @[Mux.scala 31:69:@10235.4]
  wire [5:0] _T_29896; // @[Mux.scala 31:69:@10236.4]
  wire [5:0] _T_29897; // @[Mux.scala 31:69:@10237.4]
  wire [5:0] _T_29898; // @[Mux.scala 31:69:@10238.4]
  wire [5:0] _T_29899; // @[Mux.scala 31:69:@10239.4]
  wire [5:0] _T_29900; // @[Mux.scala 31:69:@10240.4]
  wire [5:0] _T_29901; // @[Mux.scala 31:69:@10241.4]
  wire [5:0] _T_29902; // @[Mux.scala 31:69:@10242.4]
  wire [5:0] _T_29903; // @[Mux.scala 31:69:@10243.4]
  wire [5:0] _T_29904; // @[Mux.scala 31:69:@10244.4]
  wire [5:0] _T_29905; // @[Mux.scala 31:69:@10245.4]
  wire [5:0] select_31; // @[Mux.scala 31:69:@10246.4]
  wire [47:0] _GEN_1985; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_1986; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_1987; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_1988; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_1989; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_1990; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_1991; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_1992; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_1993; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_1994; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_1995; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_1996; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_1997; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_1998; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_1999; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2000; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2001; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2002; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2003; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2004; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2005; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2006; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2007; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2008; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2009; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2010; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2011; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2012; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2013; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2014; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2015; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2016; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2017; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2018; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2019; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2020; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2021; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2022; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2023; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2024; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2025; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2026; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2027; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2028; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2029; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2030; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2031; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2032; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2033; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2034; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2035; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2036; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2037; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2038; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2039; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2040; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2041; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2042; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2043; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2044; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2045; // @[Switch.scala 33:19:@10248.4]
  wire [47:0] _GEN_2046; // @[Switch.scala 33:19:@10248.4]
  wire [7:0] _T_29914; // @[Switch.scala 34:32:@10255.4]
  wire [15:0] _T_29922; // @[Switch.scala 34:32:@10263.4]
  wire [7:0] _T_29929; // @[Switch.scala 34:32:@10270.4]
  wire [31:0] _T_29938; // @[Switch.scala 34:32:@10279.4]
  wire [7:0] _T_29945; // @[Switch.scala 34:32:@10286.4]
  wire [15:0] _T_29953; // @[Switch.scala 34:32:@10294.4]
  wire [7:0] _T_29960; // @[Switch.scala 34:32:@10301.4]
  wire [31:0] _T_29969; // @[Switch.scala 34:32:@10310.4]
  wire [63:0] _T_29970; // @[Switch.scala 34:32:@10311.4]
  wire  _T_29974; // @[Switch.scala 30:53:@10314.4]
  wire  valid_32_0; // @[Switch.scala 30:36:@10315.4]
  wire  _T_29977; // @[Switch.scala 30:53:@10317.4]
  wire  valid_32_1; // @[Switch.scala 30:36:@10318.4]
  wire  _T_29980; // @[Switch.scala 30:53:@10320.4]
  wire  valid_32_2; // @[Switch.scala 30:36:@10321.4]
  wire  _T_29983; // @[Switch.scala 30:53:@10323.4]
  wire  valid_32_3; // @[Switch.scala 30:36:@10324.4]
  wire  _T_29986; // @[Switch.scala 30:53:@10326.4]
  wire  valid_32_4; // @[Switch.scala 30:36:@10327.4]
  wire  _T_29989; // @[Switch.scala 30:53:@10329.4]
  wire  valid_32_5; // @[Switch.scala 30:36:@10330.4]
  wire  _T_29992; // @[Switch.scala 30:53:@10332.4]
  wire  valid_32_6; // @[Switch.scala 30:36:@10333.4]
  wire  _T_29995; // @[Switch.scala 30:53:@10335.4]
  wire  valid_32_7; // @[Switch.scala 30:36:@10336.4]
  wire  _T_29998; // @[Switch.scala 30:53:@10338.4]
  wire  valid_32_8; // @[Switch.scala 30:36:@10339.4]
  wire  _T_30001; // @[Switch.scala 30:53:@10341.4]
  wire  valid_32_9; // @[Switch.scala 30:36:@10342.4]
  wire  _T_30004; // @[Switch.scala 30:53:@10344.4]
  wire  valid_32_10; // @[Switch.scala 30:36:@10345.4]
  wire  _T_30007; // @[Switch.scala 30:53:@10347.4]
  wire  valid_32_11; // @[Switch.scala 30:36:@10348.4]
  wire  _T_30010; // @[Switch.scala 30:53:@10350.4]
  wire  valid_32_12; // @[Switch.scala 30:36:@10351.4]
  wire  _T_30013; // @[Switch.scala 30:53:@10353.4]
  wire  valid_32_13; // @[Switch.scala 30:36:@10354.4]
  wire  _T_30016; // @[Switch.scala 30:53:@10356.4]
  wire  valid_32_14; // @[Switch.scala 30:36:@10357.4]
  wire  _T_30019; // @[Switch.scala 30:53:@10359.4]
  wire  valid_32_15; // @[Switch.scala 30:36:@10360.4]
  wire  _T_30022; // @[Switch.scala 30:53:@10362.4]
  wire  valid_32_16; // @[Switch.scala 30:36:@10363.4]
  wire  _T_30025; // @[Switch.scala 30:53:@10365.4]
  wire  valid_32_17; // @[Switch.scala 30:36:@10366.4]
  wire  _T_30028; // @[Switch.scala 30:53:@10368.4]
  wire  valid_32_18; // @[Switch.scala 30:36:@10369.4]
  wire  _T_30031; // @[Switch.scala 30:53:@10371.4]
  wire  valid_32_19; // @[Switch.scala 30:36:@10372.4]
  wire  _T_30034; // @[Switch.scala 30:53:@10374.4]
  wire  valid_32_20; // @[Switch.scala 30:36:@10375.4]
  wire  _T_30037; // @[Switch.scala 30:53:@10377.4]
  wire  valid_32_21; // @[Switch.scala 30:36:@10378.4]
  wire  _T_30040; // @[Switch.scala 30:53:@10380.4]
  wire  valid_32_22; // @[Switch.scala 30:36:@10381.4]
  wire  _T_30043; // @[Switch.scala 30:53:@10383.4]
  wire  valid_32_23; // @[Switch.scala 30:36:@10384.4]
  wire  _T_30046; // @[Switch.scala 30:53:@10386.4]
  wire  valid_32_24; // @[Switch.scala 30:36:@10387.4]
  wire  _T_30049; // @[Switch.scala 30:53:@10389.4]
  wire  valid_32_25; // @[Switch.scala 30:36:@10390.4]
  wire  _T_30052; // @[Switch.scala 30:53:@10392.4]
  wire  valid_32_26; // @[Switch.scala 30:36:@10393.4]
  wire  _T_30055; // @[Switch.scala 30:53:@10395.4]
  wire  valid_32_27; // @[Switch.scala 30:36:@10396.4]
  wire  _T_30058; // @[Switch.scala 30:53:@10398.4]
  wire  valid_32_28; // @[Switch.scala 30:36:@10399.4]
  wire  _T_30061; // @[Switch.scala 30:53:@10401.4]
  wire  valid_32_29; // @[Switch.scala 30:36:@10402.4]
  wire  _T_30064; // @[Switch.scala 30:53:@10404.4]
  wire  valid_32_30; // @[Switch.scala 30:36:@10405.4]
  wire  _T_30067; // @[Switch.scala 30:53:@10407.4]
  wire  valid_32_31; // @[Switch.scala 30:36:@10408.4]
  wire  _T_30070; // @[Switch.scala 30:53:@10410.4]
  wire  valid_32_32; // @[Switch.scala 30:36:@10411.4]
  wire  _T_30073; // @[Switch.scala 30:53:@10413.4]
  wire  valid_32_33; // @[Switch.scala 30:36:@10414.4]
  wire  _T_30076; // @[Switch.scala 30:53:@10416.4]
  wire  valid_32_34; // @[Switch.scala 30:36:@10417.4]
  wire  _T_30079; // @[Switch.scala 30:53:@10419.4]
  wire  valid_32_35; // @[Switch.scala 30:36:@10420.4]
  wire  _T_30082; // @[Switch.scala 30:53:@10422.4]
  wire  valid_32_36; // @[Switch.scala 30:36:@10423.4]
  wire  _T_30085; // @[Switch.scala 30:53:@10425.4]
  wire  valid_32_37; // @[Switch.scala 30:36:@10426.4]
  wire  _T_30088; // @[Switch.scala 30:53:@10428.4]
  wire  valid_32_38; // @[Switch.scala 30:36:@10429.4]
  wire  _T_30091; // @[Switch.scala 30:53:@10431.4]
  wire  valid_32_39; // @[Switch.scala 30:36:@10432.4]
  wire  _T_30094; // @[Switch.scala 30:53:@10434.4]
  wire  valid_32_40; // @[Switch.scala 30:36:@10435.4]
  wire  _T_30097; // @[Switch.scala 30:53:@10437.4]
  wire  valid_32_41; // @[Switch.scala 30:36:@10438.4]
  wire  _T_30100; // @[Switch.scala 30:53:@10440.4]
  wire  valid_32_42; // @[Switch.scala 30:36:@10441.4]
  wire  _T_30103; // @[Switch.scala 30:53:@10443.4]
  wire  valid_32_43; // @[Switch.scala 30:36:@10444.4]
  wire  _T_30106; // @[Switch.scala 30:53:@10446.4]
  wire  valid_32_44; // @[Switch.scala 30:36:@10447.4]
  wire  _T_30109; // @[Switch.scala 30:53:@10449.4]
  wire  valid_32_45; // @[Switch.scala 30:36:@10450.4]
  wire  _T_30112; // @[Switch.scala 30:53:@10452.4]
  wire  valid_32_46; // @[Switch.scala 30:36:@10453.4]
  wire  _T_30115; // @[Switch.scala 30:53:@10455.4]
  wire  valid_32_47; // @[Switch.scala 30:36:@10456.4]
  wire  _T_30118; // @[Switch.scala 30:53:@10458.4]
  wire  valid_32_48; // @[Switch.scala 30:36:@10459.4]
  wire  _T_30121; // @[Switch.scala 30:53:@10461.4]
  wire  valid_32_49; // @[Switch.scala 30:36:@10462.4]
  wire  _T_30124; // @[Switch.scala 30:53:@10464.4]
  wire  valid_32_50; // @[Switch.scala 30:36:@10465.4]
  wire  _T_30127; // @[Switch.scala 30:53:@10467.4]
  wire  valid_32_51; // @[Switch.scala 30:36:@10468.4]
  wire  _T_30130; // @[Switch.scala 30:53:@10470.4]
  wire  valid_32_52; // @[Switch.scala 30:36:@10471.4]
  wire  _T_30133; // @[Switch.scala 30:53:@10473.4]
  wire  valid_32_53; // @[Switch.scala 30:36:@10474.4]
  wire  _T_30136; // @[Switch.scala 30:53:@10476.4]
  wire  valid_32_54; // @[Switch.scala 30:36:@10477.4]
  wire  _T_30139; // @[Switch.scala 30:53:@10479.4]
  wire  valid_32_55; // @[Switch.scala 30:36:@10480.4]
  wire  _T_30142; // @[Switch.scala 30:53:@10482.4]
  wire  valid_32_56; // @[Switch.scala 30:36:@10483.4]
  wire  _T_30145; // @[Switch.scala 30:53:@10485.4]
  wire  valid_32_57; // @[Switch.scala 30:36:@10486.4]
  wire  _T_30148; // @[Switch.scala 30:53:@10488.4]
  wire  valid_32_58; // @[Switch.scala 30:36:@10489.4]
  wire  _T_30151; // @[Switch.scala 30:53:@10491.4]
  wire  valid_32_59; // @[Switch.scala 30:36:@10492.4]
  wire  _T_30154; // @[Switch.scala 30:53:@10494.4]
  wire  valid_32_60; // @[Switch.scala 30:36:@10495.4]
  wire  _T_30157; // @[Switch.scala 30:53:@10497.4]
  wire  valid_32_61; // @[Switch.scala 30:36:@10498.4]
  wire  _T_30160; // @[Switch.scala 30:53:@10500.4]
  wire  valid_32_62; // @[Switch.scala 30:36:@10501.4]
  wire  _T_30163; // @[Switch.scala 30:53:@10503.4]
  wire  valid_32_63; // @[Switch.scala 30:36:@10504.4]
  wire [5:0] _T_30229; // @[Mux.scala 31:69:@10506.4]
  wire [5:0] _T_30230; // @[Mux.scala 31:69:@10507.4]
  wire [5:0] _T_30231; // @[Mux.scala 31:69:@10508.4]
  wire [5:0] _T_30232; // @[Mux.scala 31:69:@10509.4]
  wire [5:0] _T_30233; // @[Mux.scala 31:69:@10510.4]
  wire [5:0] _T_30234; // @[Mux.scala 31:69:@10511.4]
  wire [5:0] _T_30235; // @[Mux.scala 31:69:@10512.4]
  wire [5:0] _T_30236; // @[Mux.scala 31:69:@10513.4]
  wire [5:0] _T_30237; // @[Mux.scala 31:69:@10514.4]
  wire [5:0] _T_30238; // @[Mux.scala 31:69:@10515.4]
  wire [5:0] _T_30239; // @[Mux.scala 31:69:@10516.4]
  wire [5:0] _T_30240; // @[Mux.scala 31:69:@10517.4]
  wire [5:0] _T_30241; // @[Mux.scala 31:69:@10518.4]
  wire [5:0] _T_30242; // @[Mux.scala 31:69:@10519.4]
  wire [5:0] _T_30243; // @[Mux.scala 31:69:@10520.4]
  wire [5:0] _T_30244; // @[Mux.scala 31:69:@10521.4]
  wire [5:0] _T_30245; // @[Mux.scala 31:69:@10522.4]
  wire [5:0] _T_30246; // @[Mux.scala 31:69:@10523.4]
  wire [5:0] _T_30247; // @[Mux.scala 31:69:@10524.4]
  wire [5:0] _T_30248; // @[Mux.scala 31:69:@10525.4]
  wire [5:0] _T_30249; // @[Mux.scala 31:69:@10526.4]
  wire [5:0] _T_30250; // @[Mux.scala 31:69:@10527.4]
  wire [5:0] _T_30251; // @[Mux.scala 31:69:@10528.4]
  wire [5:0] _T_30252; // @[Mux.scala 31:69:@10529.4]
  wire [5:0] _T_30253; // @[Mux.scala 31:69:@10530.4]
  wire [5:0] _T_30254; // @[Mux.scala 31:69:@10531.4]
  wire [5:0] _T_30255; // @[Mux.scala 31:69:@10532.4]
  wire [5:0] _T_30256; // @[Mux.scala 31:69:@10533.4]
  wire [5:0] _T_30257; // @[Mux.scala 31:69:@10534.4]
  wire [5:0] _T_30258; // @[Mux.scala 31:69:@10535.4]
  wire [5:0] _T_30259; // @[Mux.scala 31:69:@10536.4]
  wire [5:0] _T_30260; // @[Mux.scala 31:69:@10537.4]
  wire [5:0] _T_30261; // @[Mux.scala 31:69:@10538.4]
  wire [5:0] _T_30262; // @[Mux.scala 31:69:@10539.4]
  wire [5:0] _T_30263; // @[Mux.scala 31:69:@10540.4]
  wire [5:0] _T_30264; // @[Mux.scala 31:69:@10541.4]
  wire [5:0] _T_30265; // @[Mux.scala 31:69:@10542.4]
  wire [5:0] _T_30266; // @[Mux.scala 31:69:@10543.4]
  wire [5:0] _T_30267; // @[Mux.scala 31:69:@10544.4]
  wire [5:0] _T_30268; // @[Mux.scala 31:69:@10545.4]
  wire [5:0] _T_30269; // @[Mux.scala 31:69:@10546.4]
  wire [5:0] _T_30270; // @[Mux.scala 31:69:@10547.4]
  wire [5:0] _T_30271; // @[Mux.scala 31:69:@10548.4]
  wire [5:0] _T_30272; // @[Mux.scala 31:69:@10549.4]
  wire [5:0] _T_30273; // @[Mux.scala 31:69:@10550.4]
  wire [5:0] _T_30274; // @[Mux.scala 31:69:@10551.4]
  wire [5:0] _T_30275; // @[Mux.scala 31:69:@10552.4]
  wire [5:0] _T_30276; // @[Mux.scala 31:69:@10553.4]
  wire [5:0] _T_30277; // @[Mux.scala 31:69:@10554.4]
  wire [5:0] _T_30278; // @[Mux.scala 31:69:@10555.4]
  wire [5:0] _T_30279; // @[Mux.scala 31:69:@10556.4]
  wire [5:0] _T_30280; // @[Mux.scala 31:69:@10557.4]
  wire [5:0] _T_30281; // @[Mux.scala 31:69:@10558.4]
  wire [5:0] _T_30282; // @[Mux.scala 31:69:@10559.4]
  wire [5:0] _T_30283; // @[Mux.scala 31:69:@10560.4]
  wire [5:0] _T_30284; // @[Mux.scala 31:69:@10561.4]
  wire [5:0] _T_30285; // @[Mux.scala 31:69:@10562.4]
  wire [5:0] _T_30286; // @[Mux.scala 31:69:@10563.4]
  wire [5:0] _T_30287; // @[Mux.scala 31:69:@10564.4]
  wire [5:0] _T_30288; // @[Mux.scala 31:69:@10565.4]
  wire [5:0] _T_30289; // @[Mux.scala 31:69:@10566.4]
  wire [5:0] _T_30290; // @[Mux.scala 31:69:@10567.4]
  wire [5:0] select_32; // @[Mux.scala 31:69:@10568.4]
  wire [47:0] _GEN_2049; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2050; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2051; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2052; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2053; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2054; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2055; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2056; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2057; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2058; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2059; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2060; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2061; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2062; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2063; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2064; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2065; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2066; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2067; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2068; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2069; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2070; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2071; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2072; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2073; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2074; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2075; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2076; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2077; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2078; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2079; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2080; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2081; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2082; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2083; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2084; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2085; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2086; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2087; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2088; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2089; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2090; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2091; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2092; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2093; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2094; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2095; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2096; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2097; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2098; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2099; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2100; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2101; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2102; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2103; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2104; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2105; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2106; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2107; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2108; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2109; // @[Switch.scala 33:19:@10570.4]
  wire [47:0] _GEN_2110; // @[Switch.scala 33:19:@10570.4]
  wire [7:0] _T_30299; // @[Switch.scala 34:32:@10577.4]
  wire [15:0] _T_30307; // @[Switch.scala 34:32:@10585.4]
  wire [7:0] _T_30314; // @[Switch.scala 34:32:@10592.4]
  wire [31:0] _T_30323; // @[Switch.scala 34:32:@10601.4]
  wire [7:0] _T_30330; // @[Switch.scala 34:32:@10608.4]
  wire [15:0] _T_30338; // @[Switch.scala 34:32:@10616.4]
  wire [7:0] _T_30345; // @[Switch.scala 34:32:@10623.4]
  wire [31:0] _T_30354; // @[Switch.scala 34:32:@10632.4]
  wire [63:0] _T_30355; // @[Switch.scala 34:32:@10633.4]
  wire  _T_30359; // @[Switch.scala 30:53:@10636.4]
  wire  valid_33_0; // @[Switch.scala 30:36:@10637.4]
  wire  _T_30362; // @[Switch.scala 30:53:@10639.4]
  wire  valid_33_1; // @[Switch.scala 30:36:@10640.4]
  wire  _T_30365; // @[Switch.scala 30:53:@10642.4]
  wire  valid_33_2; // @[Switch.scala 30:36:@10643.4]
  wire  _T_30368; // @[Switch.scala 30:53:@10645.4]
  wire  valid_33_3; // @[Switch.scala 30:36:@10646.4]
  wire  _T_30371; // @[Switch.scala 30:53:@10648.4]
  wire  valid_33_4; // @[Switch.scala 30:36:@10649.4]
  wire  _T_30374; // @[Switch.scala 30:53:@10651.4]
  wire  valid_33_5; // @[Switch.scala 30:36:@10652.4]
  wire  _T_30377; // @[Switch.scala 30:53:@10654.4]
  wire  valid_33_6; // @[Switch.scala 30:36:@10655.4]
  wire  _T_30380; // @[Switch.scala 30:53:@10657.4]
  wire  valid_33_7; // @[Switch.scala 30:36:@10658.4]
  wire  _T_30383; // @[Switch.scala 30:53:@10660.4]
  wire  valid_33_8; // @[Switch.scala 30:36:@10661.4]
  wire  _T_30386; // @[Switch.scala 30:53:@10663.4]
  wire  valid_33_9; // @[Switch.scala 30:36:@10664.4]
  wire  _T_30389; // @[Switch.scala 30:53:@10666.4]
  wire  valid_33_10; // @[Switch.scala 30:36:@10667.4]
  wire  _T_30392; // @[Switch.scala 30:53:@10669.4]
  wire  valid_33_11; // @[Switch.scala 30:36:@10670.4]
  wire  _T_30395; // @[Switch.scala 30:53:@10672.4]
  wire  valid_33_12; // @[Switch.scala 30:36:@10673.4]
  wire  _T_30398; // @[Switch.scala 30:53:@10675.4]
  wire  valid_33_13; // @[Switch.scala 30:36:@10676.4]
  wire  _T_30401; // @[Switch.scala 30:53:@10678.4]
  wire  valid_33_14; // @[Switch.scala 30:36:@10679.4]
  wire  _T_30404; // @[Switch.scala 30:53:@10681.4]
  wire  valid_33_15; // @[Switch.scala 30:36:@10682.4]
  wire  _T_30407; // @[Switch.scala 30:53:@10684.4]
  wire  valid_33_16; // @[Switch.scala 30:36:@10685.4]
  wire  _T_30410; // @[Switch.scala 30:53:@10687.4]
  wire  valid_33_17; // @[Switch.scala 30:36:@10688.4]
  wire  _T_30413; // @[Switch.scala 30:53:@10690.4]
  wire  valid_33_18; // @[Switch.scala 30:36:@10691.4]
  wire  _T_30416; // @[Switch.scala 30:53:@10693.4]
  wire  valid_33_19; // @[Switch.scala 30:36:@10694.4]
  wire  _T_30419; // @[Switch.scala 30:53:@10696.4]
  wire  valid_33_20; // @[Switch.scala 30:36:@10697.4]
  wire  _T_30422; // @[Switch.scala 30:53:@10699.4]
  wire  valid_33_21; // @[Switch.scala 30:36:@10700.4]
  wire  _T_30425; // @[Switch.scala 30:53:@10702.4]
  wire  valid_33_22; // @[Switch.scala 30:36:@10703.4]
  wire  _T_30428; // @[Switch.scala 30:53:@10705.4]
  wire  valid_33_23; // @[Switch.scala 30:36:@10706.4]
  wire  _T_30431; // @[Switch.scala 30:53:@10708.4]
  wire  valid_33_24; // @[Switch.scala 30:36:@10709.4]
  wire  _T_30434; // @[Switch.scala 30:53:@10711.4]
  wire  valid_33_25; // @[Switch.scala 30:36:@10712.4]
  wire  _T_30437; // @[Switch.scala 30:53:@10714.4]
  wire  valid_33_26; // @[Switch.scala 30:36:@10715.4]
  wire  _T_30440; // @[Switch.scala 30:53:@10717.4]
  wire  valid_33_27; // @[Switch.scala 30:36:@10718.4]
  wire  _T_30443; // @[Switch.scala 30:53:@10720.4]
  wire  valid_33_28; // @[Switch.scala 30:36:@10721.4]
  wire  _T_30446; // @[Switch.scala 30:53:@10723.4]
  wire  valid_33_29; // @[Switch.scala 30:36:@10724.4]
  wire  _T_30449; // @[Switch.scala 30:53:@10726.4]
  wire  valid_33_30; // @[Switch.scala 30:36:@10727.4]
  wire  _T_30452; // @[Switch.scala 30:53:@10729.4]
  wire  valid_33_31; // @[Switch.scala 30:36:@10730.4]
  wire  _T_30455; // @[Switch.scala 30:53:@10732.4]
  wire  valid_33_32; // @[Switch.scala 30:36:@10733.4]
  wire  _T_30458; // @[Switch.scala 30:53:@10735.4]
  wire  valid_33_33; // @[Switch.scala 30:36:@10736.4]
  wire  _T_30461; // @[Switch.scala 30:53:@10738.4]
  wire  valid_33_34; // @[Switch.scala 30:36:@10739.4]
  wire  _T_30464; // @[Switch.scala 30:53:@10741.4]
  wire  valid_33_35; // @[Switch.scala 30:36:@10742.4]
  wire  _T_30467; // @[Switch.scala 30:53:@10744.4]
  wire  valid_33_36; // @[Switch.scala 30:36:@10745.4]
  wire  _T_30470; // @[Switch.scala 30:53:@10747.4]
  wire  valid_33_37; // @[Switch.scala 30:36:@10748.4]
  wire  _T_30473; // @[Switch.scala 30:53:@10750.4]
  wire  valid_33_38; // @[Switch.scala 30:36:@10751.4]
  wire  _T_30476; // @[Switch.scala 30:53:@10753.4]
  wire  valid_33_39; // @[Switch.scala 30:36:@10754.4]
  wire  _T_30479; // @[Switch.scala 30:53:@10756.4]
  wire  valid_33_40; // @[Switch.scala 30:36:@10757.4]
  wire  _T_30482; // @[Switch.scala 30:53:@10759.4]
  wire  valid_33_41; // @[Switch.scala 30:36:@10760.4]
  wire  _T_30485; // @[Switch.scala 30:53:@10762.4]
  wire  valid_33_42; // @[Switch.scala 30:36:@10763.4]
  wire  _T_30488; // @[Switch.scala 30:53:@10765.4]
  wire  valid_33_43; // @[Switch.scala 30:36:@10766.4]
  wire  _T_30491; // @[Switch.scala 30:53:@10768.4]
  wire  valid_33_44; // @[Switch.scala 30:36:@10769.4]
  wire  _T_30494; // @[Switch.scala 30:53:@10771.4]
  wire  valid_33_45; // @[Switch.scala 30:36:@10772.4]
  wire  _T_30497; // @[Switch.scala 30:53:@10774.4]
  wire  valid_33_46; // @[Switch.scala 30:36:@10775.4]
  wire  _T_30500; // @[Switch.scala 30:53:@10777.4]
  wire  valid_33_47; // @[Switch.scala 30:36:@10778.4]
  wire  _T_30503; // @[Switch.scala 30:53:@10780.4]
  wire  valid_33_48; // @[Switch.scala 30:36:@10781.4]
  wire  _T_30506; // @[Switch.scala 30:53:@10783.4]
  wire  valid_33_49; // @[Switch.scala 30:36:@10784.4]
  wire  _T_30509; // @[Switch.scala 30:53:@10786.4]
  wire  valid_33_50; // @[Switch.scala 30:36:@10787.4]
  wire  _T_30512; // @[Switch.scala 30:53:@10789.4]
  wire  valid_33_51; // @[Switch.scala 30:36:@10790.4]
  wire  _T_30515; // @[Switch.scala 30:53:@10792.4]
  wire  valid_33_52; // @[Switch.scala 30:36:@10793.4]
  wire  _T_30518; // @[Switch.scala 30:53:@10795.4]
  wire  valid_33_53; // @[Switch.scala 30:36:@10796.4]
  wire  _T_30521; // @[Switch.scala 30:53:@10798.4]
  wire  valid_33_54; // @[Switch.scala 30:36:@10799.4]
  wire  _T_30524; // @[Switch.scala 30:53:@10801.4]
  wire  valid_33_55; // @[Switch.scala 30:36:@10802.4]
  wire  _T_30527; // @[Switch.scala 30:53:@10804.4]
  wire  valid_33_56; // @[Switch.scala 30:36:@10805.4]
  wire  _T_30530; // @[Switch.scala 30:53:@10807.4]
  wire  valid_33_57; // @[Switch.scala 30:36:@10808.4]
  wire  _T_30533; // @[Switch.scala 30:53:@10810.4]
  wire  valid_33_58; // @[Switch.scala 30:36:@10811.4]
  wire  _T_30536; // @[Switch.scala 30:53:@10813.4]
  wire  valid_33_59; // @[Switch.scala 30:36:@10814.4]
  wire  _T_30539; // @[Switch.scala 30:53:@10816.4]
  wire  valid_33_60; // @[Switch.scala 30:36:@10817.4]
  wire  _T_30542; // @[Switch.scala 30:53:@10819.4]
  wire  valid_33_61; // @[Switch.scala 30:36:@10820.4]
  wire  _T_30545; // @[Switch.scala 30:53:@10822.4]
  wire  valid_33_62; // @[Switch.scala 30:36:@10823.4]
  wire  _T_30548; // @[Switch.scala 30:53:@10825.4]
  wire  valid_33_63; // @[Switch.scala 30:36:@10826.4]
  wire [5:0] _T_30614; // @[Mux.scala 31:69:@10828.4]
  wire [5:0] _T_30615; // @[Mux.scala 31:69:@10829.4]
  wire [5:0] _T_30616; // @[Mux.scala 31:69:@10830.4]
  wire [5:0] _T_30617; // @[Mux.scala 31:69:@10831.4]
  wire [5:0] _T_30618; // @[Mux.scala 31:69:@10832.4]
  wire [5:0] _T_30619; // @[Mux.scala 31:69:@10833.4]
  wire [5:0] _T_30620; // @[Mux.scala 31:69:@10834.4]
  wire [5:0] _T_30621; // @[Mux.scala 31:69:@10835.4]
  wire [5:0] _T_30622; // @[Mux.scala 31:69:@10836.4]
  wire [5:0] _T_30623; // @[Mux.scala 31:69:@10837.4]
  wire [5:0] _T_30624; // @[Mux.scala 31:69:@10838.4]
  wire [5:0] _T_30625; // @[Mux.scala 31:69:@10839.4]
  wire [5:0] _T_30626; // @[Mux.scala 31:69:@10840.4]
  wire [5:0] _T_30627; // @[Mux.scala 31:69:@10841.4]
  wire [5:0] _T_30628; // @[Mux.scala 31:69:@10842.4]
  wire [5:0] _T_30629; // @[Mux.scala 31:69:@10843.4]
  wire [5:0] _T_30630; // @[Mux.scala 31:69:@10844.4]
  wire [5:0] _T_30631; // @[Mux.scala 31:69:@10845.4]
  wire [5:0] _T_30632; // @[Mux.scala 31:69:@10846.4]
  wire [5:0] _T_30633; // @[Mux.scala 31:69:@10847.4]
  wire [5:0] _T_30634; // @[Mux.scala 31:69:@10848.4]
  wire [5:0] _T_30635; // @[Mux.scala 31:69:@10849.4]
  wire [5:0] _T_30636; // @[Mux.scala 31:69:@10850.4]
  wire [5:0] _T_30637; // @[Mux.scala 31:69:@10851.4]
  wire [5:0] _T_30638; // @[Mux.scala 31:69:@10852.4]
  wire [5:0] _T_30639; // @[Mux.scala 31:69:@10853.4]
  wire [5:0] _T_30640; // @[Mux.scala 31:69:@10854.4]
  wire [5:0] _T_30641; // @[Mux.scala 31:69:@10855.4]
  wire [5:0] _T_30642; // @[Mux.scala 31:69:@10856.4]
  wire [5:0] _T_30643; // @[Mux.scala 31:69:@10857.4]
  wire [5:0] _T_30644; // @[Mux.scala 31:69:@10858.4]
  wire [5:0] _T_30645; // @[Mux.scala 31:69:@10859.4]
  wire [5:0] _T_30646; // @[Mux.scala 31:69:@10860.4]
  wire [5:0] _T_30647; // @[Mux.scala 31:69:@10861.4]
  wire [5:0] _T_30648; // @[Mux.scala 31:69:@10862.4]
  wire [5:0] _T_30649; // @[Mux.scala 31:69:@10863.4]
  wire [5:0] _T_30650; // @[Mux.scala 31:69:@10864.4]
  wire [5:0] _T_30651; // @[Mux.scala 31:69:@10865.4]
  wire [5:0] _T_30652; // @[Mux.scala 31:69:@10866.4]
  wire [5:0] _T_30653; // @[Mux.scala 31:69:@10867.4]
  wire [5:0] _T_30654; // @[Mux.scala 31:69:@10868.4]
  wire [5:0] _T_30655; // @[Mux.scala 31:69:@10869.4]
  wire [5:0] _T_30656; // @[Mux.scala 31:69:@10870.4]
  wire [5:0] _T_30657; // @[Mux.scala 31:69:@10871.4]
  wire [5:0] _T_30658; // @[Mux.scala 31:69:@10872.4]
  wire [5:0] _T_30659; // @[Mux.scala 31:69:@10873.4]
  wire [5:0] _T_30660; // @[Mux.scala 31:69:@10874.4]
  wire [5:0] _T_30661; // @[Mux.scala 31:69:@10875.4]
  wire [5:0] _T_30662; // @[Mux.scala 31:69:@10876.4]
  wire [5:0] _T_30663; // @[Mux.scala 31:69:@10877.4]
  wire [5:0] _T_30664; // @[Mux.scala 31:69:@10878.4]
  wire [5:0] _T_30665; // @[Mux.scala 31:69:@10879.4]
  wire [5:0] _T_30666; // @[Mux.scala 31:69:@10880.4]
  wire [5:0] _T_30667; // @[Mux.scala 31:69:@10881.4]
  wire [5:0] _T_30668; // @[Mux.scala 31:69:@10882.4]
  wire [5:0] _T_30669; // @[Mux.scala 31:69:@10883.4]
  wire [5:0] _T_30670; // @[Mux.scala 31:69:@10884.4]
  wire [5:0] _T_30671; // @[Mux.scala 31:69:@10885.4]
  wire [5:0] _T_30672; // @[Mux.scala 31:69:@10886.4]
  wire [5:0] _T_30673; // @[Mux.scala 31:69:@10887.4]
  wire [5:0] _T_30674; // @[Mux.scala 31:69:@10888.4]
  wire [5:0] _T_30675; // @[Mux.scala 31:69:@10889.4]
  wire [5:0] select_33; // @[Mux.scala 31:69:@10890.4]
  wire [47:0] _GEN_2113; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2114; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2115; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2116; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2117; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2118; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2119; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2120; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2121; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2122; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2123; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2124; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2125; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2126; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2127; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2128; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2129; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2130; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2131; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2132; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2133; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2134; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2135; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2136; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2137; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2138; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2139; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2140; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2141; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2142; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2143; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2144; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2145; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2146; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2147; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2148; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2149; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2150; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2151; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2152; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2153; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2154; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2155; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2156; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2157; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2158; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2159; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2160; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2161; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2162; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2163; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2164; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2165; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2166; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2167; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2168; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2169; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2170; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2171; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2172; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2173; // @[Switch.scala 33:19:@10892.4]
  wire [47:0] _GEN_2174; // @[Switch.scala 33:19:@10892.4]
  wire [7:0] _T_30684; // @[Switch.scala 34:32:@10899.4]
  wire [15:0] _T_30692; // @[Switch.scala 34:32:@10907.4]
  wire [7:0] _T_30699; // @[Switch.scala 34:32:@10914.4]
  wire [31:0] _T_30708; // @[Switch.scala 34:32:@10923.4]
  wire [7:0] _T_30715; // @[Switch.scala 34:32:@10930.4]
  wire [15:0] _T_30723; // @[Switch.scala 34:32:@10938.4]
  wire [7:0] _T_30730; // @[Switch.scala 34:32:@10945.4]
  wire [31:0] _T_30739; // @[Switch.scala 34:32:@10954.4]
  wire [63:0] _T_30740; // @[Switch.scala 34:32:@10955.4]
  wire  _T_30744; // @[Switch.scala 30:53:@10958.4]
  wire  valid_34_0; // @[Switch.scala 30:36:@10959.4]
  wire  _T_30747; // @[Switch.scala 30:53:@10961.4]
  wire  valid_34_1; // @[Switch.scala 30:36:@10962.4]
  wire  _T_30750; // @[Switch.scala 30:53:@10964.4]
  wire  valid_34_2; // @[Switch.scala 30:36:@10965.4]
  wire  _T_30753; // @[Switch.scala 30:53:@10967.4]
  wire  valid_34_3; // @[Switch.scala 30:36:@10968.4]
  wire  _T_30756; // @[Switch.scala 30:53:@10970.4]
  wire  valid_34_4; // @[Switch.scala 30:36:@10971.4]
  wire  _T_30759; // @[Switch.scala 30:53:@10973.4]
  wire  valid_34_5; // @[Switch.scala 30:36:@10974.4]
  wire  _T_30762; // @[Switch.scala 30:53:@10976.4]
  wire  valid_34_6; // @[Switch.scala 30:36:@10977.4]
  wire  _T_30765; // @[Switch.scala 30:53:@10979.4]
  wire  valid_34_7; // @[Switch.scala 30:36:@10980.4]
  wire  _T_30768; // @[Switch.scala 30:53:@10982.4]
  wire  valid_34_8; // @[Switch.scala 30:36:@10983.4]
  wire  _T_30771; // @[Switch.scala 30:53:@10985.4]
  wire  valid_34_9; // @[Switch.scala 30:36:@10986.4]
  wire  _T_30774; // @[Switch.scala 30:53:@10988.4]
  wire  valid_34_10; // @[Switch.scala 30:36:@10989.4]
  wire  _T_30777; // @[Switch.scala 30:53:@10991.4]
  wire  valid_34_11; // @[Switch.scala 30:36:@10992.4]
  wire  _T_30780; // @[Switch.scala 30:53:@10994.4]
  wire  valid_34_12; // @[Switch.scala 30:36:@10995.4]
  wire  _T_30783; // @[Switch.scala 30:53:@10997.4]
  wire  valid_34_13; // @[Switch.scala 30:36:@10998.4]
  wire  _T_30786; // @[Switch.scala 30:53:@11000.4]
  wire  valid_34_14; // @[Switch.scala 30:36:@11001.4]
  wire  _T_30789; // @[Switch.scala 30:53:@11003.4]
  wire  valid_34_15; // @[Switch.scala 30:36:@11004.4]
  wire  _T_30792; // @[Switch.scala 30:53:@11006.4]
  wire  valid_34_16; // @[Switch.scala 30:36:@11007.4]
  wire  _T_30795; // @[Switch.scala 30:53:@11009.4]
  wire  valid_34_17; // @[Switch.scala 30:36:@11010.4]
  wire  _T_30798; // @[Switch.scala 30:53:@11012.4]
  wire  valid_34_18; // @[Switch.scala 30:36:@11013.4]
  wire  _T_30801; // @[Switch.scala 30:53:@11015.4]
  wire  valid_34_19; // @[Switch.scala 30:36:@11016.4]
  wire  _T_30804; // @[Switch.scala 30:53:@11018.4]
  wire  valid_34_20; // @[Switch.scala 30:36:@11019.4]
  wire  _T_30807; // @[Switch.scala 30:53:@11021.4]
  wire  valid_34_21; // @[Switch.scala 30:36:@11022.4]
  wire  _T_30810; // @[Switch.scala 30:53:@11024.4]
  wire  valid_34_22; // @[Switch.scala 30:36:@11025.4]
  wire  _T_30813; // @[Switch.scala 30:53:@11027.4]
  wire  valid_34_23; // @[Switch.scala 30:36:@11028.4]
  wire  _T_30816; // @[Switch.scala 30:53:@11030.4]
  wire  valid_34_24; // @[Switch.scala 30:36:@11031.4]
  wire  _T_30819; // @[Switch.scala 30:53:@11033.4]
  wire  valid_34_25; // @[Switch.scala 30:36:@11034.4]
  wire  _T_30822; // @[Switch.scala 30:53:@11036.4]
  wire  valid_34_26; // @[Switch.scala 30:36:@11037.4]
  wire  _T_30825; // @[Switch.scala 30:53:@11039.4]
  wire  valid_34_27; // @[Switch.scala 30:36:@11040.4]
  wire  _T_30828; // @[Switch.scala 30:53:@11042.4]
  wire  valid_34_28; // @[Switch.scala 30:36:@11043.4]
  wire  _T_30831; // @[Switch.scala 30:53:@11045.4]
  wire  valid_34_29; // @[Switch.scala 30:36:@11046.4]
  wire  _T_30834; // @[Switch.scala 30:53:@11048.4]
  wire  valid_34_30; // @[Switch.scala 30:36:@11049.4]
  wire  _T_30837; // @[Switch.scala 30:53:@11051.4]
  wire  valid_34_31; // @[Switch.scala 30:36:@11052.4]
  wire  _T_30840; // @[Switch.scala 30:53:@11054.4]
  wire  valid_34_32; // @[Switch.scala 30:36:@11055.4]
  wire  _T_30843; // @[Switch.scala 30:53:@11057.4]
  wire  valid_34_33; // @[Switch.scala 30:36:@11058.4]
  wire  _T_30846; // @[Switch.scala 30:53:@11060.4]
  wire  valid_34_34; // @[Switch.scala 30:36:@11061.4]
  wire  _T_30849; // @[Switch.scala 30:53:@11063.4]
  wire  valid_34_35; // @[Switch.scala 30:36:@11064.4]
  wire  _T_30852; // @[Switch.scala 30:53:@11066.4]
  wire  valid_34_36; // @[Switch.scala 30:36:@11067.4]
  wire  _T_30855; // @[Switch.scala 30:53:@11069.4]
  wire  valid_34_37; // @[Switch.scala 30:36:@11070.4]
  wire  _T_30858; // @[Switch.scala 30:53:@11072.4]
  wire  valid_34_38; // @[Switch.scala 30:36:@11073.4]
  wire  _T_30861; // @[Switch.scala 30:53:@11075.4]
  wire  valid_34_39; // @[Switch.scala 30:36:@11076.4]
  wire  _T_30864; // @[Switch.scala 30:53:@11078.4]
  wire  valid_34_40; // @[Switch.scala 30:36:@11079.4]
  wire  _T_30867; // @[Switch.scala 30:53:@11081.4]
  wire  valid_34_41; // @[Switch.scala 30:36:@11082.4]
  wire  _T_30870; // @[Switch.scala 30:53:@11084.4]
  wire  valid_34_42; // @[Switch.scala 30:36:@11085.4]
  wire  _T_30873; // @[Switch.scala 30:53:@11087.4]
  wire  valid_34_43; // @[Switch.scala 30:36:@11088.4]
  wire  _T_30876; // @[Switch.scala 30:53:@11090.4]
  wire  valid_34_44; // @[Switch.scala 30:36:@11091.4]
  wire  _T_30879; // @[Switch.scala 30:53:@11093.4]
  wire  valid_34_45; // @[Switch.scala 30:36:@11094.4]
  wire  _T_30882; // @[Switch.scala 30:53:@11096.4]
  wire  valid_34_46; // @[Switch.scala 30:36:@11097.4]
  wire  _T_30885; // @[Switch.scala 30:53:@11099.4]
  wire  valid_34_47; // @[Switch.scala 30:36:@11100.4]
  wire  _T_30888; // @[Switch.scala 30:53:@11102.4]
  wire  valid_34_48; // @[Switch.scala 30:36:@11103.4]
  wire  _T_30891; // @[Switch.scala 30:53:@11105.4]
  wire  valid_34_49; // @[Switch.scala 30:36:@11106.4]
  wire  _T_30894; // @[Switch.scala 30:53:@11108.4]
  wire  valid_34_50; // @[Switch.scala 30:36:@11109.4]
  wire  _T_30897; // @[Switch.scala 30:53:@11111.4]
  wire  valid_34_51; // @[Switch.scala 30:36:@11112.4]
  wire  _T_30900; // @[Switch.scala 30:53:@11114.4]
  wire  valid_34_52; // @[Switch.scala 30:36:@11115.4]
  wire  _T_30903; // @[Switch.scala 30:53:@11117.4]
  wire  valid_34_53; // @[Switch.scala 30:36:@11118.4]
  wire  _T_30906; // @[Switch.scala 30:53:@11120.4]
  wire  valid_34_54; // @[Switch.scala 30:36:@11121.4]
  wire  _T_30909; // @[Switch.scala 30:53:@11123.4]
  wire  valid_34_55; // @[Switch.scala 30:36:@11124.4]
  wire  _T_30912; // @[Switch.scala 30:53:@11126.4]
  wire  valid_34_56; // @[Switch.scala 30:36:@11127.4]
  wire  _T_30915; // @[Switch.scala 30:53:@11129.4]
  wire  valid_34_57; // @[Switch.scala 30:36:@11130.4]
  wire  _T_30918; // @[Switch.scala 30:53:@11132.4]
  wire  valid_34_58; // @[Switch.scala 30:36:@11133.4]
  wire  _T_30921; // @[Switch.scala 30:53:@11135.4]
  wire  valid_34_59; // @[Switch.scala 30:36:@11136.4]
  wire  _T_30924; // @[Switch.scala 30:53:@11138.4]
  wire  valid_34_60; // @[Switch.scala 30:36:@11139.4]
  wire  _T_30927; // @[Switch.scala 30:53:@11141.4]
  wire  valid_34_61; // @[Switch.scala 30:36:@11142.4]
  wire  _T_30930; // @[Switch.scala 30:53:@11144.4]
  wire  valid_34_62; // @[Switch.scala 30:36:@11145.4]
  wire  _T_30933; // @[Switch.scala 30:53:@11147.4]
  wire  valid_34_63; // @[Switch.scala 30:36:@11148.4]
  wire [5:0] _T_30999; // @[Mux.scala 31:69:@11150.4]
  wire [5:0] _T_31000; // @[Mux.scala 31:69:@11151.4]
  wire [5:0] _T_31001; // @[Mux.scala 31:69:@11152.4]
  wire [5:0] _T_31002; // @[Mux.scala 31:69:@11153.4]
  wire [5:0] _T_31003; // @[Mux.scala 31:69:@11154.4]
  wire [5:0] _T_31004; // @[Mux.scala 31:69:@11155.4]
  wire [5:0] _T_31005; // @[Mux.scala 31:69:@11156.4]
  wire [5:0] _T_31006; // @[Mux.scala 31:69:@11157.4]
  wire [5:0] _T_31007; // @[Mux.scala 31:69:@11158.4]
  wire [5:0] _T_31008; // @[Mux.scala 31:69:@11159.4]
  wire [5:0] _T_31009; // @[Mux.scala 31:69:@11160.4]
  wire [5:0] _T_31010; // @[Mux.scala 31:69:@11161.4]
  wire [5:0] _T_31011; // @[Mux.scala 31:69:@11162.4]
  wire [5:0] _T_31012; // @[Mux.scala 31:69:@11163.4]
  wire [5:0] _T_31013; // @[Mux.scala 31:69:@11164.4]
  wire [5:0] _T_31014; // @[Mux.scala 31:69:@11165.4]
  wire [5:0] _T_31015; // @[Mux.scala 31:69:@11166.4]
  wire [5:0] _T_31016; // @[Mux.scala 31:69:@11167.4]
  wire [5:0] _T_31017; // @[Mux.scala 31:69:@11168.4]
  wire [5:0] _T_31018; // @[Mux.scala 31:69:@11169.4]
  wire [5:0] _T_31019; // @[Mux.scala 31:69:@11170.4]
  wire [5:0] _T_31020; // @[Mux.scala 31:69:@11171.4]
  wire [5:0] _T_31021; // @[Mux.scala 31:69:@11172.4]
  wire [5:0] _T_31022; // @[Mux.scala 31:69:@11173.4]
  wire [5:0] _T_31023; // @[Mux.scala 31:69:@11174.4]
  wire [5:0] _T_31024; // @[Mux.scala 31:69:@11175.4]
  wire [5:0] _T_31025; // @[Mux.scala 31:69:@11176.4]
  wire [5:0] _T_31026; // @[Mux.scala 31:69:@11177.4]
  wire [5:0] _T_31027; // @[Mux.scala 31:69:@11178.4]
  wire [5:0] _T_31028; // @[Mux.scala 31:69:@11179.4]
  wire [5:0] _T_31029; // @[Mux.scala 31:69:@11180.4]
  wire [5:0] _T_31030; // @[Mux.scala 31:69:@11181.4]
  wire [5:0] _T_31031; // @[Mux.scala 31:69:@11182.4]
  wire [5:0] _T_31032; // @[Mux.scala 31:69:@11183.4]
  wire [5:0] _T_31033; // @[Mux.scala 31:69:@11184.4]
  wire [5:0] _T_31034; // @[Mux.scala 31:69:@11185.4]
  wire [5:0] _T_31035; // @[Mux.scala 31:69:@11186.4]
  wire [5:0] _T_31036; // @[Mux.scala 31:69:@11187.4]
  wire [5:0] _T_31037; // @[Mux.scala 31:69:@11188.4]
  wire [5:0] _T_31038; // @[Mux.scala 31:69:@11189.4]
  wire [5:0] _T_31039; // @[Mux.scala 31:69:@11190.4]
  wire [5:0] _T_31040; // @[Mux.scala 31:69:@11191.4]
  wire [5:0] _T_31041; // @[Mux.scala 31:69:@11192.4]
  wire [5:0] _T_31042; // @[Mux.scala 31:69:@11193.4]
  wire [5:0] _T_31043; // @[Mux.scala 31:69:@11194.4]
  wire [5:0] _T_31044; // @[Mux.scala 31:69:@11195.4]
  wire [5:0] _T_31045; // @[Mux.scala 31:69:@11196.4]
  wire [5:0] _T_31046; // @[Mux.scala 31:69:@11197.4]
  wire [5:0] _T_31047; // @[Mux.scala 31:69:@11198.4]
  wire [5:0] _T_31048; // @[Mux.scala 31:69:@11199.4]
  wire [5:0] _T_31049; // @[Mux.scala 31:69:@11200.4]
  wire [5:0] _T_31050; // @[Mux.scala 31:69:@11201.4]
  wire [5:0] _T_31051; // @[Mux.scala 31:69:@11202.4]
  wire [5:0] _T_31052; // @[Mux.scala 31:69:@11203.4]
  wire [5:0] _T_31053; // @[Mux.scala 31:69:@11204.4]
  wire [5:0] _T_31054; // @[Mux.scala 31:69:@11205.4]
  wire [5:0] _T_31055; // @[Mux.scala 31:69:@11206.4]
  wire [5:0] _T_31056; // @[Mux.scala 31:69:@11207.4]
  wire [5:0] _T_31057; // @[Mux.scala 31:69:@11208.4]
  wire [5:0] _T_31058; // @[Mux.scala 31:69:@11209.4]
  wire [5:0] _T_31059; // @[Mux.scala 31:69:@11210.4]
  wire [5:0] _T_31060; // @[Mux.scala 31:69:@11211.4]
  wire [5:0] select_34; // @[Mux.scala 31:69:@11212.4]
  wire [47:0] _GEN_2177; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2178; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2179; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2180; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2181; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2182; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2183; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2184; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2185; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2186; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2187; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2188; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2189; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2190; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2191; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2192; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2193; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2194; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2195; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2196; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2197; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2198; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2199; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2200; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2201; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2202; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2203; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2204; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2205; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2206; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2207; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2208; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2209; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2210; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2211; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2212; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2213; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2214; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2215; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2216; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2217; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2218; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2219; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2220; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2221; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2222; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2223; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2224; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2225; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2226; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2227; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2228; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2229; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2230; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2231; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2232; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2233; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2234; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2235; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2236; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2237; // @[Switch.scala 33:19:@11214.4]
  wire [47:0] _GEN_2238; // @[Switch.scala 33:19:@11214.4]
  wire [7:0] _T_31069; // @[Switch.scala 34:32:@11221.4]
  wire [15:0] _T_31077; // @[Switch.scala 34:32:@11229.4]
  wire [7:0] _T_31084; // @[Switch.scala 34:32:@11236.4]
  wire [31:0] _T_31093; // @[Switch.scala 34:32:@11245.4]
  wire [7:0] _T_31100; // @[Switch.scala 34:32:@11252.4]
  wire [15:0] _T_31108; // @[Switch.scala 34:32:@11260.4]
  wire [7:0] _T_31115; // @[Switch.scala 34:32:@11267.4]
  wire [31:0] _T_31124; // @[Switch.scala 34:32:@11276.4]
  wire [63:0] _T_31125; // @[Switch.scala 34:32:@11277.4]
  wire  _T_31129; // @[Switch.scala 30:53:@11280.4]
  wire  valid_35_0; // @[Switch.scala 30:36:@11281.4]
  wire  _T_31132; // @[Switch.scala 30:53:@11283.4]
  wire  valid_35_1; // @[Switch.scala 30:36:@11284.4]
  wire  _T_31135; // @[Switch.scala 30:53:@11286.4]
  wire  valid_35_2; // @[Switch.scala 30:36:@11287.4]
  wire  _T_31138; // @[Switch.scala 30:53:@11289.4]
  wire  valid_35_3; // @[Switch.scala 30:36:@11290.4]
  wire  _T_31141; // @[Switch.scala 30:53:@11292.4]
  wire  valid_35_4; // @[Switch.scala 30:36:@11293.4]
  wire  _T_31144; // @[Switch.scala 30:53:@11295.4]
  wire  valid_35_5; // @[Switch.scala 30:36:@11296.4]
  wire  _T_31147; // @[Switch.scala 30:53:@11298.4]
  wire  valid_35_6; // @[Switch.scala 30:36:@11299.4]
  wire  _T_31150; // @[Switch.scala 30:53:@11301.4]
  wire  valid_35_7; // @[Switch.scala 30:36:@11302.4]
  wire  _T_31153; // @[Switch.scala 30:53:@11304.4]
  wire  valid_35_8; // @[Switch.scala 30:36:@11305.4]
  wire  _T_31156; // @[Switch.scala 30:53:@11307.4]
  wire  valid_35_9; // @[Switch.scala 30:36:@11308.4]
  wire  _T_31159; // @[Switch.scala 30:53:@11310.4]
  wire  valid_35_10; // @[Switch.scala 30:36:@11311.4]
  wire  _T_31162; // @[Switch.scala 30:53:@11313.4]
  wire  valid_35_11; // @[Switch.scala 30:36:@11314.4]
  wire  _T_31165; // @[Switch.scala 30:53:@11316.4]
  wire  valid_35_12; // @[Switch.scala 30:36:@11317.4]
  wire  _T_31168; // @[Switch.scala 30:53:@11319.4]
  wire  valid_35_13; // @[Switch.scala 30:36:@11320.4]
  wire  _T_31171; // @[Switch.scala 30:53:@11322.4]
  wire  valid_35_14; // @[Switch.scala 30:36:@11323.4]
  wire  _T_31174; // @[Switch.scala 30:53:@11325.4]
  wire  valid_35_15; // @[Switch.scala 30:36:@11326.4]
  wire  _T_31177; // @[Switch.scala 30:53:@11328.4]
  wire  valid_35_16; // @[Switch.scala 30:36:@11329.4]
  wire  _T_31180; // @[Switch.scala 30:53:@11331.4]
  wire  valid_35_17; // @[Switch.scala 30:36:@11332.4]
  wire  _T_31183; // @[Switch.scala 30:53:@11334.4]
  wire  valid_35_18; // @[Switch.scala 30:36:@11335.4]
  wire  _T_31186; // @[Switch.scala 30:53:@11337.4]
  wire  valid_35_19; // @[Switch.scala 30:36:@11338.4]
  wire  _T_31189; // @[Switch.scala 30:53:@11340.4]
  wire  valid_35_20; // @[Switch.scala 30:36:@11341.4]
  wire  _T_31192; // @[Switch.scala 30:53:@11343.4]
  wire  valid_35_21; // @[Switch.scala 30:36:@11344.4]
  wire  _T_31195; // @[Switch.scala 30:53:@11346.4]
  wire  valid_35_22; // @[Switch.scala 30:36:@11347.4]
  wire  _T_31198; // @[Switch.scala 30:53:@11349.4]
  wire  valid_35_23; // @[Switch.scala 30:36:@11350.4]
  wire  _T_31201; // @[Switch.scala 30:53:@11352.4]
  wire  valid_35_24; // @[Switch.scala 30:36:@11353.4]
  wire  _T_31204; // @[Switch.scala 30:53:@11355.4]
  wire  valid_35_25; // @[Switch.scala 30:36:@11356.4]
  wire  _T_31207; // @[Switch.scala 30:53:@11358.4]
  wire  valid_35_26; // @[Switch.scala 30:36:@11359.4]
  wire  _T_31210; // @[Switch.scala 30:53:@11361.4]
  wire  valid_35_27; // @[Switch.scala 30:36:@11362.4]
  wire  _T_31213; // @[Switch.scala 30:53:@11364.4]
  wire  valid_35_28; // @[Switch.scala 30:36:@11365.4]
  wire  _T_31216; // @[Switch.scala 30:53:@11367.4]
  wire  valid_35_29; // @[Switch.scala 30:36:@11368.4]
  wire  _T_31219; // @[Switch.scala 30:53:@11370.4]
  wire  valid_35_30; // @[Switch.scala 30:36:@11371.4]
  wire  _T_31222; // @[Switch.scala 30:53:@11373.4]
  wire  valid_35_31; // @[Switch.scala 30:36:@11374.4]
  wire  _T_31225; // @[Switch.scala 30:53:@11376.4]
  wire  valid_35_32; // @[Switch.scala 30:36:@11377.4]
  wire  _T_31228; // @[Switch.scala 30:53:@11379.4]
  wire  valid_35_33; // @[Switch.scala 30:36:@11380.4]
  wire  _T_31231; // @[Switch.scala 30:53:@11382.4]
  wire  valid_35_34; // @[Switch.scala 30:36:@11383.4]
  wire  _T_31234; // @[Switch.scala 30:53:@11385.4]
  wire  valid_35_35; // @[Switch.scala 30:36:@11386.4]
  wire  _T_31237; // @[Switch.scala 30:53:@11388.4]
  wire  valid_35_36; // @[Switch.scala 30:36:@11389.4]
  wire  _T_31240; // @[Switch.scala 30:53:@11391.4]
  wire  valid_35_37; // @[Switch.scala 30:36:@11392.4]
  wire  _T_31243; // @[Switch.scala 30:53:@11394.4]
  wire  valid_35_38; // @[Switch.scala 30:36:@11395.4]
  wire  _T_31246; // @[Switch.scala 30:53:@11397.4]
  wire  valid_35_39; // @[Switch.scala 30:36:@11398.4]
  wire  _T_31249; // @[Switch.scala 30:53:@11400.4]
  wire  valid_35_40; // @[Switch.scala 30:36:@11401.4]
  wire  _T_31252; // @[Switch.scala 30:53:@11403.4]
  wire  valid_35_41; // @[Switch.scala 30:36:@11404.4]
  wire  _T_31255; // @[Switch.scala 30:53:@11406.4]
  wire  valid_35_42; // @[Switch.scala 30:36:@11407.4]
  wire  _T_31258; // @[Switch.scala 30:53:@11409.4]
  wire  valid_35_43; // @[Switch.scala 30:36:@11410.4]
  wire  _T_31261; // @[Switch.scala 30:53:@11412.4]
  wire  valid_35_44; // @[Switch.scala 30:36:@11413.4]
  wire  _T_31264; // @[Switch.scala 30:53:@11415.4]
  wire  valid_35_45; // @[Switch.scala 30:36:@11416.4]
  wire  _T_31267; // @[Switch.scala 30:53:@11418.4]
  wire  valid_35_46; // @[Switch.scala 30:36:@11419.4]
  wire  _T_31270; // @[Switch.scala 30:53:@11421.4]
  wire  valid_35_47; // @[Switch.scala 30:36:@11422.4]
  wire  _T_31273; // @[Switch.scala 30:53:@11424.4]
  wire  valid_35_48; // @[Switch.scala 30:36:@11425.4]
  wire  _T_31276; // @[Switch.scala 30:53:@11427.4]
  wire  valid_35_49; // @[Switch.scala 30:36:@11428.4]
  wire  _T_31279; // @[Switch.scala 30:53:@11430.4]
  wire  valid_35_50; // @[Switch.scala 30:36:@11431.4]
  wire  _T_31282; // @[Switch.scala 30:53:@11433.4]
  wire  valid_35_51; // @[Switch.scala 30:36:@11434.4]
  wire  _T_31285; // @[Switch.scala 30:53:@11436.4]
  wire  valid_35_52; // @[Switch.scala 30:36:@11437.4]
  wire  _T_31288; // @[Switch.scala 30:53:@11439.4]
  wire  valid_35_53; // @[Switch.scala 30:36:@11440.4]
  wire  _T_31291; // @[Switch.scala 30:53:@11442.4]
  wire  valid_35_54; // @[Switch.scala 30:36:@11443.4]
  wire  _T_31294; // @[Switch.scala 30:53:@11445.4]
  wire  valid_35_55; // @[Switch.scala 30:36:@11446.4]
  wire  _T_31297; // @[Switch.scala 30:53:@11448.4]
  wire  valid_35_56; // @[Switch.scala 30:36:@11449.4]
  wire  _T_31300; // @[Switch.scala 30:53:@11451.4]
  wire  valid_35_57; // @[Switch.scala 30:36:@11452.4]
  wire  _T_31303; // @[Switch.scala 30:53:@11454.4]
  wire  valid_35_58; // @[Switch.scala 30:36:@11455.4]
  wire  _T_31306; // @[Switch.scala 30:53:@11457.4]
  wire  valid_35_59; // @[Switch.scala 30:36:@11458.4]
  wire  _T_31309; // @[Switch.scala 30:53:@11460.4]
  wire  valid_35_60; // @[Switch.scala 30:36:@11461.4]
  wire  _T_31312; // @[Switch.scala 30:53:@11463.4]
  wire  valid_35_61; // @[Switch.scala 30:36:@11464.4]
  wire  _T_31315; // @[Switch.scala 30:53:@11466.4]
  wire  valid_35_62; // @[Switch.scala 30:36:@11467.4]
  wire  _T_31318; // @[Switch.scala 30:53:@11469.4]
  wire  valid_35_63; // @[Switch.scala 30:36:@11470.4]
  wire [5:0] _T_31384; // @[Mux.scala 31:69:@11472.4]
  wire [5:0] _T_31385; // @[Mux.scala 31:69:@11473.4]
  wire [5:0] _T_31386; // @[Mux.scala 31:69:@11474.4]
  wire [5:0] _T_31387; // @[Mux.scala 31:69:@11475.4]
  wire [5:0] _T_31388; // @[Mux.scala 31:69:@11476.4]
  wire [5:0] _T_31389; // @[Mux.scala 31:69:@11477.4]
  wire [5:0] _T_31390; // @[Mux.scala 31:69:@11478.4]
  wire [5:0] _T_31391; // @[Mux.scala 31:69:@11479.4]
  wire [5:0] _T_31392; // @[Mux.scala 31:69:@11480.4]
  wire [5:0] _T_31393; // @[Mux.scala 31:69:@11481.4]
  wire [5:0] _T_31394; // @[Mux.scala 31:69:@11482.4]
  wire [5:0] _T_31395; // @[Mux.scala 31:69:@11483.4]
  wire [5:0] _T_31396; // @[Mux.scala 31:69:@11484.4]
  wire [5:0] _T_31397; // @[Mux.scala 31:69:@11485.4]
  wire [5:0] _T_31398; // @[Mux.scala 31:69:@11486.4]
  wire [5:0] _T_31399; // @[Mux.scala 31:69:@11487.4]
  wire [5:0] _T_31400; // @[Mux.scala 31:69:@11488.4]
  wire [5:0] _T_31401; // @[Mux.scala 31:69:@11489.4]
  wire [5:0] _T_31402; // @[Mux.scala 31:69:@11490.4]
  wire [5:0] _T_31403; // @[Mux.scala 31:69:@11491.4]
  wire [5:0] _T_31404; // @[Mux.scala 31:69:@11492.4]
  wire [5:0] _T_31405; // @[Mux.scala 31:69:@11493.4]
  wire [5:0] _T_31406; // @[Mux.scala 31:69:@11494.4]
  wire [5:0] _T_31407; // @[Mux.scala 31:69:@11495.4]
  wire [5:0] _T_31408; // @[Mux.scala 31:69:@11496.4]
  wire [5:0] _T_31409; // @[Mux.scala 31:69:@11497.4]
  wire [5:0] _T_31410; // @[Mux.scala 31:69:@11498.4]
  wire [5:0] _T_31411; // @[Mux.scala 31:69:@11499.4]
  wire [5:0] _T_31412; // @[Mux.scala 31:69:@11500.4]
  wire [5:0] _T_31413; // @[Mux.scala 31:69:@11501.4]
  wire [5:0] _T_31414; // @[Mux.scala 31:69:@11502.4]
  wire [5:0] _T_31415; // @[Mux.scala 31:69:@11503.4]
  wire [5:0] _T_31416; // @[Mux.scala 31:69:@11504.4]
  wire [5:0] _T_31417; // @[Mux.scala 31:69:@11505.4]
  wire [5:0] _T_31418; // @[Mux.scala 31:69:@11506.4]
  wire [5:0] _T_31419; // @[Mux.scala 31:69:@11507.4]
  wire [5:0] _T_31420; // @[Mux.scala 31:69:@11508.4]
  wire [5:0] _T_31421; // @[Mux.scala 31:69:@11509.4]
  wire [5:0] _T_31422; // @[Mux.scala 31:69:@11510.4]
  wire [5:0] _T_31423; // @[Mux.scala 31:69:@11511.4]
  wire [5:0] _T_31424; // @[Mux.scala 31:69:@11512.4]
  wire [5:0] _T_31425; // @[Mux.scala 31:69:@11513.4]
  wire [5:0] _T_31426; // @[Mux.scala 31:69:@11514.4]
  wire [5:0] _T_31427; // @[Mux.scala 31:69:@11515.4]
  wire [5:0] _T_31428; // @[Mux.scala 31:69:@11516.4]
  wire [5:0] _T_31429; // @[Mux.scala 31:69:@11517.4]
  wire [5:0] _T_31430; // @[Mux.scala 31:69:@11518.4]
  wire [5:0] _T_31431; // @[Mux.scala 31:69:@11519.4]
  wire [5:0] _T_31432; // @[Mux.scala 31:69:@11520.4]
  wire [5:0] _T_31433; // @[Mux.scala 31:69:@11521.4]
  wire [5:0] _T_31434; // @[Mux.scala 31:69:@11522.4]
  wire [5:0] _T_31435; // @[Mux.scala 31:69:@11523.4]
  wire [5:0] _T_31436; // @[Mux.scala 31:69:@11524.4]
  wire [5:0] _T_31437; // @[Mux.scala 31:69:@11525.4]
  wire [5:0] _T_31438; // @[Mux.scala 31:69:@11526.4]
  wire [5:0] _T_31439; // @[Mux.scala 31:69:@11527.4]
  wire [5:0] _T_31440; // @[Mux.scala 31:69:@11528.4]
  wire [5:0] _T_31441; // @[Mux.scala 31:69:@11529.4]
  wire [5:0] _T_31442; // @[Mux.scala 31:69:@11530.4]
  wire [5:0] _T_31443; // @[Mux.scala 31:69:@11531.4]
  wire [5:0] _T_31444; // @[Mux.scala 31:69:@11532.4]
  wire [5:0] _T_31445; // @[Mux.scala 31:69:@11533.4]
  wire [5:0] select_35; // @[Mux.scala 31:69:@11534.4]
  wire [47:0] _GEN_2241; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2242; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2243; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2244; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2245; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2246; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2247; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2248; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2249; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2250; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2251; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2252; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2253; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2254; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2255; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2256; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2257; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2258; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2259; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2260; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2261; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2262; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2263; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2264; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2265; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2266; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2267; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2268; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2269; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2270; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2271; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2272; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2273; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2274; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2275; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2276; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2277; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2278; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2279; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2280; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2281; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2282; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2283; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2284; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2285; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2286; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2287; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2288; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2289; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2290; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2291; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2292; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2293; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2294; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2295; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2296; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2297; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2298; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2299; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2300; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2301; // @[Switch.scala 33:19:@11536.4]
  wire [47:0] _GEN_2302; // @[Switch.scala 33:19:@11536.4]
  wire [7:0] _T_31454; // @[Switch.scala 34:32:@11543.4]
  wire [15:0] _T_31462; // @[Switch.scala 34:32:@11551.4]
  wire [7:0] _T_31469; // @[Switch.scala 34:32:@11558.4]
  wire [31:0] _T_31478; // @[Switch.scala 34:32:@11567.4]
  wire [7:0] _T_31485; // @[Switch.scala 34:32:@11574.4]
  wire [15:0] _T_31493; // @[Switch.scala 34:32:@11582.4]
  wire [7:0] _T_31500; // @[Switch.scala 34:32:@11589.4]
  wire [31:0] _T_31509; // @[Switch.scala 34:32:@11598.4]
  wire [63:0] _T_31510; // @[Switch.scala 34:32:@11599.4]
  wire  _T_31514; // @[Switch.scala 30:53:@11602.4]
  wire  valid_36_0; // @[Switch.scala 30:36:@11603.4]
  wire  _T_31517; // @[Switch.scala 30:53:@11605.4]
  wire  valid_36_1; // @[Switch.scala 30:36:@11606.4]
  wire  _T_31520; // @[Switch.scala 30:53:@11608.4]
  wire  valid_36_2; // @[Switch.scala 30:36:@11609.4]
  wire  _T_31523; // @[Switch.scala 30:53:@11611.4]
  wire  valid_36_3; // @[Switch.scala 30:36:@11612.4]
  wire  _T_31526; // @[Switch.scala 30:53:@11614.4]
  wire  valid_36_4; // @[Switch.scala 30:36:@11615.4]
  wire  _T_31529; // @[Switch.scala 30:53:@11617.4]
  wire  valid_36_5; // @[Switch.scala 30:36:@11618.4]
  wire  _T_31532; // @[Switch.scala 30:53:@11620.4]
  wire  valid_36_6; // @[Switch.scala 30:36:@11621.4]
  wire  _T_31535; // @[Switch.scala 30:53:@11623.4]
  wire  valid_36_7; // @[Switch.scala 30:36:@11624.4]
  wire  _T_31538; // @[Switch.scala 30:53:@11626.4]
  wire  valid_36_8; // @[Switch.scala 30:36:@11627.4]
  wire  _T_31541; // @[Switch.scala 30:53:@11629.4]
  wire  valid_36_9; // @[Switch.scala 30:36:@11630.4]
  wire  _T_31544; // @[Switch.scala 30:53:@11632.4]
  wire  valid_36_10; // @[Switch.scala 30:36:@11633.4]
  wire  _T_31547; // @[Switch.scala 30:53:@11635.4]
  wire  valid_36_11; // @[Switch.scala 30:36:@11636.4]
  wire  _T_31550; // @[Switch.scala 30:53:@11638.4]
  wire  valid_36_12; // @[Switch.scala 30:36:@11639.4]
  wire  _T_31553; // @[Switch.scala 30:53:@11641.4]
  wire  valid_36_13; // @[Switch.scala 30:36:@11642.4]
  wire  _T_31556; // @[Switch.scala 30:53:@11644.4]
  wire  valid_36_14; // @[Switch.scala 30:36:@11645.4]
  wire  _T_31559; // @[Switch.scala 30:53:@11647.4]
  wire  valid_36_15; // @[Switch.scala 30:36:@11648.4]
  wire  _T_31562; // @[Switch.scala 30:53:@11650.4]
  wire  valid_36_16; // @[Switch.scala 30:36:@11651.4]
  wire  _T_31565; // @[Switch.scala 30:53:@11653.4]
  wire  valid_36_17; // @[Switch.scala 30:36:@11654.4]
  wire  _T_31568; // @[Switch.scala 30:53:@11656.4]
  wire  valid_36_18; // @[Switch.scala 30:36:@11657.4]
  wire  _T_31571; // @[Switch.scala 30:53:@11659.4]
  wire  valid_36_19; // @[Switch.scala 30:36:@11660.4]
  wire  _T_31574; // @[Switch.scala 30:53:@11662.4]
  wire  valid_36_20; // @[Switch.scala 30:36:@11663.4]
  wire  _T_31577; // @[Switch.scala 30:53:@11665.4]
  wire  valid_36_21; // @[Switch.scala 30:36:@11666.4]
  wire  _T_31580; // @[Switch.scala 30:53:@11668.4]
  wire  valid_36_22; // @[Switch.scala 30:36:@11669.4]
  wire  _T_31583; // @[Switch.scala 30:53:@11671.4]
  wire  valid_36_23; // @[Switch.scala 30:36:@11672.4]
  wire  _T_31586; // @[Switch.scala 30:53:@11674.4]
  wire  valid_36_24; // @[Switch.scala 30:36:@11675.4]
  wire  _T_31589; // @[Switch.scala 30:53:@11677.4]
  wire  valid_36_25; // @[Switch.scala 30:36:@11678.4]
  wire  _T_31592; // @[Switch.scala 30:53:@11680.4]
  wire  valid_36_26; // @[Switch.scala 30:36:@11681.4]
  wire  _T_31595; // @[Switch.scala 30:53:@11683.4]
  wire  valid_36_27; // @[Switch.scala 30:36:@11684.4]
  wire  _T_31598; // @[Switch.scala 30:53:@11686.4]
  wire  valid_36_28; // @[Switch.scala 30:36:@11687.4]
  wire  _T_31601; // @[Switch.scala 30:53:@11689.4]
  wire  valid_36_29; // @[Switch.scala 30:36:@11690.4]
  wire  _T_31604; // @[Switch.scala 30:53:@11692.4]
  wire  valid_36_30; // @[Switch.scala 30:36:@11693.4]
  wire  _T_31607; // @[Switch.scala 30:53:@11695.4]
  wire  valid_36_31; // @[Switch.scala 30:36:@11696.4]
  wire  _T_31610; // @[Switch.scala 30:53:@11698.4]
  wire  valid_36_32; // @[Switch.scala 30:36:@11699.4]
  wire  _T_31613; // @[Switch.scala 30:53:@11701.4]
  wire  valid_36_33; // @[Switch.scala 30:36:@11702.4]
  wire  _T_31616; // @[Switch.scala 30:53:@11704.4]
  wire  valid_36_34; // @[Switch.scala 30:36:@11705.4]
  wire  _T_31619; // @[Switch.scala 30:53:@11707.4]
  wire  valid_36_35; // @[Switch.scala 30:36:@11708.4]
  wire  _T_31622; // @[Switch.scala 30:53:@11710.4]
  wire  valid_36_36; // @[Switch.scala 30:36:@11711.4]
  wire  _T_31625; // @[Switch.scala 30:53:@11713.4]
  wire  valid_36_37; // @[Switch.scala 30:36:@11714.4]
  wire  _T_31628; // @[Switch.scala 30:53:@11716.4]
  wire  valid_36_38; // @[Switch.scala 30:36:@11717.4]
  wire  _T_31631; // @[Switch.scala 30:53:@11719.4]
  wire  valid_36_39; // @[Switch.scala 30:36:@11720.4]
  wire  _T_31634; // @[Switch.scala 30:53:@11722.4]
  wire  valid_36_40; // @[Switch.scala 30:36:@11723.4]
  wire  _T_31637; // @[Switch.scala 30:53:@11725.4]
  wire  valid_36_41; // @[Switch.scala 30:36:@11726.4]
  wire  _T_31640; // @[Switch.scala 30:53:@11728.4]
  wire  valid_36_42; // @[Switch.scala 30:36:@11729.4]
  wire  _T_31643; // @[Switch.scala 30:53:@11731.4]
  wire  valid_36_43; // @[Switch.scala 30:36:@11732.4]
  wire  _T_31646; // @[Switch.scala 30:53:@11734.4]
  wire  valid_36_44; // @[Switch.scala 30:36:@11735.4]
  wire  _T_31649; // @[Switch.scala 30:53:@11737.4]
  wire  valid_36_45; // @[Switch.scala 30:36:@11738.4]
  wire  _T_31652; // @[Switch.scala 30:53:@11740.4]
  wire  valid_36_46; // @[Switch.scala 30:36:@11741.4]
  wire  _T_31655; // @[Switch.scala 30:53:@11743.4]
  wire  valid_36_47; // @[Switch.scala 30:36:@11744.4]
  wire  _T_31658; // @[Switch.scala 30:53:@11746.4]
  wire  valid_36_48; // @[Switch.scala 30:36:@11747.4]
  wire  _T_31661; // @[Switch.scala 30:53:@11749.4]
  wire  valid_36_49; // @[Switch.scala 30:36:@11750.4]
  wire  _T_31664; // @[Switch.scala 30:53:@11752.4]
  wire  valid_36_50; // @[Switch.scala 30:36:@11753.4]
  wire  _T_31667; // @[Switch.scala 30:53:@11755.4]
  wire  valid_36_51; // @[Switch.scala 30:36:@11756.4]
  wire  _T_31670; // @[Switch.scala 30:53:@11758.4]
  wire  valid_36_52; // @[Switch.scala 30:36:@11759.4]
  wire  _T_31673; // @[Switch.scala 30:53:@11761.4]
  wire  valid_36_53; // @[Switch.scala 30:36:@11762.4]
  wire  _T_31676; // @[Switch.scala 30:53:@11764.4]
  wire  valid_36_54; // @[Switch.scala 30:36:@11765.4]
  wire  _T_31679; // @[Switch.scala 30:53:@11767.4]
  wire  valid_36_55; // @[Switch.scala 30:36:@11768.4]
  wire  _T_31682; // @[Switch.scala 30:53:@11770.4]
  wire  valid_36_56; // @[Switch.scala 30:36:@11771.4]
  wire  _T_31685; // @[Switch.scala 30:53:@11773.4]
  wire  valid_36_57; // @[Switch.scala 30:36:@11774.4]
  wire  _T_31688; // @[Switch.scala 30:53:@11776.4]
  wire  valid_36_58; // @[Switch.scala 30:36:@11777.4]
  wire  _T_31691; // @[Switch.scala 30:53:@11779.4]
  wire  valid_36_59; // @[Switch.scala 30:36:@11780.4]
  wire  _T_31694; // @[Switch.scala 30:53:@11782.4]
  wire  valid_36_60; // @[Switch.scala 30:36:@11783.4]
  wire  _T_31697; // @[Switch.scala 30:53:@11785.4]
  wire  valid_36_61; // @[Switch.scala 30:36:@11786.4]
  wire  _T_31700; // @[Switch.scala 30:53:@11788.4]
  wire  valid_36_62; // @[Switch.scala 30:36:@11789.4]
  wire  _T_31703; // @[Switch.scala 30:53:@11791.4]
  wire  valid_36_63; // @[Switch.scala 30:36:@11792.4]
  wire [5:0] _T_31769; // @[Mux.scala 31:69:@11794.4]
  wire [5:0] _T_31770; // @[Mux.scala 31:69:@11795.4]
  wire [5:0] _T_31771; // @[Mux.scala 31:69:@11796.4]
  wire [5:0] _T_31772; // @[Mux.scala 31:69:@11797.4]
  wire [5:0] _T_31773; // @[Mux.scala 31:69:@11798.4]
  wire [5:0] _T_31774; // @[Mux.scala 31:69:@11799.4]
  wire [5:0] _T_31775; // @[Mux.scala 31:69:@11800.4]
  wire [5:0] _T_31776; // @[Mux.scala 31:69:@11801.4]
  wire [5:0] _T_31777; // @[Mux.scala 31:69:@11802.4]
  wire [5:0] _T_31778; // @[Mux.scala 31:69:@11803.4]
  wire [5:0] _T_31779; // @[Mux.scala 31:69:@11804.4]
  wire [5:0] _T_31780; // @[Mux.scala 31:69:@11805.4]
  wire [5:0] _T_31781; // @[Mux.scala 31:69:@11806.4]
  wire [5:0] _T_31782; // @[Mux.scala 31:69:@11807.4]
  wire [5:0] _T_31783; // @[Mux.scala 31:69:@11808.4]
  wire [5:0] _T_31784; // @[Mux.scala 31:69:@11809.4]
  wire [5:0] _T_31785; // @[Mux.scala 31:69:@11810.4]
  wire [5:0] _T_31786; // @[Mux.scala 31:69:@11811.4]
  wire [5:0] _T_31787; // @[Mux.scala 31:69:@11812.4]
  wire [5:0] _T_31788; // @[Mux.scala 31:69:@11813.4]
  wire [5:0] _T_31789; // @[Mux.scala 31:69:@11814.4]
  wire [5:0] _T_31790; // @[Mux.scala 31:69:@11815.4]
  wire [5:0] _T_31791; // @[Mux.scala 31:69:@11816.4]
  wire [5:0] _T_31792; // @[Mux.scala 31:69:@11817.4]
  wire [5:0] _T_31793; // @[Mux.scala 31:69:@11818.4]
  wire [5:0] _T_31794; // @[Mux.scala 31:69:@11819.4]
  wire [5:0] _T_31795; // @[Mux.scala 31:69:@11820.4]
  wire [5:0] _T_31796; // @[Mux.scala 31:69:@11821.4]
  wire [5:0] _T_31797; // @[Mux.scala 31:69:@11822.4]
  wire [5:0] _T_31798; // @[Mux.scala 31:69:@11823.4]
  wire [5:0] _T_31799; // @[Mux.scala 31:69:@11824.4]
  wire [5:0] _T_31800; // @[Mux.scala 31:69:@11825.4]
  wire [5:0] _T_31801; // @[Mux.scala 31:69:@11826.4]
  wire [5:0] _T_31802; // @[Mux.scala 31:69:@11827.4]
  wire [5:0] _T_31803; // @[Mux.scala 31:69:@11828.4]
  wire [5:0] _T_31804; // @[Mux.scala 31:69:@11829.4]
  wire [5:0] _T_31805; // @[Mux.scala 31:69:@11830.4]
  wire [5:0] _T_31806; // @[Mux.scala 31:69:@11831.4]
  wire [5:0] _T_31807; // @[Mux.scala 31:69:@11832.4]
  wire [5:0] _T_31808; // @[Mux.scala 31:69:@11833.4]
  wire [5:0] _T_31809; // @[Mux.scala 31:69:@11834.4]
  wire [5:0] _T_31810; // @[Mux.scala 31:69:@11835.4]
  wire [5:0] _T_31811; // @[Mux.scala 31:69:@11836.4]
  wire [5:0] _T_31812; // @[Mux.scala 31:69:@11837.4]
  wire [5:0] _T_31813; // @[Mux.scala 31:69:@11838.4]
  wire [5:0] _T_31814; // @[Mux.scala 31:69:@11839.4]
  wire [5:0] _T_31815; // @[Mux.scala 31:69:@11840.4]
  wire [5:0] _T_31816; // @[Mux.scala 31:69:@11841.4]
  wire [5:0] _T_31817; // @[Mux.scala 31:69:@11842.4]
  wire [5:0] _T_31818; // @[Mux.scala 31:69:@11843.4]
  wire [5:0] _T_31819; // @[Mux.scala 31:69:@11844.4]
  wire [5:0] _T_31820; // @[Mux.scala 31:69:@11845.4]
  wire [5:0] _T_31821; // @[Mux.scala 31:69:@11846.4]
  wire [5:0] _T_31822; // @[Mux.scala 31:69:@11847.4]
  wire [5:0] _T_31823; // @[Mux.scala 31:69:@11848.4]
  wire [5:0] _T_31824; // @[Mux.scala 31:69:@11849.4]
  wire [5:0] _T_31825; // @[Mux.scala 31:69:@11850.4]
  wire [5:0] _T_31826; // @[Mux.scala 31:69:@11851.4]
  wire [5:0] _T_31827; // @[Mux.scala 31:69:@11852.4]
  wire [5:0] _T_31828; // @[Mux.scala 31:69:@11853.4]
  wire [5:0] _T_31829; // @[Mux.scala 31:69:@11854.4]
  wire [5:0] _T_31830; // @[Mux.scala 31:69:@11855.4]
  wire [5:0] select_36; // @[Mux.scala 31:69:@11856.4]
  wire [47:0] _GEN_2305; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2306; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2307; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2308; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2309; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2310; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2311; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2312; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2313; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2314; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2315; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2316; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2317; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2318; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2319; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2320; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2321; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2322; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2323; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2324; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2325; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2326; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2327; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2328; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2329; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2330; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2331; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2332; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2333; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2334; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2335; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2336; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2337; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2338; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2339; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2340; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2341; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2342; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2343; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2344; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2345; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2346; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2347; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2348; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2349; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2350; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2351; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2352; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2353; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2354; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2355; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2356; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2357; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2358; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2359; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2360; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2361; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2362; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2363; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2364; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2365; // @[Switch.scala 33:19:@11858.4]
  wire [47:0] _GEN_2366; // @[Switch.scala 33:19:@11858.4]
  wire [7:0] _T_31839; // @[Switch.scala 34:32:@11865.4]
  wire [15:0] _T_31847; // @[Switch.scala 34:32:@11873.4]
  wire [7:0] _T_31854; // @[Switch.scala 34:32:@11880.4]
  wire [31:0] _T_31863; // @[Switch.scala 34:32:@11889.4]
  wire [7:0] _T_31870; // @[Switch.scala 34:32:@11896.4]
  wire [15:0] _T_31878; // @[Switch.scala 34:32:@11904.4]
  wire [7:0] _T_31885; // @[Switch.scala 34:32:@11911.4]
  wire [31:0] _T_31894; // @[Switch.scala 34:32:@11920.4]
  wire [63:0] _T_31895; // @[Switch.scala 34:32:@11921.4]
  wire  _T_31899; // @[Switch.scala 30:53:@11924.4]
  wire  valid_37_0; // @[Switch.scala 30:36:@11925.4]
  wire  _T_31902; // @[Switch.scala 30:53:@11927.4]
  wire  valid_37_1; // @[Switch.scala 30:36:@11928.4]
  wire  _T_31905; // @[Switch.scala 30:53:@11930.4]
  wire  valid_37_2; // @[Switch.scala 30:36:@11931.4]
  wire  _T_31908; // @[Switch.scala 30:53:@11933.4]
  wire  valid_37_3; // @[Switch.scala 30:36:@11934.4]
  wire  _T_31911; // @[Switch.scala 30:53:@11936.4]
  wire  valid_37_4; // @[Switch.scala 30:36:@11937.4]
  wire  _T_31914; // @[Switch.scala 30:53:@11939.4]
  wire  valid_37_5; // @[Switch.scala 30:36:@11940.4]
  wire  _T_31917; // @[Switch.scala 30:53:@11942.4]
  wire  valid_37_6; // @[Switch.scala 30:36:@11943.4]
  wire  _T_31920; // @[Switch.scala 30:53:@11945.4]
  wire  valid_37_7; // @[Switch.scala 30:36:@11946.4]
  wire  _T_31923; // @[Switch.scala 30:53:@11948.4]
  wire  valid_37_8; // @[Switch.scala 30:36:@11949.4]
  wire  _T_31926; // @[Switch.scala 30:53:@11951.4]
  wire  valid_37_9; // @[Switch.scala 30:36:@11952.4]
  wire  _T_31929; // @[Switch.scala 30:53:@11954.4]
  wire  valid_37_10; // @[Switch.scala 30:36:@11955.4]
  wire  _T_31932; // @[Switch.scala 30:53:@11957.4]
  wire  valid_37_11; // @[Switch.scala 30:36:@11958.4]
  wire  _T_31935; // @[Switch.scala 30:53:@11960.4]
  wire  valid_37_12; // @[Switch.scala 30:36:@11961.4]
  wire  _T_31938; // @[Switch.scala 30:53:@11963.4]
  wire  valid_37_13; // @[Switch.scala 30:36:@11964.4]
  wire  _T_31941; // @[Switch.scala 30:53:@11966.4]
  wire  valid_37_14; // @[Switch.scala 30:36:@11967.4]
  wire  _T_31944; // @[Switch.scala 30:53:@11969.4]
  wire  valid_37_15; // @[Switch.scala 30:36:@11970.4]
  wire  _T_31947; // @[Switch.scala 30:53:@11972.4]
  wire  valid_37_16; // @[Switch.scala 30:36:@11973.4]
  wire  _T_31950; // @[Switch.scala 30:53:@11975.4]
  wire  valid_37_17; // @[Switch.scala 30:36:@11976.4]
  wire  _T_31953; // @[Switch.scala 30:53:@11978.4]
  wire  valid_37_18; // @[Switch.scala 30:36:@11979.4]
  wire  _T_31956; // @[Switch.scala 30:53:@11981.4]
  wire  valid_37_19; // @[Switch.scala 30:36:@11982.4]
  wire  _T_31959; // @[Switch.scala 30:53:@11984.4]
  wire  valid_37_20; // @[Switch.scala 30:36:@11985.4]
  wire  _T_31962; // @[Switch.scala 30:53:@11987.4]
  wire  valid_37_21; // @[Switch.scala 30:36:@11988.4]
  wire  _T_31965; // @[Switch.scala 30:53:@11990.4]
  wire  valid_37_22; // @[Switch.scala 30:36:@11991.4]
  wire  _T_31968; // @[Switch.scala 30:53:@11993.4]
  wire  valid_37_23; // @[Switch.scala 30:36:@11994.4]
  wire  _T_31971; // @[Switch.scala 30:53:@11996.4]
  wire  valid_37_24; // @[Switch.scala 30:36:@11997.4]
  wire  _T_31974; // @[Switch.scala 30:53:@11999.4]
  wire  valid_37_25; // @[Switch.scala 30:36:@12000.4]
  wire  _T_31977; // @[Switch.scala 30:53:@12002.4]
  wire  valid_37_26; // @[Switch.scala 30:36:@12003.4]
  wire  _T_31980; // @[Switch.scala 30:53:@12005.4]
  wire  valid_37_27; // @[Switch.scala 30:36:@12006.4]
  wire  _T_31983; // @[Switch.scala 30:53:@12008.4]
  wire  valid_37_28; // @[Switch.scala 30:36:@12009.4]
  wire  _T_31986; // @[Switch.scala 30:53:@12011.4]
  wire  valid_37_29; // @[Switch.scala 30:36:@12012.4]
  wire  _T_31989; // @[Switch.scala 30:53:@12014.4]
  wire  valid_37_30; // @[Switch.scala 30:36:@12015.4]
  wire  _T_31992; // @[Switch.scala 30:53:@12017.4]
  wire  valid_37_31; // @[Switch.scala 30:36:@12018.4]
  wire  _T_31995; // @[Switch.scala 30:53:@12020.4]
  wire  valid_37_32; // @[Switch.scala 30:36:@12021.4]
  wire  _T_31998; // @[Switch.scala 30:53:@12023.4]
  wire  valid_37_33; // @[Switch.scala 30:36:@12024.4]
  wire  _T_32001; // @[Switch.scala 30:53:@12026.4]
  wire  valid_37_34; // @[Switch.scala 30:36:@12027.4]
  wire  _T_32004; // @[Switch.scala 30:53:@12029.4]
  wire  valid_37_35; // @[Switch.scala 30:36:@12030.4]
  wire  _T_32007; // @[Switch.scala 30:53:@12032.4]
  wire  valid_37_36; // @[Switch.scala 30:36:@12033.4]
  wire  _T_32010; // @[Switch.scala 30:53:@12035.4]
  wire  valid_37_37; // @[Switch.scala 30:36:@12036.4]
  wire  _T_32013; // @[Switch.scala 30:53:@12038.4]
  wire  valid_37_38; // @[Switch.scala 30:36:@12039.4]
  wire  _T_32016; // @[Switch.scala 30:53:@12041.4]
  wire  valid_37_39; // @[Switch.scala 30:36:@12042.4]
  wire  _T_32019; // @[Switch.scala 30:53:@12044.4]
  wire  valid_37_40; // @[Switch.scala 30:36:@12045.4]
  wire  _T_32022; // @[Switch.scala 30:53:@12047.4]
  wire  valid_37_41; // @[Switch.scala 30:36:@12048.4]
  wire  _T_32025; // @[Switch.scala 30:53:@12050.4]
  wire  valid_37_42; // @[Switch.scala 30:36:@12051.4]
  wire  _T_32028; // @[Switch.scala 30:53:@12053.4]
  wire  valid_37_43; // @[Switch.scala 30:36:@12054.4]
  wire  _T_32031; // @[Switch.scala 30:53:@12056.4]
  wire  valid_37_44; // @[Switch.scala 30:36:@12057.4]
  wire  _T_32034; // @[Switch.scala 30:53:@12059.4]
  wire  valid_37_45; // @[Switch.scala 30:36:@12060.4]
  wire  _T_32037; // @[Switch.scala 30:53:@12062.4]
  wire  valid_37_46; // @[Switch.scala 30:36:@12063.4]
  wire  _T_32040; // @[Switch.scala 30:53:@12065.4]
  wire  valid_37_47; // @[Switch.scala 30:36:@12066.4]
  wire  _T_32043; // @[Switch.scala 30:53:@12068.4]
  wire  valid_37_48; // @[Switch.scala 30:36:@12069.4]
  wire  _T_32046; // @[Switch.scala 30:53:@12071.4]
  wire  valid_37_49; // @[Switch.scala 30:36:@12072.4]
  wire  _T_32049; // @[Switch.scala 30:53:@12074.4]
  wire  valid_37_50; // @[Switch.scala 30:36:@12075.4]
  wire  _T_32052; // @[Switch.scala 30:53:@12077.4]
  wire  valid_37_51; // @[Switch.scala 30:36:@12078.4]
  wire  _T_32055; // @[Switch.scala 30:53:@12080.4]
  wire  valid_37_52; // @[Switch.scala 30:36:@12081.4]
  wire  _T_32058; // @[Switch.scala 30:53:@12083.4]
  wire  valid_37_53; // @[Switch.scala 30:36:@12084.4]
  wire  _T_32061; // @[Switch.scala 30:53:@12086.4]
  wire  valid_37_54; // @[Switch.scala 30:36:@12087.4]
  wire  _T_32064; // @[Switch.scala 30:53:@12089.4]
  wire  valid_37_55; // @[Switch.scala 30:36:@12090.4]
  wire  _T_32067; // @[Switch.scala 30:53:@12092.4]
  wire  valid_37_56; // @[Switch.scala 30:36:@12093.4]
  wire  _T_32070; // @[Switch.scala 30:53:@12095.4]
  wire  valid_37_57; // @[Switch.scala 30:36:@12096.4]
  wire  _T_32073; // @[Switch.scala 30:53:@12098.4]
  wire  valid_37_58; // @[Switch.scala 30:36:@12099.4]
  wire  _T_32076; // @[Switch.scala 30:53:@12101.4]
  wire  valid_37_59; // @[Switch.scala 30:36:@12102.4]
  wire  _T_32079; // @[Switch.scala 30:53:@12104.4]
  wire  valid_37_60; // @[Switch.scala 30:36:@12105.4]
  wire  _T_32082; // @[Switch.scala 30:53:@12107.4]
  wire  valid_37_61; // @[Switch.scala 30:36:@12108.4]
  wire  _T_32085; // @[Switch.scala 30:53:@12110.4]
  wire  valid_37_62; // @[Switch.scala 30:36:@12111.4]
  wire  _T_32088; // @[Switch.scala 30:53:@12113.4]
  wire  valid_37_63; // @[Switch.scala 30:36:@12114.4]
  wire [5:0] _T_32154; // @[Mux.scala 31:69:@12116.4]
  wire [5:0] _T_32155; // @[Mux.scala 31:69:@12117.4]
  wire [5:0] _T_32156; // @[Mux.scala 31:69:@12118.4]
  wire [5:0] _T_32157; // @[Mux.scala 31:69:@12119.4]
  wire [5:0] _T_32158; // @[Mux.scala 31:69:@12120.4]
  wire [5:0] _T_32159; // @[Mux.scala 31:69:@12121.4]
  wire [5:0] _T_32160; // @[Mux.scala 31:69:@12122.4]
  wire [5:0] _T_32161; // @[Mux.scala 31:69:@12123.4]
  wire [5:0] _T_32162; // @[Mux.scala 31:69:@12124.4]
  wire [5:0] _T_32163; // @[Mux.scala 31:69:@12125.4]
  wire [5:0] _T_32164; // @[Mux.scala 31:69:@12126.4]
  wire [5:0] _T_32165; // @[Mux.scala 31:69:@12127.4]
  wire [5:0] _T_32166; // @[Mux.scala 31:69:@12128.4]
  wire [5:0] _T_32167; // @[Mux.scala 31:69:@12129.4]
  wire [5:0] _T_32168; // @[Mux.scala 31:69:@12130.4]
  wire [5:0] _T_32169; // @[Mux.scala 31:69:@12131.4]
  wire [5:0] _T_32170; // @[Mux.scala 31:69:@12132.4]
  wire [5:0] _T_32171; // @[Mux.scala 31:69:@12133.4]
  wire [5:0] _T_32172; // @[Mux.scala 31:69:@12134.4]
  wire [5:0] _T_32173; // @[Mux.scala 31:69:@12135.4]
  wire [5:0] _T_32174; // @[Mux.scala 31:69:@12136.4]
  wire [5:0] _T_32175; // @[Mux.scala 31:69:@12137.4]
  wire [5:0] _T_32176; // @[Mux.scala 31:69:@12138.4]
  wire [5:0] _T_32177; // @[Mux.scala 31:69:@12139.4]
  wire [5:0] _T_32178; // @[Mux.scala 31:69:@12140.4]
  wire [5:0] _T_32179; // @[Mux.scala 31:69:@12141.4]
  wire [5:0] _T_32180; // @[Mux.scala 31:69:@12142.4]
  wire [5:0] _T_32181; // @[Mux.scala 31:69:@12143.4]
  wire [5:0] _T_32182; // @[Mux.scala 31:69:@12144.4]
  wire [5:0] _T_32183; // @[Mux.scala 31:69:@12145.4]
  wire [5:0] _T_32184; // @[Mux.scala 31:69:@12146.4]
  wire [5:0] _T_32185; // @[Mux.scala 31:69:@12147.4]
  wire [5:0] _T_32186; // @[Mux.scala 31:69:@12148.4]
  wire [5:0] _T_32187; // @[Mux.scala 31:69:@12149.4]
  wire [5:0] _T_32188; // @[Mux.scala 31:69:@12150.4]
  wire [5:0] _T_32189; // @[Mux.scala 31:69:@12151.4]
  wire [5:0] _T_32190; // @[Mux.scala 31:69:@12152.4]
  wire [5:0] _T_32191; // @[Mux.scala 31:69:@12153.4]
  wire [5:0] _T_32192; // @[Mux.scala 31:69:@12154.4]
  wire [5:0] _T_32193; // @[Mux.scala 31:69:@12155.4]
  wire [5:0] _T_32194; // @[Mux.scala 31:69:@12156.4]
  wire [5:0] _T_32195; // @[Mux.scala 31:69:@12157.4]
  wire [5:0] _T_32196; // @[Mux.scala 31:69:@12158.4]
  wire [5:0] _T_32197; // @[Mux.scala 31:69:@12159.4]
  wire [5:0] _T_32198; // @[Mux.scala 31:69:@12160.4]
  wire [5:0] _T_32199; // @[Mux.scala 31:69:@12161.4]
  wire [5:0] _T_32200; // @[Mux.scala 31:69:@12162.4]
  wire [5:0] _T_32201; // @[Mux.scala 31:69:@12163.4]
  wire [5:0] _T_32202; // @[Mux.scala 31:69:@12164.4]
  wire [5:0] _T_32203; // @[Mux.scala 31:69:@12165.4]
  wire [5:0] _T_32204; // @[Mux.scala 31:69:@12166.4]
  wire [5:0] _T_32205; // @[Mux.scala 31:69:@12167.4]
  wire [5:0] _T_32206; // @[Mux.scala 31:69:@12168.4]
  wire [5:0] _T_32207; // @[Mux.scala 31:69:@12169.4]
  wire [5:0] _T_32208; // @[Mux.scala 31:69:@12170.4]
  wire [5:0] _T_32209; // @[Mux.scala 31:69:@12171.4]
  wire [5:0] _T_32210; // @[Mux.scala 31:69:@12172.4]
  wire [5:0] _T_32211; // @[Mux.scala 31:69:@12173.4]
  wire [5:0] _T_32212; // @[Mux.scala 31:69:@12174.4]
  wire [5:0] _T_32213; // @[Mux.scala 31:69:@12175.4]
  wire [5:0] _T_32214; // @[Mux.scala 31:69:@12176.4]
  wire [5:0] _T_32215; // @[Mux.scala 31:69:@12177.4]
  wire [5:0] select_37; // @[Mux.scala 31:69:@12178.4]
  wire [47:0] _GEN_2369; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2370; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2371; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2372; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2373; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2374; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2375; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2376; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2377; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2378; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2379; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2380; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2381; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2382; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2383; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2384; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2385; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2386; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2387; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2388; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2389; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2390; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2391; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2392; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2393; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2394; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2395; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2396; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2397; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2398; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2399; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2400; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2401; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2402; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2403; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2404; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2405; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2406; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2407; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2408; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2409; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2410; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2411; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2412; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2413; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2414; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2415; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2416; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2417; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2418; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2419; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2420; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2421; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2422; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2423; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2424; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2425; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2426; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2427; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2428; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2429; // @[Switch.scala 33:19:@12180.4]
  wire [47:0] _GEN_2430; // @[Switch.scala 33:19:@12180.4]
  wire [7:0] _T_32224; // @[Switch.scala 34:32:@12187.4]
  wire [15:0] _T_32232; // @[Switch.scala 34:32:@12195.4]
  wire [7:0] _T_32239; // @[Switch.scala 34:32:@12202.4]
  wire [31:0] _T_32248; // @[Switch.scala 34:32:@12211.4]
  wire [7:0] _T_32255; // @[Switch.scala 34:32:@12218.4]
  wire [15:0] _T_32263; // @[Switch.scala 34:32:@12226.4]
  wire [7:0] _T_32270; // @[Switch.scala 34:32:@12233.4]
  wire [31:0] _T_32279; // @[Switch.scala 34:32:@12242.4]
  wire [63:0] _T_32280; // @[Switch.scala 34:32:@12243.4]
  wire  _T_32284; // @[Switch.scala 30:53:@12246.4]
  wire  valid_38_0; // @[Switch.scala 30:36:@12247.4]
  wire  _T_32287; // @[Switch.scala 30:53:@12249.4]
  wire  valid_38_1; // @[Switch.scala 30:36:@12250.4]
  wire  _T_32290; // @[Switch.scala 30:53:@12252.4]
  wire  valid_38_2; // @[Switch.scala 30:36:@12253.4]
  wire  _T_32293; // @[Switch.scala 30:53:@12255.4]
  wire  valid_38_3; // @[Switch.scala 30:36:@12256.4]
  wire  _T_32296; // @[Switch.scala 30:53:@12258.4]
  wire  valid_38_4; // @[Switch.scala 30:36:@12259.4]
  wire  _T_32299; // @[Switch.scala 30:53:@12261.4]
  wire  valid_38_5; // @[Switch.scala 30:36:@12262.4]
  wire  _T_32302; // @[Switch.scala 30:53:@12264.4]
  wire  valid_38_6; // @[Switch.scala 30:36:@12265.4]
  wire  _T_32305; // @[Switch.scala 30:53:@12267.4]
  wire  valid_38_7; // @[Switch.scala 30:36:@12268.4]
  wire  _T_32308; // @[Switch.scala 30:53:@12270.4]
  wire  valid_38_8; // @[Switch.scala 30:36:@12271.4]
  wire  _T_32311; // @[Switch.scala 30:53:@12273.4]
  wire  valid_38_9; // @[Switch.scala 30:36:@12274.4]
  wire  _T_32314; // @[Switch.scala 30:53:@12276.4]
  wire  valid_38_10; // @[Switch.scala 30:36:@12277.4]
  wire  _T_32317; // @[Switch.scala 30:53:@12279.4]
  wire  valid_38_11; // @[Switch.scala 30:36:@12280.4]
  wire  _T_32320; // @[Switch.scala 30:53:@12282.4]
  wire  valid_38_12; // @[Switch.scala 30:36:@12283.4]
  wire  _T_32323; // @[Switch.scala 30:53:@12285.4]
  wire  valid_38_13; // @[Switch.scala 30:36:@12286.4]
  wire  _T_32326; // @[Switch.scala 30:53:@12288.4]
  wire  valid_38_14; // @[Switch.scala 30:36:@12289.4]
  wire  _T_32329; // @[Switch.scala 30:53:@12291.4]
  wire  valid_38_15; // @[Switch.scala 30:36:@12292.4]
  wire  _T_32332; // @[Switch.scala 30:53:@12294.4]
  wire  valid_38_16; // @[Switch.scala 30:36:@12295.4]
  wire  _T_32335; // @[Switch.scala 30:53:@12297.4]
  wire  valid_38_17; // @[Switch.scala 30:36:@12298.4]
  wire  _T_32338; // @[Switch.scala 30:53:@12300.4]
  wire  valid_38_18; // @[Switch.scala 30:36:@12301.4]
  wire  _T_32341; // @[Switch.scala 30:53:@12303.4]
  wire  valid_38_19; // @[Switch.scala 30:36:@12304.4]
  wire  _T_32344; // @[Switch.scala 30:53:@12306.4]
  wire  valid_38_20; // @[Switch.scala 30:36:@12307.4]
  wire  _T_32347; // @[Switch.scala 30:53:@12309.4]
  wire  valid_38_21; // @[Switch.scala 30:36:@12310.4]
  wire  _T_32350; // @[Switch.scala 30:53:@12312.4]
  wire  valid_38_22; // @[Switch.scala 30:36:@12313.4]
  wire  _T_32353; // @[Switch.scala 30:53:@12315.4]
  wire  valid_38_23; // @[Switch.scala 30:36:@12316.4]
  wire  _T_32356; // @[Switch.scala 30:53:@12318.4]
  wire  valid_38_24; // @[Switch.scala 30:36:@12319.4]
  wire  _T_32359; // @[Switch.scala 30:53:@12321.4]
  wire  valid_38_25; // @[Switch.scala 30:36:@12322.4]
  wire  _T_32362; // @[Switch.scala 30:53:@12324.4]
  wire  valid_38_26; // @[Switch.scala 30:36:@12325.4]
  wire  _T_32365; // @[Switch.scala 30:53:@12327.4]
  wire  valid_38_27; // @[Switch.scala 30:36:@12328.4]
  wire  _T_32368; // @[Switch.scala 30:53:@12330.4]
  wire  valid_38_28; // @[Switch.scala 30:36:@12331.4]
  wire  _T_32371; // @[Switch.scala 30:53:@12333.4]
  wire  valid_38_29; // @[Switch.scala 30:36:@12334.4]
  wire  _T_32374; // @[Switch.scala 30:53:@12336.4]
  wire  valid_38_30; // @[Switch.scala 30:36:@12337.4]
  wire  _T_32377; // @[Switch.scala 30:53:@12339.4]
  wire  valid_38_31; // @[Switch.scala 30:36:@12340.4]
  wire  _T_32380; // @[Switch.scala 30:53:@12342.4]
  wire  valid_38_32; // @[Switch.scala 30:36:@12343.4]
  wire  _T_32383; // @[Switch.scala 30:53:@12345.4]
  wire  valid_38_33; // @[Switch.scala 30:36:@12346.4]
  wire  _T_32386; // @[Switch.scala 30:53:@12348.4]
  wire  valid_38_34; // @[Switch.scala 30:36:@12349.4]
  wire  _T_32389; // @[Switch.scala 30:53:@12351.4]
  wire  valid_38_35; // @[Switch.scala 30:36:@12352.4]
  wire  _T_32392; // @[Switch.scala 30:53:@12354.4]
  wire  valid_38_36; // @[Switch.scala 30:36:@12355.4]
  wire  _T_32395; // @[Switch.scala 30:53:@12357.4]
  wire  valid_38_37; // @[Switch.scala 30:36:@12358.4]
  wire  _T_32398; // @[Switch.scala 30:53:@12360.4]
  wire  valid_38_38; // @[Switch.scala 30:36:@12361.4]
  wire  _T_32401; // @[Switch.scala 30:53:@12363.4]
  wire  valid_38_39; // @[Switch.scala 30:36:@12364.4]
  wire  _T_32404; // @[Switch.scala 30:53:@12366.4]
  wire  valid_38_40; // @[Switch.scala 30:36:@12367.4]
  wire  _T_32407; // @[Switch.scala 30:53:@12369.4]
  wire  valid_38_41; // @[Switch.scala 30:36:@12370.4]
  wire  _T_32410; // @[Switch.scala 30:53:@12372.4]
  wire  valid_38_42; // @[Switch.scala 30:36:@12373.4]
  wire  _T_32413; // @[Switch.scala 30:53:@12375.4]
  wire  valid_38_43; // @[Switch.scala 30:36:@12376.4]
  wire  _T_32416; // @[Switch.scala 30:53:@12378.4]
  wire  valid_38_44; // @[Switch.scala 30:36:@12379.4]
  wire  _T_32419; // @[Switch.scala 30:53:@12381.4]
  wire  valid_38_45; // @[Switch.scala 30:36:@12382.4]
  wire  _T_32422; // @[Switch.scala 30:53:@12384.4]
  wire  valid_38_46; // @[Switch.scala 30:36:@12385.4]
  wire  _T_32425; // @[Switch.scala 30:53:@12387.4]
  wire  valid_38_47; // @[Switch.scala 30:36:@12388.4]
  wire  _T_32428; // @[Switch.scala 30:53:@12390.4]
  wire  valid_38_48; // @[Switch.scala 30:36:@12391.4]
  wire  _T_32431; // @[Switch.scala 30:53:@12393.4]
  wire  valid_38_49; // @[Switch.scala 30:36:@12394.4]
  wire  _T_32434; // @[Switch.scala 30:53:@12396.4]
  wire  valid_38_50; // @[Switch.scala 30:36:@12397.4]
  wire  _T_32437; // @[Switch.scala 30:53:@12399.4]
  wire  valid_38_51; // @[Switch.scala 30:36:@12400.4]
  wire  _T_32440; // @[Switch.scala 30:53:@12402.4]
  wire  valid_38_52; // @[Switch.scala 30:36:@12403.4]
  wire  _T_32443; // @[Switch.scala 30:53:@12405.4]
  wire  valid_38_53; // @[Switch.scala 30:36:@12406.4]
  wire  _T_32446; // @[Switch.scala 30:53:@12408.4]
  wire  valid_38_54; // @[Switch.scala 30:36:@12409.4]
  wire  _T_32449; // @[Switch.scala 30:53:@12411.4]
  wire  valid_38_55; // @[Switch.scala 30:36:@12412.4]
  wire  _T_32452; // @[Switch.scala 30:53:@12414.4]
  wire  valid_38_56; // @[Switch.scala 30:36:@12415.4]
  wire  _T_32455; // @[Switch.scala 30:53:@12417.4]
  wire  valid_38_57; // @[Switch.scala 30:36:@12418.4]
  wire  _T_32458; // @[Switch.scala 30:53:@12420.4]
  wire  valid_38_58; // @[Switch.scala 30:36:@12421.4]
  wire  _T_32461; // @[Switch.scala 30:53:@12423.4]
  wire  valid_38_59; // @[Switch.scala 30:36:@12424.4]
  wire  _T_32464; // @[Switch.scala 30:53:@12426.4]
  wire  valid_38_60; // @[Switch.scala 30:36:@12427.4]
  wire  _T_32467; // @[Switch.scala 30:53:@12429.4]
  wire  valid_38_61; // @[Switch.scala 30:36:@12430.4]
  wire  _T_32470; // @[Switch.scala 30:53:@12432.4]
  wire  valid_38_62; // @[Switch.scala 30:36:@12433.4]
  wire  _T_32473; // @[Switch.scala 30:53:@12435.4]
  wire  valid_38_63; // @[Switch.scala 30:36:@12436.4]
  wire [5:0] _T_32539; // @[Mux.scala 31:69:@12438.4]
  wire [5:0] _T_32540; // @[Mux.scala 31:69:@12439.4]
  wire [5:0] _T_32541; // @[Mux.scala 31:69:@12440.4]
  wire [5:0] _T_32542; // @[Mux.scala 31:69:@12441.4]
  wire [5:0] _T_32543; // @[Mux.scala 31:69:@12442.4]
  wire [5:0] _T_32544; // @[Mux.scala 31:69:@12443.4]
  wire [5:0] _T_32545; // @[Mux.scala 31:69:@12444.4]
  wire [5:0] _T_32546; // @[Mux.scala 31:69:@12445.4]
  wire [5:0] _T_32547; // @[Mux.scala 31:69:@12446.4]
  wire [5:0] _T_32548; // @[Mux.scala 31:69:@12447.4]
  wire [5:0] _T_32549; // @[Mux.scala 31:69:@12448.4]
  wire [5:0] _T_32550; // @[Mux.scala 31:69:@12449.4]
  wire [5:0] _T_32551; // @[Mux.scala 31:69:@12450.4]
  wire [5:0] _T_32552; // @[Mux.scala 31:69:@12451.4]
  wire [5:0] _T_32553; // @[Mux.scala 31:69:@12452.4]
  wire [5:0] _T_32554; // @[Mux.scala 31:69:@12453.4]
  wire [5:0] _T_32555; // @[Mux.scala 31:69:@12454.4]
  wire [5:0] _T_32556; // @[Mux.scala 31:69:@12455.4]
  wire [5:0] _T_32557; // @[Mux.scala 31:69:@12456.4]
  wire [5:0] _T_32558; // @[Mux.scala 31:69:@12457.4]
  wire [5:0] _T_32559; // @[Mux.scala 31:69:@12458.4]
  wire [5:0] _T_32560; // @[Mux.scala 31:69:@12459.4]
  wire [5:0] _T_32561; // @[Mux.scala 31:69:@12460.4]
  wire [5:0] _T_32562; // @[Mux.scala 31:69:@12461.4]
  wire [5:0] _T_32563; // @[Mux.scala 31:69:@12462.4]
  wire [5:0] _T_32564; // @[Mux.scala 31:69:@12463.4]
  wire [5:0] _T_32565; // @[Mux.scala 31:69:@12464.4]
  wire [5:0] _T_32566; // @[Mux.scala 31:69:@12465.4]
  wire [5:0] _T_32567; // @[Mux.scala 31:69:@12466.4]
  wire [5:0] _T_32568; // @[Mux.scala 31:69:@12467.4]
  wire [5:0] _T_32569; // @[Mux.scala 31:69:@12468.4]
  wire [5:0] _T_32570; // @[Mux.scala 31:69:@12469.4]
  wire [5:0] _T_32571; // @[Mux.scala 31:69:@12470.4]
  wire [5:0] _T_32572; // @[Mux.scala 31:69:@12471.4]
  wire [5:0] _T_32573; // @[Mux.scala 31:69:@12472.4]
  wire [5:0] _T_32574; // @[Mux.scala 31:69:@12473.4]
  wire [5:0] _T_32575; // @[Mux.scala 31:69:@12474.4]
  wire [5:0] _T_32576; // @[Mux.scala 31:69:@12475.4]
  wire [5:0] _T_32577; // @[Mux.scala 31:69:@12476.4]
  wire [5:0] _T_32578; // @[Mux.scala 31:69:@12477.4]
  wire [5:0] _T_32579; // @[Mux.scala 31:69:@12478.4]
  wire [5:0] _T_32580; // @[Mux.scala 31:69:@12479.4]
  wire [5:0] _T_32581; // @[Mux.scala 31:69:@12480.4]
  wire [5:0] _T_32582; // @[Mux.scala 31:69:@12481.4]
  wire [5:0] _T_32583; // @[Mux.scala 31:69:@12482.4]
  wire [5:0] _T_32584; // @[Mux.scala 31:69:@12483.4]
  wire [5:0] _T_32585; // @[Mux.scala 31:69:@12484.4]
  wire [5:0] _T_32586; // @[Mux.scala 31:69:@12485.4]
  wire [5:0] _T_32587; // @[Mux.scala 31:69:@12486.4]
  wire [5:0] _T_32588; // @[Mux.scala 31:69:@12487.4]
  wire [5:0] _T_32589; // @[Mux.scala 31:69:@12488.4]
  wire [5:0] _T_32590; // @[Mux.scala 31:69:@12489.4]
  wire [5:0] _T_32591; // @[Mux.scala 31:69:@12490.4]
  wire [5:0] _T_32592; // @[Mux.scala 31:69:@12491.4]
  wire [5:0] _T_32593; // @[Mux.scala 31:69:@12492.4]
  wire [5:0] _T_32594; // @[Mux.scala 31:69:@12493.4]
  wire [5:0] _T_32595; // @[Mux.scala 31:69:@12494.4]
  wire [5:0] _T_32596; // @[Mux.scala 31:69:@12495.4]
  wire [5:0] _T_32597; // @[Mux.scala 31:69:@12496.4]
  wire [5:0] _T_32598; // @[Mux.scala 31:69:@12497.4]
  wire [5:0] _T_32599; // @[Mux.scala 31:69:@12498.4]
  wire [5:0] _T_32600; // @[Mux.scala 31:69:@12499.4]
  wire [5:0] select_38; // @[Mux.scala 31:69:@12500.4]
  wire [47:0] _GEN_2433; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2434; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2435; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2436; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2437; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2438; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2439; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2440; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2441; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2442; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2443; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2444; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2445; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2446; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2447; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2448; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2449; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2450; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2451; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2452; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2453; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2454; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2455; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2456; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2457; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2458; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2459; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2460; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2461; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2462; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2463; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2464; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2465; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2466; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2467; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2468; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2469; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2470; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2471; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2472; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2473; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2474; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2475; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2476; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2477; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2478; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2479; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2480; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2481; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2482; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2483; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2484; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2485; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2486; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2487; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2488; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2489; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2490; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2491; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2492; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2493; // @[Switch.scala 33:19:@12502.4]
  wire [47:0] _GEN_2494; // @[Switch.scala 33:19:@12502.4]
  wire [7:0] _T_32609; // @[Switch.scala 34:32:@12509.4]
  wire [15:0] _T_32617; // @[Switch.scala 34:32:@12517.4]
  wire [7:0] _T_32624; // @[Switch.scala 34:32:@12524.4]
  wire [31:0] _T_32633; // @[Switch.scala 34:32:@12533.4]
  wire [7:0] _T_32640; // @[Switch.scala 34:32:@12540.4]
  wire [15:0] _T_32648; // @[Switch.scala 34:32:@12548.4]
  wire [7:0] _T_32655; // @[Switch.scala 34:32:@12555.4]
  wire [31:0] _T_32664; // @[Switch.scala 34:32:@12564.4]
  wire [63:0] _T_32665; // @[Switch.scala 34:32:@12565.4]
  wire  _T_32669; // @[Switch.scala 30:53:@12568.4]
  wire  valid_39_0; // @[Switch.scala 30:36:@12569.4]
  wire  _T_32672; // @[Switch.scala 30:53:@12571.4]
  wire  valid_39_1; // @[Switch.scala 30:36:@12572.4]
  wire  _T_32675; // @[Switch.scala 30:53:@12574.4]
  wire  valid_39_2; // @[Switch.scala 30:36:@12575.4]
  wire  _T_32678; // @[Switch.scala 30:53:@12577.4]
  wire  valid_39_3; // @[Switch.scala 30:36:@12578.4]
  wire  _T_32681; // @[Switch.scala 30:53:@12580.4]
  wire  valid_39_4; // @[Switch.scala 30:36:@12581.4]
  wire  _T_32684; // @[Switch.scala 30:53:@12583.4]
  wire  valid_39_5; // @[Switch.scala 30:36:@12584.4]
  wire  _T_32687; // @[Switch.scala 30:53:@12586.4]
  wire  valid_39_6; // @[Switch.scala 30:36:@12587.4]
  wire  _T_32690; // @[Switch.scala 30:53:@12589.4]
  wire  valid_39_7; // @[Switch.scala 30:36:@12590.4]
  wire  _T_32693; // @[Switch.scala 30:53:@12592.4]
  wire  valid_39_8; // @[Switch.scala 30:36:@12593.4]
  wire  _T_32696; // @[Switch.scala 30:53:@12595.4]
  wire  valid_39_9; // @[Switch.scala 30:36:@12596.4]
  wire  _T_32699; // @[Switch.scala 30:53:@12598.4]
  wire  valid_39_10; // @[Switch.scala 30:36:@12599.4]
  wire  _T_32702; // @[Switch.scala 30:53:@12601.4]
  wire  valid_39_11; // @[Switch.scala 30:36:@12602.4]
  wire  _T_32705; // @[Switch.scala 30:53:@12604.4]
  wire  valid_39_12; // @[Switch.scala 30:36:@12605.4]
  wire  _T_32708; // @[Switch.scala 30:53:@12607.4]
  wire  valid_39_13; // @[Switch.scala 30:36:@12608.4]
  wire  _T_32711; // @[Switch.scala 30:53:@12610.4]
  wire  valid_39_14; // @[Switch.scala 30:36:@12611.4]
  wire  _T_32714; // @[Switch.scala 30:53:@12613.4]
  wire  valid_39_15; // @[Switch.scala 30:36:@12614.4]
  wire  _T_32717; // @[Switch.scala 30:53:@12616.4]
  wire  valid_39_16; // @[Switch.scala 30:36:@12617.4]
  wire  _T_32720; // @[Switch.scala 30:53:@12619.4]
  wire  valid_39_17; // @[Switch.scala 30:36:@12620.4]
  wire  _T_32723; // @[Switch.scala 30:53:@12622.4]
  wire  valid_39_18; // @[Switch.scala 30:36:@12623.4]
  wire  _T_32726; // @[Switch.scala 30:53:@12625.4]
  wire  valid_39_19; // @[Switch.scala 30:36:@12626.4]
  wire  _T_32729; // @[Switch.scala 30:53:@12628.4]
  wire  valid_39_20; // @[Switch.scala 30:36:@12629.4]
  wire  _T_32732; // @[Switch.scala 30:53:@12631.4]
  wire  valid_39_21; // @[Switch.scala 30:36:@12632.4]
  wire  _T_32735; // @[Switch.scala 30:53:@12634.4]
  wire  valid_39_22; // @[Switch.scala 30:36:@12635.4]
  wire  _T_32738; // @[Switch.scala 30:53:@12637.4]
  wire  valid_39_23; // @[Switch.scala 30:36:@12638.4]
  wire  _T_32741; // @[Switch.scala 30:53:@12640.4]
  wire  valid_39_24; // @[Switch.scala 30:36:@12641.4]
  wire  _T_32744; // @[Switch.scala 30:53:@12643.4]
  wire  valid_39_25; // @[Switch.scala 30:36:@12644.4]
  wire  _T_32747; // @[Switch.scala 30:53:@12646.4]
  wire  valid_39_26; // @[Switch.scala 30:36:@12647.4]
  wire  _T_32750; // @[Switch.scala 30:53:@12649.4]
  wire  valid_39_27; // @[Switch.scala 30:36:@12650.4]
  wire  _T_32753; // @[Switch.scala 30:53:@12652.4]
  wire  valid_39_28; // @[Switch.scala 30:36:@12653.4]
  wire  _T_32756; // @[Switch.scala 30:53:@12655.4]
  wire  valid_39_29; // @[Switch.scala 30:36:@12656.4]
  wire  _T_32759; // @[Switch.scala 30:53:@12658.4]
  wire  valid_39_30; // @[Switch.scala 30:36:@12659.4]
  wire  _T_32762; // @[Switch.scala 30:53:@12661.4]
  wire  valid_39_31; // @[Switch.scala 30:36:@12662.4]
  wire  _T_32765; // @[Switch.scala 30:53:@12664.4]
  wire  valid_39_32; // @[Switch.scala 30:36:@12665.4]
  wire  _T_32768; // @[Switch.scala 30:53:@12667.4]
  wire  valid_39_33; // @[Switch.scala 30:36:@12668.4]
  wire  _T_32771; // @[Switch.scala 30:53:@12670.4]
  wire  valid_39_34; // @[Switch.scala 30:36:@12671.4]
  wire  _T_32774; // @[Switch.scala 30:53:@12673.4]
  wire  valid_39_35; // @[Switch.scala 30:36:@12674.4]
  wire  _T_32777; // @[Switch.scala 30:53:@12676.4]
  wire  valid_39_36; // @[Switch.scala 30:36:@12677.4]
  wire  _T_32780; // @[Switch.scala 30:53:@12679.4]
  wire  valid_39_37; // @[Switch.scala 30:36:@12680.4]
  wire  _T_32783; // @[Switch.scala 30:53:@12682.4]
  wire  valid_39_38; // @[Switch.scala 30:36:@12683.4]
  wire  _T_32786; // @[Switch.scala 30:53:@12685.4]
  wire  valid_39_39; // @[Switch.scala 30:36:@12686.4]
  wire  _T_32789; // @[Switch.scala 30:53:@12688.4]
  wire  valid_39_40; // @[Switch.scala 30:36:@12689.4]
  wire  _T_32792; // @[Switch.scala 30:53:@12691.4]
  wire  valid_39_41; // @[Switch.scala 30:36:@12692.4]
  wire  _T_32795; // @[Switch.scala 30:53:@12694.4]
  wire  valid_39_42; // @[Switch.scala 30:36:@12695.4]
  wire  _T_32798; // @[Switch.scala 30:53:@12697.4]
  wire  valid_39_43; // @[Switch.scala 30:36:@12698.4]
  wire  _T_32801; // @[Switch.scala 30:53:@12700.4]
  wire  valid_39_44; // @[Switch.scala 30:36:@12701.4]
  wire  _T_32804; // @[Switch.scala 30:53:@12703.4]
  wire  valid_39_45; // @[Switch.scala 30:36:@12704.4]
  wire  _T_32807; // @[Switch.scala 30:53:@12706.4]
  wire  valid_39_46; // @[Switch.scala 30:36:@12707.4]
  wire  _T_32810; // @[Switch.scala 30:53:@12709.4]
  wire  valid_39_47; // @[Switch.scala 30:36:@12710.4]
  wire  _T_32813; // @[Switch.scala 30:53:@12712.4]
  wire  valid_39_48; // @[Switch.scala 30:36:@12713.4]
  wire  _T_32816; // @[Switch.scala 30:53:@12715.4]
  wire  valid_39_49; // @[Switch.scala 30:36:@12716.4]
  wire  _T_32819; // @[Switch.scala 30:53:@12718.4]
  wire  valid_39_50; // @[Switch.scala 30:36:@12719.4]
  wire  _T_32822; // @[Switch.scala 30:53:@12721.4]
  wire  valid_39_51; // @[Switch.scala 30:36:@12722.4]
  wire  _T_32825; // @[Switch.scala 30:53:@12724.4]
  wire  valid_39_52; // @[Switch.scala 30:36:@12725.4]
  wire  _T_32828; // @[Switch.scala 30:53:@12727.4]
  wire  valid_39_53; // @[Switch.scala 30:36:@12728.4]
  wire  _T_32831; // @[Switch.scala 30:53:@12730.4]
  wire  valid_39_54; // @[Switch.scala 30:36:@12731.4]
  wire  _T_32834; // @[Switch.scala 30:53:@12733.4]
  wire  valid_39_55; // @[Switch.scala 30:36:@12734.4]
  wire  _T_32837; // @[Switch.scala 30:53:@12736.4]
  wire  valid_39_56; // @[Switch.scala 30:36:@12737.4]
  wire  _T_32840; // @[Switch.scala 30:53:@12739.4]
  wire  valid_39_57; // @[Switch.scala 30:36:@12740.4]
  wire  _T_32843; // @[Switch.scala 30:53:@12742.4]
  wire  valid_39_58; // @[Switch.scala 30:36:@12743.4]
  wire  _T_32846; // @[Switch.scala 30:53:@12745.4]
  wire  valid_39_59; // @[Switch.scala 30:36:@12746.4]
  wire  _T_32849; // @[Switch.scala 30:53:@12748.4]
  wire  valid_39_60; // @[Switch.scala 30:36:@12749.4]
  wire  _T_32852; // @[Switch.scala 30:53:@12751.4]
  wire  valid_39_61; // @[Switch.scala 30:36:@12752.4]
  wire  _T_32855; // @[Switch.scala 30:53:@12754.4]
  wire  valid_39_62; // @[Switch.scala 30:36:@12755.4]
  wire  _T_32858; // @[Switch.scala 30:53:@12757.4]
  wire  valid_39_63; // @[Switch.scala 30:36:@12758.4]
  wire [5:0] _T_32924; // @[Mux.scala 31:69:@12760.4]
  wire [5:0] _T_32925; // @[Mux.scala 31:69:@12761.4]
  wire [5:0] _T_32926; // @[Mux.scala 31:69:@12762.4]
  wire [5:0] _T_32927; // @[Mux.scala 31:69:@12763.4]
  wire [5:0] _T_32928; // @[Mux.scala 31:69:@12764.4]
  wire [5:0] _T_32929; // @[Mux.scala 31:69:@12765.4]
  wire [5:0] _T_32930; // @[Mux.scala 31:69:@12766.4]
  wire [5:0] _T_32931; // @[Mux.scala 31:69:@12767.4]
  wire [5:0] _T_32932; // @[Mux.scala 31:69:@12768.4]
  wire [5:0] _T_32933; // @[Mux.scala 31:69:@12769.4]
  wire [5:0] _T_32934; // @[Mux.scala 31:69:@12770.4]
  wire [5:0] _T_32935; // @[Mux.scala 31:69:@12771.4]
  wire [5:0] _T_32936; // @[Mux.scala 31:69:@12772.4]
  wire [5:0] _T_32937; // @[Mux.scala 31:69:@12773.4]
  wire [5:0] _T_32938; // @[Mux.scala 31:69:@12774.4]
  wire [5:0] _T_32939; // @[Mux.scala 31:69:@12775.4]
  wire [5:0] _T_32940; // @[Mux.scala 31:69:@12776.4]
  wire [5:0] _T_32941; // @[Mux.scala 31:69:@12777.4]
  wire [5:0] _T_32942; // @[Mux.scala 31:69:@12778.4]
  wire [5:0] _T_32943; // @[Mux.scala 31:69:@12779.4]
  wire [5:0] _T_32944; // @[Mux.scala 31:69:@12780.4]
  wire [5:0] _T_32945; // @[Mux.scala 31:69:@12781.4]
  wire [5:0] _T_32946; // @[Mux.scala 31:69:@12782.4]
  wire [5:0] _T_32947; // @[Mux.scala 31:69:@12783.4]
  wire [5:0] _T_32948; // @[Mux.scala 31:69:@12784.4]
  wire [5:0] _T_32949; // @[Mux.scala 31:69:@12785.4]
  wire [5:0] _T_32950; // @[Mux.scala 31:69:@12786.4]
  wire [5:0] _T_32951; // @[Mux.scala 31:69:@12787.4]
  wire [5:0] _T_32952; // @[Mux.scala 31:69:@12788.4]
  wire [5:0] _T_32953; // @[Mux.scala 31:69:@12789.4]
  wire [5:0] _T_32954; // @[Mux.scala 31:69:@12790.4]
  wire [5:0] _T_32955; // @[Mux.scala 31:69:@12791.4]
  wire [5:0] _T_32956; // @[Mux.scala 31:69:@12792.4]
  wire [5:0] _T_32957; // @[Mux.scala 31:69:@12793.4]
  wire [5:0] _T_32958; // @[Mux.scala 31:69:@12794.4]
  wire [5:0] _T_32959; // @[Mux.scala 31:69:@12795.4]
  wire [5:0] _T_32960; // @[Mux.scala 31:69:@12796.4]
  wire [5:0] _T_32961; // @[Mux.scala 31:69:@12797.4]
  wire [5:0] _T_32962; // @[Mux.scala 31:69:@12798.4]
  wire [5:0] _T_32963; // @[Mux.scala 31:69:@12799.4]
  wire [5:0] _T_32964; // @[Mux.scala 31:69:@12800.4]
  wire [5:0] _T_32965; // @[Mux.scala 31:69:@12801.4]
  wire [5:0] _T_32966; // @[Mux.scala 31:69:@12802.4]
  wire [5:0] _T_32967; // @[Mux.scala 31:69:@12803.4]
  wire [5:0] _T_32968; // @[Mux.scala 31:69:@12804.4]
  wire [5:0] _T_32969; // @[Mux.scala 31:69:@12805.4]
  wire [5:0] _T_32970; // @[Mux.scala 31:69:@12806.4]
  wire [5:0] _T_32971; // @[Mux.scala 31:69:@12807.4]
  wire [5:0] _T_32972; // @[Mux.scala 31:69:@12808.4]
  wire [5:0] _T_32973; // @[Mux.scala 31:69:@12809.4]
  wire [5:0] _T_32974; // @[Mux.scala 31:69:@12810.4]
  wire [5:0] _T_32975; // @[Mux.scala 31:69:@12811.4]
  wire [5:0] _T_32976; // @[Mux.scala 31:69:@12812.4]
  wire [5:0] _T_32977; // @[Mux.scala 31:69:@12813.4]
  wire [5:0] _T_32978; // @[Mux.scala 31:69:@12814.4]
  wire [5:0] _T_32979; // @[Mux.scala 31:69:@12815.4]
  wire [5:0] _T_32980; // @[Mux.scala 31:69:@12816.4]
  wire [5:0] _T_32981; // @[Mux.scala 31:69:@12817.4]
  wire [5:0] _T_32982; // @[Mux.scala 31:69:@12818.4]
  wire [5:0] _T_32983; // @[Mux.scala 31:69:@12819.4]
  wire [5:0] _T_32984; // @[Mux.scala 31:69:@12820.4]
  wire [5:0] _T_32985; // @[Mux.scala 31:69:@12821.4]
  wire [5:0] select_39; // @[Mux.scala 31:69:@12822.4]
  wire [47:0] _GEN_2497; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2498; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2499; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2500; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2501; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2502; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2503; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2504; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2505; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2506; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2507; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2508; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2509; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2510; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2511; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2512; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2513; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2514; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2515; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2516; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2517; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2518; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2519; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2520; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2521; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2522; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2523; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2524; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2525; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2526; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2527; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2528; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2529; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2530; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2531; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2532; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2533; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2534; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2535; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2536; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2537; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2538; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2539; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2540; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2541; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2542; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2543; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2544; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2545; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2546; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2547; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2548; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2549; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2550; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2551; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2552; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2553; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2554; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2555; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2556; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2557; // @[Switch.scala 33:19:@12824.4]
  wire [47:0] _GEN_2558; // @[Switch.scala 33:19:@12824.4]
  wire [7:0] _T_32994; // @[Switch.scala 34:32:@12831.4]
  wire [15:0] _T_33002; // @[Switch.scala 34:32:@12839.4]
  wire [7:0] _T_33009; // @[Switch.scala 34:32:@12846.4]
  wire [31:0] _T_33018; // @[Switch.scala 34:32:@12855.4]
  wire [7:0] _T_33025; // @[Switch.scala 34:32:@12862.4]
  wire [15:0] _T_33033; // @[Switch.scala 34:32:@12870.4]
  wire [7:0] _T_33040; // @[Switch.scala 34:32:@12877.4]
  wire [31:0] _T_33049; // @[Switch.scala 34:32:@12886.4]
  wire [63:0] _T_33050; // @[Switch.scala 34:32:@12887.4]
  wire  _T_33054; // @[Switch.scala 30:53:@12890.4]
  wire  valid_40_0; // @[Switch.scala 30:36:@12891.4]
  wire  _T_33057; // @[Switch.scala 30:53:@12893.4]
  wire  valid_40_1; // @[Switch.scala 30:36:@12894.4]
  wire  _T_33060; // @[Switch.scala 30:53:@12896.4]
  wire  valid_40_2; // @[Switch.scala 30:36:@12897.4]
  wire  _T_33063; // @[Switch.scala 30:53:@12899.4]
  wire  valid_40_3; // @[Switch.scala 30:36:@12900.4]
  wire  _T_33066; // @[Switch.scala 30:53:@12902.4]
  wire  valid_40_4; // @[Switch.scala 30:36:@12903.4]
  wire  _T_33069; // @[Switch.scala 30:53:@12905.4]
  wire  valid_40_5; // @[Switch.scala 30:36:@12906.4]
  wire  _T_33072; // @[Switch.scala 30:53:@12908.4]
  wire  valid_40_6; // @[Switch.scala 30:36:@12909.4]
  wire  _T_33075; // @[Switch.scala 30:53:@12911.4]
  wire  valid_40_7; // @[Switch.scala 30:36:@12912.4]
  wire  _T_33078; // @[Switch.scala 30:53:@12914.4]
  wire  valid_40_8; // @[Switch.scala 30:36:@12915.4]
  wire  _T_33081; // @[Switch.scala 30:53:@12917.4]
  wire  valid_40_9; // @[Switch.scala 30:36:@12918.4]
  wire  _T_33084; // @[Switch.scala 30:53:@12920.4]
  wire  valid_40_10; // @[Switch.scala 30:36:@12921.4]
  wire  _T_33087; // @[Switch.scala 30:53:@12923.4]
  wire  valid_40_11; // @[Switch.scala 30:36:@12924.4]
  wire  _T_33090; // @[Switch.scala 30:53:@12926.4]
  wire  valid_40_12; // @[Switch.scala 30:36:@12927.4]
  wire  _T_33093; // @[Switch.scala 30:53:@12929.4]
  wire  valid_40_13; // @[Switch.scala 30:36:@12930.4]
  wire  _T_33096; // @[Switch.scala 30:53:@12932.4]
  wire  valid_40_14; // @[Switch.scala 30:36:@12933.4]
  wire  _T_33099; // @[Switch.scala 30:53:@12935.4]
  wire  valid_40_15; // @[Switch.scala 30:36:@12936.4]
  wire  _T_33102; // @[Switch.scala 30:53:@12938.4]
  wire  valid_40_16; // @[Switch.scala 30:36:@12939.4]
  wire  _T_33105; // @[Switch.scala 30:53:@12941.4]
  wire  valid_40_17; // @[Switch.scala 30:36:@12942.4]
  wire  _T_33108; // @[Switch.scala 30:53:@12944.4]
  wire  valid_40_18; // @[Switch.scala 30:36:@12945.4]
  wire  _T_33111; // @[Switch.scala 30:53:@12947.4]
  wire  valid_40_19; // @[Switch.scala 30:36:@12948.4]
  wire  _T_33114; // @[Switch.scala 30:53:@12950.4]
  wire  valid_40_20; // @[Switch.scala 30:36:@12951.4]
  wire  _T_33117; // @[Switch.scala 30:53:@12953.4]
  wire  valid_40_21; // @[Switch.scala 30:36:@12954.4]
  wire  _T_33120; // @[Switch.scala 30:53:@12956.4]
  wire  valid_40_22; // @[Switch.scala 30:36:@12957.4]
  wire  _T_33123; // @[Switch.scala 30:53:@12959.4]
  wire  valid_40_23; // @[Switch.scala 30:36:@12960.4]
  wire  _T_33126; // @[Switch.scala 30:53:@12962.4]
  wire  valid_40_24; // @[Switch.scala 30:36:@12963.4]
  wire  _T_33129; // @[Switch.scala 30:53:@12965.4]
  wire  valid_40_25; // @[Switch.scala 30:36:@12966.4]
  wire  _T_33132; // @[Switch.scala 30:53:@12968.4]
  wire  valid_40_26; // @[Switch.scala 30:36:@12969.4]
  wire  _T_33135; // @[Switch.scala 30:53:@12971.4]
  wire  valid_40_27; // @[Switch.scala 30:36:@12972.4]
  wire  _T_33138; // @[Switch.scala 30:53:@12974.4]
  wire  valid_40_28; // @[Switch.scala 30:36:@12975.4]
  wire  _T_33141; // @[Switch.scala 30:53:@12977.4]
  wire  valid_40_29; // @[Switch.scala 30:36:@12978.4]
  wire  _T_33144; // @[Switch.scala 30:53:@12980.4]
  wire  valid_40_30; // @[Switch.scala 30:36:@12981.4]
  wire  _T_33147; // @[Switch.scala 30:53:@12983.4]
  wire  valid_40_31; // @[Switch.scala 30:36:@12984.4]
  wire  _T_33150; // @[Switch.scala 30:53:@12986.4]
  wire  valid_40_32; // @[Switch.scala 30:36:@12987.4]
  wire  _T_33153; // @[Switch.scala 30:53:@12989.4]
  wire  valid_40_33; // @[Switch.scala 30:36:@12990.4]
  wire  _T_33156; // @[Switch.scala 30:53:@12992.4]
  wire  valid_40_34; // @[Switch.scala 30:36:@12993.4]
  wire  _T_33159; // @[Switch.scala 30:53:@12995.4]
  wire  valid_40_35; // @[Switch.scala 30:36:@12996.4]
  wire  _T_33162; // @[Switch.scala 30:53:@12998.4]
  wire  valid_40_36; // @[Switch.scala 30:36:@12999.4]
  wire  _T_33165; // @[Switch.scala 30:53:@13001.4]
  wire  valid_40_37; // @[Switch.scala 30:36:@13002.4]
  wire  _T_33168; // @[Switch.scala 30:53:@13004.4]
  wire  valid_40_38; // @[Switch.scala 30:36:@13005.4]
  wire  _T_33171; // @[Switch.scala 30:53:@13007.4]
  wire  valid_40_39; // @[Switch.scala 30:36:@13008.4]
  wire  _T_33174; // @[Switch.scala 30:53:@13010.4]
  wire  valid_40_40; // @[Switch.scala 30:36:@13011.4]
  wire  _T_33177; // @[Switch.scala 30:53:@13013.4]
  wire  valid_40_41; // @[Switch.scala 30:36:@13014.4]
  wire  _T_33180; // @[Switch.scala 30:53:@13016.4]
  wire  valid_40_42; // @[Switch.scala 30:36:@13017.4]
  wire  _T_33183; // @[Switch.scala 30:53:@13019.4]
  wire  valid_40_43; // @[Switch.scala 30:36:@13020.4]
  wire  _T_33186; // @[Switch.scala 30:53:@13022.4]
  wire  valid_40_44; // @[Switch.scala 30:36:@13023.4]
  wire  _T_33189; // @[Switch.scala 30:53:@13025.4]
  wire  valid_40_45; // @[Switch.scala 30:36:@13026.4]
  wire  _T_33192; // @[Switch.scala 30:53:@13028.4]
  wire  valid_40_46; // @[Switch.scala 30:36:@13029.4]
  wire  _T_33195; // @[Switch.scala 30:53:@13031.4]
  wire  valid_40_47; // @[Switch.scala 30:36:@13032.4]
  wire  _T_33198; // @[Switch.scala 30:53:@13034.4]
  wire  valid_40_48; // @[Switch.scala 30:36:@13035.4]
  wire  _T_33201; // @[Switch.scala 30:53:@13037.4]
  wire  valid_40_49; // @[Switch.scala 30:36:@13038.4]
  wire  _T_33204; // @[Switch.scala 30:53:@13040.4]
  wire  valid_40_50; // @[Switch.scala 30:36:@13041.4]
  wire  _T_33207; // @[Switch.scala 30:53:@13043.4]
  wire  valid_40_51; // @[Switch.scala 30:36:@13044.4]
  wire  _T_33210; // @[Switch.scala 30:53:@13046.4]
  wire  valid_40_52; // @[Switch.scala 30:36:@13047.4]
  wire  _T_33213; // @[Switch.scala 30:53:@13049.4]
  wire  valid_40_53; // @[Switch.scala 30:36:@13050.4]
  wire  _T_33216; // @[Switch.scala 30:53:@13052.4]
  wire  valid_40_54; // @[Switch.scala 30:36:@13053.4]
  wire  _T_33219; // @[Switch.scala 30:53:@13055.4]
  wire  valid_40_55; // @[Switch.scala 30:36:@13056.4]
  wire  _T_33222; // @[Switch.scala 30:53:@13058.4]
  wire  valid_40_56; // @[Switch.scala 30:36:@13059.4]
  wire  _T_33225; // @[Switch.scala 30:53:@13061.4]
  wire  valid_40_57; // @[Switch.scala 30:36:@13062.4]
  wire  _T_33228; // @[Switch.scala 30:53:@13064.4]
  wire  valid_40_58; // @[Switch.scala 30:36:@13065.4]
  wire  _T_33231; // @[Switch.scala 30:53:@13067.4]
  wire  valid_40_59; // @[Switch.scala 30:36:@13068.4]
  wire  _T_33234; // @[Switch.scala 30:53:@13070.4]
  wire  valid_40_60; // @[Switch.scala 30:36:@13071.4]
  wire  _T_33237; // @[Switch.scala 30:53:@13073.4]
  wire  valid_40_61; // @[Switch.scala 30:36:@13074.4]
  wire  _T_33240; // @[Switch.scala 30:53:@13076.4]
  wire  valid_40_62; // @[Switch.scala 30:36:@13077.4]
  wire  _T_33243; // @[Switch.scala 30:53:@13079.4]
  wire  valid_40_63; // @[Switch.scala 30:36:@13080.4]
  wire [5:0] _T_33309; // @[Mux.scala 31:69:@13082.4]
  wire [5:0] _T_33310; // @[Mux.scala 31:69:@13083.4]
  wire [5:0] _T_33311; // @[Mux.scala 31:69:@13084.4]
  wire [5:0] _T_33312; // @[Mux.scala 31:69:@13085.4]
  wire [5:0] _T_33313; // @[Mux.scala 31:69:@13086.4]
  wire [5:0] _T_33314; // @[Mux.scala 31:69:@13087.4]
  wire [5:0] _T_33315; // @[Mux.scala 31:69:@13088.4]
  wire [5:0] _T_33316; // @[Mux.scala 31:69:@13089.4]
  wire [5:0] _T_33317; // @[Mux.scala 31:69:@13090.4]
  wire [5:0] _T_33318; // @[Mux.scala 31:69:@13091.4]
  wire [5:0] _T_33319; // @[Mux.scala 31:69:@13092.4]
  wire [5:0] _T_33320; // @[Mux.scala 31:69:@13093.4]
  wire [5:0] _T_33321; // @[Mux.scala 31:69:@13094.4]
  wire [5:0] _T_33322; // @[Mux.scala 31:69:@13095.4]
  wire [5:0] _T_33323; // @[Mux.scala 31:69:@13096.4]
  wire [5:0] _T_33324; // @[Mux.scala 31:69:@13097.4]
  wire [5:0] _T_33325; // @[Mux.scala 31:69:@13098.4]
  wire [5:0] _T_33326; // @[Mux.scala 31:69:@13099.4]
  wire [5:0] _T_33327; // @[Mux.scala 31:69:@13100.4]
  wire [5:0] _T_33328; // @[Mux.scala 31:69:@13101.4]
  wire [5:0] _T_33329; // @[Mux.scala 31:69:@13102.4]
  wire [5:0] _T_33330; // @[Mux.scala 31:69:@13103.4]
  wire [5:0] _T_33331; // @[Mux.scala 31:69:@13104.4]
  wire [5:0] _T_33332; // @[Mux.scala 31:69:@13105.4]
  wire [5:0] _T_33333; // @[Mux.scala 31:69:@13106.4]
  wire [5:0] _T_33334; // @[Mux.scala 31:69:@13107.4]
  wire [5:0] _T_33335; // @[Mux.scala 31:69:@13108.4]
  wire [5:0] _T_33336; // @[Mux.scala 31:69:@13109.4]
  wire [5:0] _T_33337; // @[Mux.scala 31:69:@13110.4]
  wire [5:0] _T_33338; // @[Mux.scala 31:69:@13111.4]
  wire [5:0] _T_33339; // @[Mux.scala 31:69:@13112.4]
  wire [5:0] _T_33340; // @[Mux.scala 31:69:@13113.4]
  wire [5:0] _T_33341; // @[Mux.scala 31:69:@13114.4]
  wire [5:0] _T_33342; // @[Mux.scala 31:69:@13115.4]
  wire [5:0] _T_33343; // @[Mux.scala 31:69:@13116.4]
  wire [5:0] _T_33344; // @[Mux.scala 31:69:@13117.4]
  wire [5:0] _T_33345; // @[Mux.scala 31:69:@13118.4]
  wire [5:0] _T_33346; // @[Mux.scala 31:69:@13119.4]
  wire [5:0] _T_33347; // @[Mux.scala 31:69:@13120.4]
  wire [5:0] _T_33348; // @[Mux.scala 31:69:@13121.4]
  wire [5:0] _T_33349; // @[Mux.scala 31:69:@13122.4]
  wire [5:0] _T_33350; // @[Mux.scala 31:69:@13123.4]
  wire [5:0] _T_33351; // @[Mux.scala 31:69:@13124.4]
  wire [5:0] _T_33352; // @[Mux.scala 31:69:@13125.4]
  wire [5:0] _T_33353; // @[Mux.scala 31:69:@13126.4]
  wire [5:0] _T_33354; // @[Mux.scala 31:69:@13127.4]
  wire [5:0] _T_33355; // @[Mux.scala 31:69:@13128.4]
  wire [5:0] _T_33356; // @[Mux.scala 31:69:@13129.4]
  wire [5:0] _T_33357; // @[Mux.scala 31:69:@13130.4]
  wire [5:0] _T_33358; // @[Mux.scala 31:69:@13131.4]
  wire [5:0] _T_33359; // @[Mux.scala 31:69:@13132.4]
  wire [5:0] _T_33360; // @[Mux.scala 31:69:@13133.4]
  wire [5:0] _T_33361; // @[Mux.scala 31:69:@13134.4]
  wire [5:0] _T_33362; // @[Mux.scala 31:69:@13135.4]
  wire [5:0] _T_33363; // @[Mux.scala 31:69:@13136.4]
  wire [5:0] _T_33364; // @[Mux.scala 31:69:@13137.4]
  wire [5:0] _T_33365; // @[Mux.scala 31:69:@13138.4]
  wire [5:0] _T_33366; // @[Mux.scala 31:69:@13139.4]
  wire [5:0] _T_33367; // @[Mux.scala 31:69:@13140.4]
  wire [5:0] _T_33368; // @[Mux.scala 31:69:@13141.4]
  wire [5:0] _T_33369; // @[Mux.scala 31:69:@13142.4]
  wire [5:0] _T_33370; // @[Mux.scala 31:69:@13143.4]
  wire [5:0] select_40; // @[Mux.scala 31:69:@13144.4]
  wire [47:0] _GEN_2561; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2562; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2563; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2564; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2565; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2566; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2567; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2568; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2569; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2570; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2571; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2572; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2573; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2574; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2575; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2576; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2577; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2578; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2579; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2580; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2581; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2582; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2583; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2584; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2585; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2586; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2587; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2588; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2589; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2590; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2591; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2592; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2593; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2594; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2595; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2596; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2597; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2598; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2599; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2600; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2601; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2602; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2603; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2604; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2605; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2606; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2607; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2608; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2609; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2610; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2611; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2612; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2613; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2614; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2615; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2616; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2617; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2618; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2619; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2620; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2621; // @[Switch.scala 33:19:@13146.4]
  wire [47:0] _GEN_2622; // @[Switch.scala 33:19:@13146.4]
  wire [7:0] _T_33379; // @[Switch.scala 34:32:@13153.4]
  wire [15:0] _T_33387; // @[Switch.scala 34:32:@13161.4]
  wire [7:0] _T_33394; // @[Switch.scala 34:32:@13168.4]
  wire [31:0] _T_33403; // @[Switch.scala 34:32:@13177.4]
  wire [7:0] _T_33410; // @[Switch.scala 34:32:@13184.4]
  wire [15:0] _T_33418; // @[Switch.scala 34:32:@13192.4]
  wire [7:0] _T_33425; // @[Switch.scala 34:32:@13199.4]
  wire [31:0] _T_33434; // @[Switch.scala 34:32:@13208.4]
  wire [63:0] _T_33435; // @[Switch.scala 34:32:@13209.4]
  wire  _T_33439; // @[Switch.scala 30:53:@13212.4]
  wire  valid_41_0; // @[Switch.scala 30:36:@13213.4]
  wire  _T_33442; // @[Switch.scala 30:53:@13215.4]
  wire  valid_41_1; // @[Switch.scala 30:36:@13216.4]
  wire  _T_33445; // @[Switch.scala 30:53:@13218.4]
  wire  valid_41_2; // @[Switch.scala 30:36:@13219.4]
  wire  _T_33448; // @[Switch.scala 30:53:@13221.4]
  wire  valid_41_3; // @[Switch.scala 30:36:@13222.4]
  wire  _T_33451; // @[Switch.scala 30:53:@13224.4]
  wire  valid_41_4; // @[Switch.scala 30:36:@13225.4]
  wire  _T_33454; // @[Switch.scala 30:53:@13227.4]
  wire  valid_41_5; // @[Switch.scala 30:36:@13228.4]
  wire  _T_33457; // @[Switch.scala 30:53:@13230.4]
  wire  valid_41_6; // @[Switch.scala 30:36:@13231.4]
  wire  _T_33460; // @[Switch.scala 30:53:@13233.4]
  wire  valid_41_7; // @[Switch.scala 30:36:@13234.4]
  wire  _T_33463; // @[Switch.scala 30:53:@13236.4]
  wire  valid_41_8; // @[Switch.scala 30:36:@13237.4]
  wire  _T_33466; // @[Switch.scala 30:53:@13239.4]
  wire  valid_41_9; // @[Switch.scala 30:36:@13240.4]
  wire  _T_33469; // @[Switch.scala 30:53:@13242.4]
  wire  valid_41_10; // @[Switch.scala 30:36:@13243.4]
  wire  _T_33472; // @[Switch.scala 30:53:@13245.4]
  wire  valid_41_11; // @[Switch.scala 30:36:@13246.4]
  wire  _T_33475; // @[Switch.scala 30:53:@13248.4]
  wire  valid_41_12; // @[Switch.scala 30:36:@13249.4]
  wire  _T_33478; // @[Switch.scala 30:53:@13251.4]
  wire  valid_41_13; // @[Switch.scala 30:36:@13252.4]
  wire  _T_33481; // @[Switch.scala 30:53:@13254.4]
  wire  valid_41_14; // @[Switch.scala 30:36:@13255.4]
  wire  _T_33484; // @[Switch.scala 30:53:@13257.4]
  wire  valid_41_15; // @[Switch.scala 30:36:@13258.4]
  wire  _T_33487; // @[Switch.scala 30:53:@13260.4]
  wire  valid_41_16; // @[Switch.scala 30:36:@13261.4]
  wire  _T_33490; // @[Switch.scala 30:53:@13263.4]
  wire  valid_41_17; // @[Switch.scala 30:36:@13264.4]
  wire  _T_33493; // @[Switch.scala 30:53:@13266.4]
  wire  valid_41_18; // @[Switch.scala 30:36:@13267.4]
  wire  _T_33496; // @[Switch.scala 30:53:@13269.4]
  wire  valid_41_19; // @[Switch.scala 30:36:@13270.4]
  wire  _T_33499; // @[Switch.scala 30:53:@13272.4]
  wire  valid_41_20; // @[Switch.scala 30:36:@13273.4]
  wire  _T_33502; // @[Switch.scala 30:53:@13275.4]
  wire  valid_41_21; // @[Switch.scala 30:36:@13276.4]
  wire  _T_33505; // @[Switch.scala 30:53:@13278.4]
  wire  valid_41_22; // @[Switch.scala 30:36:@13279.4]
  wire  _T_33508; // @[Switch.scala 30:53:@13281.4]
  wire  valid_41_23; // @[Switch.scala 30:36:@13282.4]
  wire  _T_33511; // @[Switch.scala 30:53:@13284.4]
  wire  valid_41_24; // @[Switch.scala 30:36:@13285.4]
  wire  _T_33514; // @[Switch.scala 30:53:@13287.4]
  wire  valid_41_25; // @[Switch.scala 30:36:@13288.4]
  wire  _T_33517; // @[Switch.scala 30:53:@13290.4]
  wire  valid_41_26; // @[Switch.scala 30:36:@13291.4]
  wire  _T_33520; // @[Switch.scala 30:53:@13293.4]
  wire  valid_41_27; // @[Switch.scala 30:36:@13294.4]
  wire  _T_33523; // @[Switch.scala 30:53:@13296.4]
  wire  valid_41_28; // @[Switch.scala 30:36:@13297.4]
  wire  _T_33526; // @[Switch.scala 30:53:@13299.4]
  wire  valid_41_29; // @[Switch.scala 30:36:@13300.4]
  wire  _T_33529; // @[Switch.scala 30:53:@13302.4]
  wire  valid_41_30; // @[Switch.scala 30:36:@13303.4]
  wire  _T_33532; // @[Switch.scala 30:53:@13305.4]
  wire  valid_41_31; // @[Switch.scala 30:36:@13306.4]
  wire  _T_33535; // @[Switch.scala 30:53:@13308.4]
  wire  valid_41_32; // @[Switch.scala 30:36:@13309.4]
  wire  _T_33538; // @[Switch.scala 30:53:@13311.4]
  wire  valid_41_33; // @[Switch.scala 30:36:@13312.4]
  wire  _T_33541; // @[Switch.scala 30:53:@13314.4]
  wire  valid_41_34; // @[Switch.scala 30:36:@13315.4]
  wire  _T_33544; // @[Switch.scala 30:53:@13317.4]
  wire  valid_41_35; // @[Switch.scala 30:36:@13318.4]
  wire  _T_33547; // @[Switch.scala 30:53:@13320.4]
  wire  valid_41_36; // @[Switch.scala 30:36:@13321.4]
  wire  _T_33550; // @[Switch.scala 30:53:@13323.4]
  wire  valid_41_37; // @[Switch.scala 30:36:@13324.4]
  wire  _T_33553; // @[Switch.scala 30:53:@13326.4]
  wire  valid_41_38; // @[Switch.scala 30:36:@13327.4]
  wire  _T_33556; // @[Switch.scala 30:53:@13329.4]
  wire  valid_41_39; // @[Switch.scala 30:36:@13330.4]
  wire  _T_33559; // @[Switch.scala 30:53:@13332.4]
  wire  valid_41_40; // @[Switch.scala 30:36:@13333.4]
  wire  _T_33562; // @[Switch.scala 30:53:@13335.4]
  wire  valid_41_41; // @[Switch.scala 30:36:@13336.4]
  wire  _T_33565; // @[Switch.scala 30:53:@13338.4]
  wire  valid_41_42; // @[Switch.scala 30:36:@13339.4]
  wire  _T_33568; // @[Switch.scala 30:53:@13341.4]
  wire  valid_41_43; // @[Switch.scala 30:36:@13342.4]
  wire  _T_33571; // @[Switch.scala 30:53:@13344.4]
  wire  valid_41_44; // @[Switch.scala 30:36:@13345.4]
  wire  _T_33574; // @[Switch.scala 30:53:@13347.4]
  wire  valid_41_45; // @[Switch.scala 30:36:@13348.4]
  wire  _T_33577; // @[Switch.scala 30:53:@13350.4]
  wire  valid_41_46; // @[Switch.scala 30:36:@13351.4]
  wire  _T_33580; // @[Switch.scala 30:53:@13353.4]
  wire  valid_41_47; // @[Switch.scala 30:36:@13354.4]
  wire  _T_33583; // @[Switch.scala 30:53:@13356.4]
  wire  valid_41_48; // @[Switch.scala 30:36:@13357.4]
  wire  _T_33586; // @[Switch.scala 30:53:@13359.4]
  wire  valid_41_49; // @[Switch.scala 30:36:@13360.4]
  wire  _T_33589; // @[Switch.scala 30:53:@13362.4]
  wire  valid_41_50; // @[Switch.scala 30:36:@13363.4]
  wire  _T_33592; // @[Switch.scala 30:53:@13365.4]
  wire  valid_41_51; // @[Switch.scala 30:36:@13366.4]
  wire  _T_33595; // @[Switch.scala 30:53:@13368.4]
  wire  valid_41_52; // @[Switch.scala 30:36:@13369.4]
  wire  _T_33598; // @[Switch.scala 30:53:@13371.4]
  wire  valid_41_53; // @[Switch.scala 30:36:@13372.4]
  wire  _T_33601; // @[Switch.scala 30:53:@13374.4]
  wire  valid_41_54; // @[Switch.scala 30:36:@13375.4]
  wire  _T_33604; // @[Switch.scala 30:53:@13377.4]
  wire  valid_41_55; // @[Switch.scala 30:36:@13378.4]
  wire  _T_33607; // @[Switch.scala 30:53:@13380.4]
  wire  valid_41_56; // @[Switch.scala 30:36:@13381.4]
  wire  _T_33610; // @[Switch.scala 30:53:@13383.4]
  wire  valid_41_57; // @[Switch.scala 30:36:@13384.4]
  wire  _T_33613; // @[Switch.scala 30:53:@13386.4]
  wire  valid_41_58; // @[Switch.scala 30:36:@13387.4]
  wire  _T_33616; // @[Switch.scala 30:53:@13389.4]
  wire  valid_41_59; // @[Switch.scala 30:36:@13390.4]
  wire  _T_33619; // @[Switch.scala 30:53:@13392.4]
  wire  valid_41_60; // @[Switch.scala 30:36:@13393.4]
  wire  _T_33622; // @[Switch.scala 30:53:@13395.4]
  wire  valid_41_61; // @[Switch.scala 30:36:@13396.4]
  wire  _T_33625; // @[Switch.scala 30:53:@13398.4]
  wire  valid_41_62; // @[Switch.scala 30:36:@13399.4]
  wire  _T_33628; // @[Switch.scala 30:53:@13401.4]
  wire  valid_41_63; // @[Switch.scala 30:36:@13402.4]
  wire [5:0] _T_33694; // @[Mux.scala 31:69:@13404.4]
  wire [5:0] _T_33695; // @[Mux.scala 31:69:@13405.4]
  wire [5:0] _T_33696; // @[Mux.scala 31:69:@13406.4]
  wire [5:0] _T_33697; // @[Mux.scala 31:69:@13407.4]
  wire [5:0] _T_33698; // @[Mux.scala 31:69:@13408.4]
  wire [5:0] _T_33699; // @[Mux.scala 31:69:@13409.4]
  wire [5:0] _T_33700; // @[Mux.scala 31:69:@13410.4]
  wire [5:0] _T_33701; // @[Mux.scala 31:69:@13411.4]
  wire [5:0] _T_33702; // @[Mux.scala 31:69:@13412.4]
  wire [5:0] _T_33703; // @[Mux.scala 31:69:@13413.4]
  wire [5:0] _T_33704; // @[Mux.scala 31:69:@13414.4]
  wire [5:0] _T_33705; // @[Mux.scala 31:69:@13415.4]
  wire [5:0] _T_33706; // @[Mux.scala 31:69:@13416.4]
  wire [5:0] _T_33707; // @[Mux.scala 31:69:@13417.4]
  wire [5:0] _T_33708; // @[Mux.scala 31:69:@13418.4]
  wire [5:0] _T_33709; // @[Mux.scala 31:69:@13419.4]
  wire [5:0] _T_33710; // @[Mux.scala 31:69:@13420.4]
  wire [5:0] _T_33711; // @[Mux.scala 31:69:@13421.4]
  wire [5:0] _T_33712; // @[Mux.scala 31:69:@13422.4]
  wire [5:0] _T_33713; // @[Mux.scala 31:69:@13423.4]
  wire [5:0] _T_33714; // @[Mux.scala 31:69:@13424.4]
  wire [5:0] _T_33715; // @[Mux.scala 31:69:@13425.4]
  wire [5:0] _T_33716; // @[Mux.scala 31:69:@13426.4]
  wire [5:0] _T_33717; // @[Mux.scala 31:69:@13427.4]
  wire [5:0] _T_33718; // @[Mux.scala 31:69:@13428.4]
  wire [5:0] _T_33719; // @[Mux.scala 31:69:@13429.4]
  wire [5:0] _T_33720; // @[Mux.scala 31:69:@13430.4]
  wire [5:0] _T_33721; // @[Mux.scala 31:69:@13431.4]
  wire [5:0] _T_33722; // @[Mux.scala 31:69:@13432.4]
  wire [5:0] _T_33723; // @[Mux.scala 31:69:@13433.4]
  wire [5:0] _T_33724; // @[Mux.scala 31:69:@13434.4]
  wire [5:0] _T_33725; // @[Mux.scala 31:69:@13435.4]
  wire [5:0] _T_33726; // @[Mux.scala 31:69:@13436.4]
  wire [5:0] _T_33727; // @[Mux.scala 31:69:@13437.4]
  wire [5:0] _T_33728; // @[Mux.scala 31:69:@13438.4]
  wire [5:0] _T_33729; // @[Mux.scala 31:69:@13439.4]
  wire [5:0] _T_33730; // @[Mux.scala 31:69:@13440.4]
  wire [5:0] _T_33731; // @[Mux.scala 31:69:@13441.4]
  wire [5:0] _T_33732; // @[Mux.scala 31:69:@13442.4]
  wire [5:0] _T_33733; // @[Mux.scala 31:69:@13443.4]
  wire [5:0] _T_33734; // @[Mux.scala 31:69:@13444.4]
  wire [5:0] _T_33735; // @[Mux.scala 31:69:@13445.4]
  wire [5:0] _T_33736; // @[Mux.scala 31:69:@13446.4]
  wire [5:0] _T_33737; // @[Mux.scala 31:69:@13447.4]
  wire [5:0] _T_33738; // @[Mux.scala 31:69:@13448.4]
  wire [5:0] _T_33739; // @[Mux.scala 31:69:@13449.4]
  wire [5:0] _T_33740; // @[Mux.scala 31:69:@13450.4]
  wire [5:0] _T_33741; // @[Mux.scala 31:69:@13451.4]
  wire [5:0] _T_33742; // @[Mux.scala 31:69:@13452.4]
  wire [5:0] _T_33743; // @[Mux.scala 31:69:@13453.4]
  wire [5:0] _T_33744; // @[Mux.scala 31:69:@13454.4]
  wire [5:0] _T_33745; // @[Mux.scala 31:69:@13455.4]
  wire [5:0] _T_33746; // @[Mux.scala 31:69:@13456.4]
  wire [5:0] _T_33747; // @[Mux.scala 31:69:@13457.4]
  wire [5:0] _T_33748; // @[Mux.scala 31:69:@13458.4]
  wire [5:0] _T_33749; // @[Mux.scala 31:69:@13459.4]
  wire [5:0] _T_33750; // @[Mux.scala 31:69:@13460.4]
  wire [5:0] _T_33751; // @[Mux.scala 31:69:@13461.4]
  wire [5:0] _T_33752; // @[Mux.scala 31:69:@13462.4]
  wire [5:0] _T_33753; // @[Mux.scala 31:69:@13463.4]
  wire [5:0] _T_33754; // @[Mux.scala 31:69:@13464.4]
  wire [5:0] _T_33755; // @[Mux.scala 31:69:@13465.4]
  wire [5:0] select_41; // @[Mux.scala 31:69:@13466.4]
  wire [47:0] _GEN_2625; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2626; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2627; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2628; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2629; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2630; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2631; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2632; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2633; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2634; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2635; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2636; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2637; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2638; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2639; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2640; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2641; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2642; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2643; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2644; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2645; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2646; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2647; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2648; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2649; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2650; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2651; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2652; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2653; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2654; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2655; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2656; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2657; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2658; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2659; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2660; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2661; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2662; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2663; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2664; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2665; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2666; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2667; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2668; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2669; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2670; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2671; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2672; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2673; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2674; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2675; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2676; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2677; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2678; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2679; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2680; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2681; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2682; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2683; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2684; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2685; // @[Switch.scala 33:19:@13468.4]
  wire [47:0] _GEN_2686; // @[Switch.scala 33:19:@13468.4]
  wire [7:0] _T_33764; // @[Switch.scala 34:32:@13475.4]
  wire [15:0] _T_33772; // @[Switch.scala 34:32:@13483.4]
  wire [7:0] _T_33779; // @[Switch.scala 34:32:@13490.4]
  wire [31:0] _T_33788; // @[Switch.scala 34:32:@13499.4]
  wire [7:0] _T_33795; // @[Switch.scala 34:32:@13506.4]
  wire [15:0] _T_33803; // @[Switch.scala 34:32:@13514.4]
  wire [7:0] _T_33810; // @[Switch.scala 34:32:@13521.4]
  wire [31:0] _T_33819; // @[Switch.scala 34:32:@13530.4]
  wire [63:0] _T_33820; // @[Switch.scala 34:32:@13531.4]
  wire  _T_33824; // @[Switch.scala 30:53:@13534.4]
  wire  valid_42_0; // @[Switch.scala 30:36:@13535.4]
  wire  _T_33827; // @[Switch.scala 30:53:@13537.4]
  wire  valid_42_1; // @[Switch.scala 30:36:@13538.4]
  wire  _T_33830; // @[Switch.scala 30:53:@13540.4]
  wire  valid_42_2; // @[Switch.scala 30:36:@13541.4]
  wire  _T_33833; // @[Switch.scala 30:53:@13543.4]
  wire  valid_42_3; // @[Switch.scala 30:36:@13544.4]
  wire  _T_33836; // @[Switch.scala 30:53:@13546.4]
  wire  valid_42_4; // @[Switch.scala 30:36:@13547.4]
  wire  _T_33839; // @[Switch.scala 30:53:@13549.4]
  wire  valid_42_5; // @[Switch.scala 30:36:@13550.4]
  wire  _T_33842; // @[Switch.scala 30:53:@13552.4]
  wire  valid_42_6; // @[Switch.scala 30:36:@13553.4]
  wire  _T_33845; // @[Switch.scala 30:53:@13555.4]
  wire  valid_42_7; // @[Switch.scala 30:36:@13556.4]
  wire  _T_33848; // @[Switch.scala 30:53:@13558.4]
  wire  valid_42_8; // @[Switch.scala 30:36:@13559.4]
  wire  _T_33851; // @[Switch.scala 30:53:@13561.4]
  wire  valid_42_9; // @[Switch.scala 30:36:@13562.4]
  wire  _T_33854; // @[Switch.scala 30:53:@13564.4]
  wire  valid_42_10; // @[Switch.scala 30:36:@13565.4]
  wire  _T_33857; // @[Switch.scala 30:53:@13567.4]
  wire  valid_42_11; // @[Switch.scala 30:36:@13568.4]
  wire  _T_33860; // @[Switch.scala 30:53:@13570.4]
  wire  valid_42_12; // @[Switch.scala 30:36:@13571.4]
  wire  _T_33863; // @[Switch.scala 30:53:@13573.4]
  wire  valid_42_13; // @[Switch.scala 30:36:@13574.4]
  wire  _T_33866; // @[Switch.scala 30:53:@13576.4]
  wire  valid_42_14; // @[Switch.scala 30:36:@13577.4]
  wire  _T_33869; // @[Switch.scala 30:53:@13579.4]
  wire  valid_42_15; // @[Switch.scala 30:36:@13580.4]
  wire  _T_33872; // @[Switch.scala 30:53:@13582.4]
  wire  valid_42_16; // @[Switch.scala 30:36:@13583.4]
  wire  _T_33875; // @[Switch.scala 30:53:@13585.4]
  wire  valid_42_17; // @[Switch.scala 30:36:@13586.4]
  wire  _T_33878; // @[Switch.scala 30:53:@13588.4]
  wire  valid_42_18; // @[Switch.scala 30:36:@13589.4]
  wire  _T_33881; // @[Switch.scala 30:53:@13591.4]
  wire  valid_42_19; // @[Switch.scala 30:36:@13592.4]
  wire  _T_33884; // @[Switch.scala 30:53:@13594.4]
  wire  valid_42_20; // @[Switch.scala 30:36:@13595.4]
  wire  _T_33887; // @[Switch.scala 30:53:@13597.4]
  wire  valid_42_21; // @[Switch.scala 30:36:@13598.4]
  wire  _T_33890; // @[Switch.scala 30:53:@13600.4]
  wire  valid_42_22; // @[Switch.scala 30:36:@13601.4]
  wire  _T_33893; // @[Switch.scala 30:53:@13603.4]
  wire  valid_42_23; // @[Switch.scala 30:36:@13604.4]
  wire  _T_33896; // @[Switch.scala 30:53:@13606.4]
  wire  valid_42_24; // @[Switch.scala 30:36:@13607.4]
  wire  _T_33899; // @[Switch.scala 30:53:@13609.4]
  wire  valid_42_25; // @[Switch.scala 30:36:@13610.4]
  wire  _T_33902; // @[Switch.scala 30:53:@13612.4]
  wire  valid_42_26; // @[Switch.scala 30:36:@13613.4]
  wire  _T_33905; // @[Switch.scala 30:53:@13615.4]
  wire  valid_42_27; // @[Switch.scala 30:36:@13616.4]
  wire  _T_33908; // @[Switch.scala 30:53:@13618.4]
  wire  valid_42_28; // @[Switch.scala 30:36:@13619.4]
  wire  _T_33911; // @[Switch.scala 30:53:@13621.4]
  wire  valid_42_29; // @[Switch.scala 30:36:@13622.4]
  wire  _T_33914; // @[Switch.scala 30:53:@13624.4]
  wire  valid_42_30; // @[Switch.scala 30:36:@13625.4]
  wire  _T_33917; // @[Switch.scala 30:53:@13627.4]
  wire  valid_42_31; // @[Switch.scala 30:36:@13628.4]
  wire  _T_33920; // @[Switch.scala 30:53:@13630.4]
  wire  valid_42_32; // @[Switch.scala 30:36:@13631.4]
  wire  _T_33923; // @[Switch.scala 30:53:@13633.4]
  wire  valid_42_33; // @[Switch.scala 30:36:@13634.4]
  wire  _T_33926; // @[Switch.scala 30:53:@13636.4]
  wire  valid_42_34; // @[Switch.scala 30:36:@13637.4]
  wire  _T_33929; // @[Switch.scala 30:53:@13639.4]
  wire  valid_42_35; // @[Switch.scala 30:36:@13640.4]
  wire  _T_33932; // @[Switch.scala 30:53:@13642.4]
  wire  valid_42_36; // @[Switch.scala 30:36:@13643.4]
  wire  _T_33935; // @[Switch.scala 30:53:@13645.4]
  wire  valid_42_37; // @[Switch.scala 30:36:@13646.4]
  wire  _T_33938; // @[Switch.scala 30:53:@13648.4]
  wire  valid_42_38; // @[Switch.scala 30:36:@13649.4]
  wire  _T_33941; // @[Switch.scala 30:53:@13651.4]
  wire  valid_42_39; // @[Switch.scala 30:36:@13652.4]
  wire  _T_33944; // @[Switch.scala 30:53:@13654.4]
  wire  valid_42_40; // @[Switch.scala 30:36:@13655.4]
  wire  _T_33947; // @[Switch.scala 30:53:@13657.4]
  wire  valid_42_41; // @[Switch.scala 30:36:@13658.4]
  wire  _T_33950; // @[Switch.scala 30:53:@13660.4]
  wire  valid_42_42; // @[Switch.scala 30:36:@13661.4]
  wire  _T_33953; // @[Switch.scala 30:53:@13663.4]
  wire  valid_42_43; // @[Switch.scala 30:36:@13664.4]
  wire  _T_33956; // @[Switch.scala 30:53:@13666.4]
  wire  valid_42_44; // @[Switch.scala 30:36:@13667.4]
  wire  _T_33959; // @[Switch.scala 30:53:@13669.4]
  wire  valid_42_45; // @[Switch.scala 30:36:@13670.4]
  wire  _T_33962; // @[Switch.scala 30:53:@13672.4]
  wire  valid_42_46; // @[Switch.scala 30:36:@13673.4]
  wire  _T_33965; // @[Switch.scala 30:53:@13675.4]
  wire  valid_42_47; // @[Switch.scala 30:36:@13676.4]
  wire  _T_33968; // @[Switch.scala 30:53:@13678.4]
  wire  valid_42_48; // @[Switch.scala 30:36:@13679.4]
  wire  _T_33971; // @[Switch.scala 30:53:@13681.4]
  wire  valid_42_49; // @[Switch.scala 30:36:@13682.4]
  wire  _T_33974; // @[Switch.scala 30:53:@13684.4]
  wire  valid_42_50; // @[Switch.scala 30:36:@13685.4]
  wire  _T_33977; // @[Switch.scala 30:53:@13687.4]
  wire  valid_42_51; // @[Switch.scala 30:36:@13688.4]
  wire  _T_33980; // @[Switch.scala 30:53:@13690.4]
  wire  valid_42_52; // @[Switch.scala 30:36:@13691.4]
  wire  _T_33983; // @[Switch.scala 30:53:@13693.4]
  wire  valid_42_53; // @[Switch.scala 30:36:@13694.4]
  wire  _T_33986; // @[Switch.scala 30:53:@13696.4]
  wire  valid_42_54; // @[Switch.scala 30:36:@13697.4]
  wire  _T_33989; // @[Switch.scala 30:53:@13699.4]
  wire  valid_42_55; // @[Switch.scala 30:36:@13700.4]
  wire  _T_33992; // @[Switch.scala 30:53:@13702.4]
  wire  valid_42_56; // @[Switch.scala 30:36:@13703.4]
  wire  _T_33995; // @[Switch.scala 30:53:@13705.4]
  wire  valid_42_57; // @[Switch.scala 30:36:@13706.4]
  wire  _T_33998; // @[Switch.scala 30:53:@13708.4]
  wire  valid_42_58; // @[Switch.scala 30:36:@13709.4]
  wire  _T_34001; // @[Switch.scala 30:53:@13711.4]
  wire  valid_42_59; // @[Switch.scala 30:36:@13712.4]
  wire  _T_34004; // @[Switch.scala 30:53:@13714.4]
  wire  valid_42_60; // @[Switch.scala 30:36:@13715.4]
  wire  _T_34007; // @[Switch.scala 30:53:@13717.4]
  wire  valid_42_61; // @[Switch.scala 30:36:@13718.4]
  wire  _T_34010; // @[Switch.scala 30:53:@13720.4]
  wire  valid_42_62; // @[Switch.scala 30:36:@13721.4]
  wire  _T_34013; // @[Switch.scala 30:53:@13723.4]
  wire  valid_42_63; // @[Switch.scala 30:36:@13724.4]
  wire [5:0] _T_34079; // @[Mux.scala 31:69:@13726.4]
  wire [5:0] _T_34080; // @[Mux.scala 31:69:@13727.4]
  wire [5:0] _T_34081; // @[Mux.scala 31:69:@13728.4]
  wire [5:0] _T_34082; // @[Mux.scala 31:69:@13729.4]
  wire [5:0] _T_34083; // @[Mux.scala 31:69:@13730.4]
  wire [5:0] _T_34084; // @[Mux.scala 31:69:@13731.4]
  wire [5:0] _T_34085; // @[Mux.scala 31:69:@13732.4]
  wire [5:0] _T_34086; // @[Mux.scala 31:69:@13733.4]
  wire [5:0] _T_34087; // @[Mux.scala 31:69:@13734.4]
  wire [5:0] _T_34088; // @[Mux.scala 31:69:@13735.4]
  wire [5:0] _T_34089; // @[Mux.scala 31:69:@13736.4]
  wire [5:0] _T_34090; // @[Mux.scala 31:69:@13737.4]
  wire [5:0] _T_34091; // @[Mux.scala 31:69:@13738.4]
  wire [5:0] _T_34092; // @[Mux.scala 31:69:@13739.4]
  wire [5:0] _T_34093; // @[Mux.scala 31:69:@13740.4]
  wire [5:0] _T_34094; // @[Mux.scala 31:69:@13741.4]
  wire [5:0] _T_34095; // @[Mux.scala 31:69:@13742.4]
  wire [5:0] _T_34096; // @[Mux.scala 31:69:@13743.4]
  wire [5:0] _T_34097; // @[Mux.scala 31:69:@13744.4]
  wire [5:0] _T_34098; // @[Mux.scala 31:69:@13745.4]
  wire [5:0] _T_34099; // @[Mux.scala 31:69:@13746.4]
  wire [5:0] _T_34100; // @[Mux.scala 31:69:@13747.4]
  wire [5:0] _T_34101; // @[Mux.scala 31:69:@13748.4]
  wire [5:0] _T_34102; // @[Mux.scala 31:69:@13749.4]
  wire [5:0] _T_34103; // @[Mux.scala 31:69:@13750.4]
  wire [5:0] _T_34104; // @[Mux.scala 31:69:@13751.4]
  wire [5:0] _T_34105; // @[Mux.scala 31:69:@13752.4]
  wire [5:0] _T_34106; // @[Mux.scala 31:69:@13753.4]
  wire [5:0] _T_34107; // @[Mux.scala 31:69:@13754.4]
  wire [5:0] _T_34108; // @[Mux.scala 31:69:@13755.4]
  wire [5:0] _T_34109; // @[Mux.scala 31:69:@13756.4]
  wire [5:0] _T_34110; // @[Mux.scala 31:69:@13757.4]
  wire [5:0] _T_34111; // @[Mux.scala 31:69:@13758.4]
  wire [5:0] _T_34112; // @[Mux.scala 31:69:@13759.4]
  wire [5:0] _T_34113; // @[Mux.scala 31:69:@13760.4]
  wire [5:0] _T_34114; // @[Mux.scala 31:69:@13761.4]
  wire [5:0] _T_34115; // @[Mux.scala 31:69:@13762.4]
  wire [5:0] _T_34116; // @[Mux.scala 31:69:@13763.4]
  wire [5:0] _T_34117; // @[Mux.scala 31:69:@13764.4]
  wire [5:0] _T_34118; // @[Mux.scala 31:69:@13765.4]
  wire [5:0] _T_34119; // @[Mux.scala 31:69:@13766.4]
  wire [5:0] _T_34120; // @[Mux.scala 31:69:@13767.4]
  wire [5:0] _T_34121; // @[Mux.scala 31:69:@13768.4]
  wire [5:0] _T_34122; // @[Mux.scala 31:69:@13769.4]
  wire [5:0] _T_34123; // @[Mux.scala 31:69:@13770.4]
  wire [5:0] _T_34124; // @[Mux.scala 31:69:@13771.4]
  wire [5:0] _T_34125; // @[Mux.scala 31:69:@13772.4]
  wire [5:0] _T_34126; // @[Mux.scala 31:69:@13773.4]
  wire [5:0] _T_34127; // @[Mux.scala 31:69:@13774.4]
  wire [5:0] _T_34128; // @[Mux.scala 31:69:@13775.4]
  wire [5:0] _T_34129; // @[Mux.scala 31:69:@13776.4]
  wire [5:0] _T_34130; // @[Mux.scala 31:69:@13777.4]
  wire [5:0] _T_34131; // @[Mux.scala 31:69:@13778.4]
  wire [5:0] _T_34132; // @[Mux.scala 31:69:@13779.4]
  wire [5:0] _T_34133; // @[Mux.scala 31:69:@13780.4]
  wire [5:0] _T_34134; // @[Mux.scala 31:69:@13781.4]
  wire [5:0] _T_34135; // @[Mux.scala 31:69:@13782.4]
  wire [5:0] _T_34136; // @[Mux.scala 31:69:@13783.4]
  wire [5:0] _T_34137; // @[Mux.scala 31:69:@13784.4]
  wire [5:0] _T_34138; // @[Mux.scala 31:69:@13785.4]
  wire [5:0] _T_34139; // @[Mux.scala 31:69:@13786.4]
  wire [5:0] _T_34140; // @[Mux.scala 31:69:@13787.4]
  wire [5:0] select_42; // @[Mux.scala 31:69:@13788.4]
  wire [47:0] _GEN_2689; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2690; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2691; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2692; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2693; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2694; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2695; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2696; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2697; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2698; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2699; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2700; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2701; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2702; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2703; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2704; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2705; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2706; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2707; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2708; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2709; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2710; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2711; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2712; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2713; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2714; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2715; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2716; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2717; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2718; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2719; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2720; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2721; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2722; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2723; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2724; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2725; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2726; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2727; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2728; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2729; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2730; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2731; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2732; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2733; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2734; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2735; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2736; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2737; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2738; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2739; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2740; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2741; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2742; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2743; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2744; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2745; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2746; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2747; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2748; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2749; // @[Switch.scala 33:19:@13790.4]
  wire [47:0] _GEN_2750; // @[Switch.scala 33:19:@13790.4]
  wire [7:0] _T_34149; // @[Switch.scala 34:32:@13797.4]
  wire [15:0] _T_34157; // @[Switch.scala 34:32:@13805.4]
  wire [7:0] _T_34164; // @[Switch.scala 34:32:@13812.4]
  wire [31:0] _T_34173; // @[Switch.scala 34:32:@13821.4]
  wire [7:0] _T_34180; // @[Switch.scala 34:32:@13828.4]
  wire [15:0] _T_34188; // @[Switch.scala 34:32:@13836.4]
  wire [7:0] _T_34195; // @[Switch.scala 34:32:@13843.4]
  wire [31:0] _T_34204; // @[Switch.scala 34:32:@13852.4]
  wire [63:0] _T_34205; // @[Switch.scala 34:32:@13853.4]
  wire  _T_34209; // @[Switch.scala 30:53:@13856.4]
  wire  valid_43_0; // @[Switch.scala 30:36:@13857.4]
  wire  _T_34212; // @[Switch.scala 30:53:@13859.4]
  wire  valid_43_1; // @[Switch.scala 30:36:@13860.4]
  wire  _T_34215; // @[Switch.scala 30:53:@13862.4]
  wire  valid_43_2; // @[Switch.scala 30:36:@13863.4]
  wire  _T_34218; // @[Switch.scala 30:53:@13865.4]
  wire  valid_43_3; // @[Switch.scala 30:36:@13866.4]
  wire  _T_34221; // @[Switch.scala 30:53:@13868.4]
  wire  valid_43_4; // @[Switch.scala 30:36:@13869.4]
  wire  _T_34224; // @[Switch.scala 30:53:@13871.4]
  wire  valid_43_5; // @[Switch.scala 30:36:@13872.4]
  wire  _T_34227; // @[Switch.scala 30:53:@13874.4]
  wire  valid_43_6; // @[Switch.scala 30:36:@13875.4]
  wire  _T_34230; // @[Switch.scala 30:53:@13877.4]
  wire  valid_43_7; // @[Switch.scala 30:36:@13878.4]
  wire  _T_34233; // @[Switch.scala 30:53:@13880.4]
  wire  valid_43_8; // @[Switch.scala 30:36:@13881.4]
  wire  _T_34236; // @[Switch.scala 30:53:@13883.4]
  wire  valid_43_9; // @[Switch.scala 30:36:@13884.4]
  wire  _T_34239; // @[Switch.scala 30:53:@13886.4]
  wire  valid_43_10; // @[Switch.scala 30:36:@13887.4]
  wire  _T_34242; // @[Switch.scala 30:53:@13889.4]
  wire  valid_43_11; // @[Switch.scala 30:36:@13890.4]
  wire  _T_34245; // @[Switch.scala 30:53:@13892.4]
  wire  valid_43_12; // @[Switch.scala 30:36:@13893.4]
  wire  _T_34248; // @[Switch.scala 30:53:@13895.4]
  wire  valid_43_13; // @[Switch.scala 30:36:@13896.4]
  wire  _T_34251; // @[Switch.scala 30:53:@13898.4]
  wire  valid_43_14; // @[Switch.scala 30:36:@13899.4]
  wire  _T_34254; // @[Switch.scala 30:53:@13901.4]
  wire  valid_43_15; // @[Switch.scala 30:36:@13902.4]
  wire  _T_34257; // @[Switch.scala 30:53:@13904.4]
  wire  valid_43_16; // @[Switch.scala 30:36:@13905.4]
  wire  _T_34260; // @[Switch.scala 30:53:@13907.4]
  wire  valid_43_17; // @[Switch.scala 30:36:@13908.4]
  wire  _T_34263; // @[Switch.scala 30:53:@13910.4]
  wire  valid_43_18; // @[Switch.scala 30:36:@13911.4]
  wire  _T_34266; // @[Switch.scala 30:53:@13913.4]
  wire  valid_43_19; // @[Switch.scala 30:36:@13914.4]
  wire  _T_34269; // @[Switch.scala 30:53:@13916.4]
  wire  valid_43_20; // @[Switch.scala 30:36:@13917.4]
  wire  _T_34272; // @[Switch.scala 30:53:@13919.4]
  wire  valid_43_21; // @[Switch.scala 30:36:@13920.4]
  wire  _T_34275; // @[Switch.scala 30:53:@13922.4]
  wire  valid_43_22; // @[Switch.scala 30:36:@13923.4]
  wire  _T_34278; // @[Switch.scala 30:53:@13925.4]
  wire  valid_43_23; // @[Switch.scala 30:36:@13926.4]
  wire  _T_34281; // @[Switch.scala 30:53:@13928.4]
  wire  valid_43_24; // @[Switch.scala 30:36:@13929.4]
  wire  _T_34284; // @[Switch.scala 30:53:@13931.4]
  wire  valid_43_25; // @[Switch.scala 30:36:@13932.4]
  wire  _T_34287; // @[Switch.scala 30:53:@13934.4]
  wire  valid_43_26; // @[Switch.scala 30:36:@13935.4]
  wire  _T_34290; // @[Switch.scala 30:53:@13937.4]
  wire  valid_43_27; // @[Switch.scala 30:36:@13938.4]
  wire  _T_34293; // @[Switch.scala 30:53:@13940.4]
  wire  valid_43_28; // @[Switch.scala 30:36:@13941.4]
  wire  _T_34296; // @[Switch.scala 30:53:@13943.4]
  wire  valid_43_29; // @[Switch.scala 30:36:@13944.4]
  wire  _T_34299; // @[Switch.scala 30:53:@13946.4]
  wire  valid_43_30; // @[Switch.scala 30:36:@13947.4]
  wire  _T_34302; // @[Switch.scala 30:53:@13949.4]
  wire  valid_43_31; // @[Switch.scala 30:36:@13950.4]
  wire  _T_34305; // @[Switch.scala 30:53:@13952.4]
  wire  valid_43_32; // @[Switch.scala 30:36:@13953.4]
  wire  _T_34308; // @[Switch.scala 30:53:@13955.4]
  wire  valid_43_33; // @[Switch.scala 30:36:@13956.4]
  wire  _T_34311; // @[Switch.scala 30:53:@13958.4]
  wire  valid_43_34; // @[Switch.scala 30:36:@13959.4]
  wire  _T_34314; // @[Switch.scala 30:53:@13961.4]
  wire  valid_43_35; // @[Switch.scala 30:36:@13962.4]
  wire  _T_34317; // @[Switch.scala 30:53:@13964.4]
  wire  valid_43_36; // @[Switch.scala 30:36:@13965.4]
  wire  _T_34320; // @[Switch.scala 30:53:@13967.4]
  wire  valid_43_37; // @[Switch.scala 30:36:@13968.4]
  wire  _T_34323; // @[Switch.scala 30:53:@13970.4]
  wire  valid_43_38; // @[Switch.scala 30:36:@13971.4]
  wire  _T_34326; // @[Switch.scala 30:53:@13973.4]
  wire  valid_43_39; // @[Switch.scala 30:36:@13974.4]
  wire  _T_34329; // @[Switch.scala 30:53:@13976.4]
  wire  valid_43_40; // @[Switch.scala 30:36:@13977.4]
  wire  _T_34332; // @[Switch.scala 30:53:@13979.4]
  wire  valid_43_41; // @[Switch.scala 30:36:@13980.4]
  wire  _T_34335; // @[Switch.scala 30:53:@13982.4]
  wire  valid_43_42; // @[Switch.scala 30:36:@13983.4]
  wire  _T_34338; // @[Switch.scala 30:53:@13985.4]
  wire  valid_43_43; // @[Switch.scala 30:36:@13986.4]
  wire  _T_34341; // @[Switch.scala 30:53:@13988.4]
  wire  valid_43_44; // @[Switch.scala 30:36:@13989.4]
  wire  _T_34344; // @[Switch.scala 30:53:@13991.4]
  wire  valid_43_45; // @[Switch.scala 30:36:@13992.4]
  wire  _T_34347; // @[Switch.scala 30:53:@13994.4]
  wire  valid_43_46; // @[Switch.scala 30:36:@13995.4]
  wire  _T_34350; // @[Switch.scala 30:53:@13997.4]
  wire  valid_43_47; // @[Switch.scala 30:36:@13998.4]
  wire  _T_34353; // @[Switch.scala 30:53:@14000.4]
  wire  valid_43_48; // @[Switch.scala 30:36:@14001.4]
  wire  _T_34356; // @[Switch.scala 30:53:@14003.4]
  wire  valid_43_49; // @[Switch.scala 30:36:@14004.4]
  wire  _T_34359; // @[Switch.scala 30:53:@14006.4]
  wire  valid_43_50; // @[Switch.scala 30:36:@14007.4]
  wire  _T_34362; // @[Switch.scala 30:53:@14009.4]
  wire  valid_43_51; // @[Switch.scala 30:36:@14010.4]
  wire  _T_34365; // @[Switch.scala 30:53:@14012.4]
  wire  valid_43_52; // @[Switch.scala 30:36:@14013.4]
  wire  _T_34368; // @[Switch.scala 30:53:@14015.4]
  wire  valid_43_53; // @[Switch.scala 30:36:@14016.4]
  wire  _T_34371; // @[Switch.scala 30:53:@14018.4]
  wire  valid_43_54; // @[Switch.scala 30:36:@14019.4]
  wire  _T_34374; // @[Switch.scala 30:53:@14021.4]
  wire  valid_43_55; // @[Switch.scala 30:36:@14022.4]
  wire  _T_34377; // @[Switch.scala 30:53:@14024.4]
  wire  valid_43_56; // @[Switch.scala 30:36:@14025.4]
  wire  _T_34380; // @[Switch.scala 30:53:@14027.4]
  wire  valid_43_57; // @[Switch.scala 30:36:@14028.4]
  wire  _T_34383; // @[Switch.scala 30:53:@14030.4]
  wire  valid_43_58; // @[Switch.scala 30:36:@14031.4]
  wire  _T_34386; // @[Switch.scala 30:53:@14033.4]
  wire  valid_43_59; // @[Switch.scala 30:36:@14034.4]
  wire  _T_34389; // @[Switch.scala 30:53:@14036.4]
  wire  valid_43_60; // @[Switch.scala 30:36:@14037.4]
  wire  _T_34392; // @[Switch.scala 30:53:@14039.4]
  wire  valid_43_61; // @[Switch.scala 30:36:@14040.4]
  wire  _T_34395; // @[Switch.scala 30:53:@14042.4]
  wire  valid_43_62; // @[Switch.scala 30:36:@14043.4]
  wire  _T_34398; // @[Switch.scala 30:53:@14045.4]
  wire  valid_43_63; // @[Switch.scala 30:36:@14046.4]
  wire [5:0] _T_34464; // @[Mux.scala 31:69:@14048.4]
  wire [5:0] _T_34465; // @[Mux.scala 31:69:@14049.4]
  wire [5:0] _T_34466; // @[Mux.scala 31:69:@14050.4]
  wire [5:0] _T_34467; // @[Mux.scala 31:69:@14051.4]
  wire [5:0] _T_34468; // @[Mux.scala 31:69:@14052.4]
  wire [5:0] _T_34469; // @[Mux.scala 31:69:@14053.4]
  wire [5:0] _T_34470; // @[Mux.scala 31:69:@14054.4]
  wire [5:0] _T_34471; // @[Mux.scala 31:69:@14055.4]
  wire [5:0] _T_34472; // @[Mux.scala 31:69:@14056.4]
  wire [5:0] _T_34473; // @[Mux.scala 31:69:@14057.4]
  wire [5:0] _T_34474; // @[Mux.scala 31:69:@14058.4]
  wire [5:0] _T_34475; // @[Mux.scala 31:69:@14059.4]
  wire [5:0] _T_34476; // @[Mux.scala 31:69:@14060.4]
  wire [5:0] _T_34477; // @[Mux.scala 31:69:@14061.4]
  wire [5:0] _T_34478; // @[Mux.scala 31:69:@14062.4]
  wire [5:0] _T_34479; // @[Mux.scala 31:69:@14063.4]
  wire [5:0] _T_34480; // @[Mux.scala 31:69:@14064.4]
  wire [5:0] _T_34481; // @[Mux.scala 31:69:@14065.4]
  wire [5:0] _T_34482; // @[Mux.scala 31:69:@14066.4]
  wire [5:0] _T_34483; // @[Mux.scala 31:69:@14067.4]
  wire [5:0] _T_34484; // @[Mux.scala 31:69:@14068.4]
  wire [5:0] _T_34485; // @[Mux.scala 31:69:@14069.4]
  wire [5:0] _T_34486; // @[Mux.scala 31:69:@14070.4]
  wire [5:0] _T_34487; // @[Mux.scala 31:69:@14071.4]
  wire [5:0] _T_34488; // @[Mux.scala 31:69:@14072.4]
  wire [5:0] _T_34489; // @[Mux.scala 31:69:@14073.4]
  wire [5:0] _T_34490; // @[Mux.scala 31:69:@14074.4]
  wire [5:0] _T_34491; // @[Mux.scala 31:69:@14075.4]
  wire [5:0] _T_34492; // @[Mux.scala 31:69:@14076.4]
  wire [5:0] _T_34493; // @[Mux.scala 31:69:@14077.4]
  wire [5:0] _T_34494; // @[Mux.scala 31:69:@14078.4]
  wire [5:0] _T_34495; // @[Mux.scala 31:69:@14079.4]
  wire [5:0] _T_34496; // @[Mux.scala 31:69:@14080.4]
  wire [5:0] _T_34497; // @[Mux.scala 31:69:@14081.4]
  wire [5:0] _T_34498; // @[Mux.scala 31:69:@14082.4]
  wire [5:0] _T_34499; // @[Mux.scala 31:69:@14083.4]
  wire [5:0] _T_34500; // @[Mux.scala 31:69:@14084.4]
  wire [5:0] _T_34501; // @[Mux.scala 31:69:@14085.4]
  wire [5:0] _T_34502; // @[Mux.scala 31:69:@14086.4]
  wire [5:0] _T_34503; // @[Mux.scala 31:69:@14087.4]
  wire [5:0] _T_34504; // @[Mux.scala 31:69:@14088.4]
  wire [5:0] _T_34505; // @[Mux.scala 31:69:@14089.4]
  wire [5:0] _T_34506; // @[Mux.scala 31:69:@14090.4]
  wire [5:0] _T_34507; // @[Mux.scala 31:69:@14091.4]
  wire [5:0] _T_34508; // @[Mux.scala 31:69:@14092.4]
  wire [5:0] _T_34509; // @[Mux.scala 31:69:@14093.4]
  wire [5:0] _T_34510; // @[Mux.scala 31:69:@14094.4]
  wire [5:0] _T_34511; // @[Mux.scala 31:69:@14095.4]
  wire [5:0] _T_34512; // @[Mux.scala 31:69:@14096.4]
  wire [5:0] _T_34513; // @[Mux.scala 31:69:@14097.4]
  wire [5:0] _T_34514; // @[Mux.scala 31:69:@14098.4]
  wire [5:0] _T_34515; // @[Mux.scala 31:69:@14099.4]
  wire [5:0] _T_34516; // @[Mux.scala 31:69:@14100.4]
  wire [5:0] _T_34517; // @[Mux.scala 31:69:@14101.4]
  wire [5:0] _T_34518; // @[Mux.scala 31:69:@14102.4]
  wire [5:0] _T_34519; // @[Mux.scala 31:69:@14103.4]
  wire [5:0] _T_34520; // @[Mux.scala 31:69:@14104.4]
  wire [5:0] _T_34521; // @[Mux.scala 31:69:@14105.4]
  wire [5:0] _T_34522; // @[Mux.scala 31:69:@14106.4]
  wire [5:0] _T_34523; // @[Mux.scala 31:69:@14107.4]
  wire [5:0] _T_34524; // @[Mux.scala 31:69:@14108.4]
  wire [5:0] _T_34525; // @[Mux.scala 31:69:@14109.4]
  wire [5:0] select_43; // @[Mux.scala 31:69:@14110.4]
  wire [47:0] _GEN_2753; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2754; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2755; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2756; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2757; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2758; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2759; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2760; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2761; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2762; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2763; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2764; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2765; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2766; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2767; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2768; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2769; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2770; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2771; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2772; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2773; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2774; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2775; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2776; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2777; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2778; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2779; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2780; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2781; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2782; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2783; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2784; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2785; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2786; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2787; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2788; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2789; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2790; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2791; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2792; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2793; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2794; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2795; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2796; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2797; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2798; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2799; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2800; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2801; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2802; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2803; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2804; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2805; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2806; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2807; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2808; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2809; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2810; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2811; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2812; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2813; // @[Switch.scala 33:19:@14112.4]
  wire [47:0] _GEN_2814; // @[Switch.scala 33:19:@14112.4]
  wire [7:0] _T_34534; // @[Switch.scala 34:32:@14119.4]
  wire [15:0] _T_34542; // @[Switch.scala 34:32:@14127.4]
  wire [7:0] _T_34549; // @[Switch.scala 34:32:@14134.4]
  wire [31:0] _T_34558; // @[Switch.scala 34:32:@14143.4]
  wire [7:0] _T_34565; // @[Switch.scala 34:32:@14150.4]
  wire [15:0] _T_34573; // @[Switch.scala 34:32:@14158.4]
  wire [7:0] _T_34580; // @[Switch.scala 34:32:@14165.4]
  wire [31:0] _T_34589; // @[Switch.scala 34:32:@14174.4]
  wire [63:0] _T_34590; // @[Switch.scala 34:32:@14175.4]
  wire  _T_34594; // @[Switch.scala 30:53:@14178.4]
  wire  valid_44_0; // @[Switch.scala 30:36:@14179.4]
  wire  _T_34597; // @[Switch.scala 30:53:@14181.4]
  wire  valid_44_1; // @[Switch.scala 30:36:@14182.4]
  wire  _T_34600; // @[Switch.scala 30:53:@14184.4]
  wire  valid_44_2; // @[Switch.scala 30:36:@14185.4]
  wire  _T_34603; // @[Switch.scala 30:53:@14187.4]
  wire  valid_44_3; // @[Switch.scala 30:36:@14188.4]
  wire  _T_34606; // @[Switch.scala 30:53:@14190.4]
  wire  valid_44_4; // @[Switch.scala 30:36:@14191.4]
  wire  _T_34609; // @[Switch.scala 30:53:@14193.4]
  wire  valid_44_5; // @[Switch.scala 30:36:@14194.4]
  wire  _T_34612; // @[Switch.scala 30:53:@14196.4]
  wire  valid_44_6; // @[Switch.scala 30:36:@14197.4]
  wire  _T_34615; // @[Switch.scala 30:53:@14199.4]
  wire  valid_44_7; // @[Switch.scala 30:36:@14200.4]
  wire  _T_34618; // @[Switch.scala 30:53:@14202.4]
  wire  valid_44_8; // @[Switch.scala 30:36:@14203.4]
  wire  _T_34621; // @[Switch.scala 30:53:@14205.4]
  wire  valid_44_9; // @[Switch.scala 30:36:@14206.4]
  wire  _T_34624; // @[Switch.scala 30:53:@14208.4]
  wire  valid_44_10; // @[Switch.scala 30:36:@14209.4]
  wire  _T_34627; // @[Switch.scala 30:53:@14211.4]
  wire  valid_44_11; // @[Switch.scala 30:36:@14212.4]
  wire  _T_34630; // @[Switch.scala 30:53:@14214.4]
  wire  valid_44_12; // @[Switch.scala 30:36:@14215.4]
  wire  _T_34633; // @[Switch.scala 30:53:@14217.4]
  wire  valid_44_13; // @[Switch.scala 30:36:@14218.4]
  wire  _T_34636; // @[Switch.scala 30:53:@14220.4]
  wire  valid_44_14; // @[Switch.scala 30:36:@14221.4]
  wire  _T_34639; // @[Switch.scala 30:53:@14223.4]
  wire  valid_44_15; // @[Switch.scala 30:36:@14224.4]
  wire  _T_34642; // @[Switch.scala 30:53:@14226.4]
  wire  valid_44_16; // @[Switch.scala 30:36:@14227.4]
  wire  _T_34645; // @[Switch.scala 30:53:@14229.4]
  wire  valid_44_17; // @[Switch.scala 30:36:@14230.4]
  wire  _T_34648; // @[Switch.scala 30:53:@14232.4]
  wire  valid_44_18; // @[Switch.scala 30:36:@14233.4]
  wire  _T_34651; // @[Switch.scala 30:53:@14235.4]
  wire  valid_44_19; // @[Switch.scala 30:36:@14236.4]
  wire  _T_34654; // @[Switch.scala 30:53:@14238.4]
  wire  valid_44_20; // @[Switch.scala 30:36:@14239.4]
  wire  _T_34657; // @[Switch.scala 30:53:@14241.4]
  wire  valid_44_21; // @[Switch.scala 30:36:@14242.4]
  wire  _T_34660; // @[Switch.scala 30:53:@14244.4]
  wire  valid_44_22; // @[Switch.scala 30:36:@14245.4]
  wire  _T_34663; // @[Switch.scala 30:53:@14247.4]
  wire  valid_44_23; // @[Switch.scala 30:36:@14248.4]
  wire  _T_34666; // @[Switch.scala 30:53:@14250.4]
  wire  valid_44_24; // @[Switch.scala 30:36:@14251.4]
  wire  _T_34669; // @[Switch.scala 30:53:@14253.4]
  wire  valid_44_25; // @[Switch.scala 30:36:@14254.4]
  wire  _T_34672; // @[Switch.scala 30:53:@14256.4]
  wire  valid_44_26; // @[Switch.scala 30:36:@14257.4]
  wire  _T_34675; // @[Switch.scala 30:53:@14259.4]
  wire  valid_44_27; // @[Switch.scala 30:36:@14260.4]
  wire  _T_34678; // @[Switch.scala 30:53:@14262.4]
  wire  valid_44_28; // @[Switch.scala 30:36:@14263.4]
  wire  _T_34681; // @[Switch.scala 30:53:@14265.4]
  wire  valid_44_29; // @[Switch.scala 30:36:@14266.4]
  wire  _T_34684; // @[Switch.scala 30:53:@14268.4]
  wire  valid_44_30; // @[Switch.scala 30:36:@14269.4]
  wire  _T_34687; // @[Switch.scala 30:53:@14271.4]
  wire  valid_44_31; // @[Switch.scala 30:36:@14272.4]
  wire  _T_34690; // @[Switch.scala 30:53:@14274.4]
  wire  valid_44_32; // @[Switch.scala 30:36:@14275.4]
  wire  _T_34693; // @[Switch.scala 30:53:@14277.4]
  wire  valid_44_33; // @[Switch.scala 30:36:@14278.4]
  wire  _T_34696; // @[Switch.scala 30:53:@14280.4]
  wire  valid_44_34; // @[Switch.scala 30:36:@14281.4]
  wire  _T_34699; // @[Switch.scala 30:53:@14283.4]
  wire  valid_44_35; // @[Switch.scala 30:36:@14284.4]
  wire  _T_34702; // @[Switch.scala 30:53:@14286.4]
  wire  valid_44_36; // @[Switch.scala 30:36:@14287.4]
  wire  _T_34705; // @[Switch.scala 30:53:@14289.4]
  wire  valid_44_37; // @[Switch.scala 30:36:@14290.4]
  wire  _T_34708; // @[Switch.scala 30:53:@14292.4]
  wire  valid_44_38; // @[Switch.scala 30:36:@14293.4]
  wire  _T_34711; // @[Switch.scala 30:53:@14295.4]
  wire  valid_44_39; // @[Switch.scala 30:36:@14296.4]
  wire  _T_34714; // @[Switch.scala 30:53:@14298.4]
  wire  valid_44_40; // @[Switch.scala 30:36:@14299.4]
  wire  _T_34717; // @[Switch.scala 30:53:@14301.4]
  wire  valid_44_41; // @[Switch.scala 30:36:@14302.4]
  wire  _T_34720; // @[Switch.scala 30:53:@14304.4]
  wire  valid_44_42; // @[Switch.scala 30:36:@14305.4]
  wire  _T_34723; // @[Switch.scala 30:53:@14307.4]
  wire  valid_44_43; // @[Switch.scala 30:36:@14308.4]
  wire  _T_34726; // @[Switch.scala 30:53:@14310.4]
  wire  valid_44_44; // @[Switch.scala 30:36:@14311.4]
  wire  _T_34729; // @[Switch.scala 30:53:@14313.4]
  wire  valid_44_45; // @[Switch.scala 30:36:@14314.4]
  wire  _T_34732; // @[Switch.scala 30:53:@14316.4]
  wire  valid_44_46; // @[Switch.scala 30:36:@14317.4]
  wire  _T_34735; // @[Switch.scala 30:53:@14319.4]
  wire  valid_44_47; // @[Switch.scala 30:36:@14320.4]
  wire  _T_34738; // @[Switch.scala 30:53:@14322.4]
  wire  valid_44_48; // @[Switch.scala 30:36:@14323.4]
  wire  _T_34741; // @[Switch.scala 30:53:@14325.4]
  wire  valid_44_49; // @[Switch.scala 30:36:@14326.4]
  wire  _T_34744; // @[Switch.scala 30:53:@14328.4]
  wire  valid_44_50; // @[Switch.scala 30:36:@14329.4]
  wire  _T_34747; // @[Switch.scala 30:53:@14331.4]
  wire  valid_44_51; // @[Switch.scala 30:36:@14332.4]
  wire  _T_34750; // @[Switch.scala 30:53:@14334.4]
  wire  valid_44_52; // @[Switch.scala 30:36:@14335.4]
  wire  _T_34753; // @[Switch.scala 30:53:@14337.4]
  wire  valid_44_53; // @[Switch.scala 30:36:@14338.4]
  wire  _T_34756; // @[Switch.scala 30:53:@14340.4]
  wire  valid_44_54; // @[Switch.scala 30:36:@14341.4]
  wire  _T_34759; // @[Switch.scala 30:53:@14343.4]
  wire  valid_44_55; // @[Switch.scala 30:36:@14344.4]
  wire  _T_34762; // @[Switch.scala 30:53:@14346.4]
  wire  valid_44_56; // @[Switch.scala 30:36:@14347.4]
  wire  _T_34765; // @[Switch.scala 30:53:@14349.4]
  wire  valid_44_57; // @[Switch.scala 30:36:@14350.4]
  wire  _T_34768; // @[Switch.scala 30:53:@14352.4]
  wire  valid_44_58; // @[Switch.scala 30:36:@14353.4]
  wire  _T_34771; // @[Switch.scala 30:53:@14355.4]
  wire  valid_44_59; // @[Switch.scala 30:36:@14356.4]
  wire  _T_34774; // @[Switch.scala 30:53:@14358.4]
  wire  valid_44_60; // @[Switch.scala 30:36:@14359.4]
  wire  _T_34777; // @[Switch.scala 30:53:@14361.4]
  wire  valid_44_61; // @[Switch.scala 30:36:@14362.4]
  wire  _T_34780; // @[Switch.scala 30:53:@14364.4]
  wire  valid_44_62; // @[Switch.scala 30:36:@14365.4]
  wire  _T_34783; // @[Switch.scala 30:53:@14367.4]
  wire  valid_44_63; // @[Switch.scala 30:36:@14368.4]
  wire [5:0] _T_34849; // @[Mux.scala 31:69:@14370.4]
  wire [5:0] _T_34850; // @[Mux.scala 31:69:@14371.4]
  wire [5:0] _T_34851; // @[Mux.scala 31:69:@14372.4]
  wire [5:0] _T_34852; // @[Mux.scala 31:69:@14373.4]
  wire [5:0] _T_34853; // @[Mux.scala 31:69:@14374.4]
  wire [5:0] _T_34854; // @[Mux.scala 31:69:@14375.4]
  wire [5:0] _T_34855; // @[Mux.scala 31:69:@14376.4]
  wire [5:0] _T_34856; // @[Mux.scala 31:69:@14377.4]
  wire [5:0] _T_34857; // @[Mux.scala 31:69:@14378.4]
  wire [5:0] _T_34858; // @[Mux.scala 31:69:@14379.4]
  wire [5:0] _T_34859; // @[Mux.scala 31:69:@14380.4]
  wire [5:0] _T_34860; // @[Mux.scala 31:69:@14381.4]
  wire [5:0] _T_34861; // @[Mux.scala 31:69:@14382.4]
  wire [5:0] _T_34862; // @[Mux.scala 31:69:@14383.4]
  wire [5:0] _T_34863; // @[Mux.scala 31:69:@14384.4]
  wire [5:0] _T_34864; // @[Mux.scala 31:69:@14385.4]
  wire [5:0] _T_34865; // @[Mux.scala 31:69:@14386.4]
  wire [5:0] _T_34866; // @[Mux.scala 31:69:@14387.4]
  wire [5:0] _T_34867; // @[Mux.scala 31:69:@14388.4]
  wire [5:0] _T_34868; // @[Mux.scala 31:69:@14389.4]
  wire [5:0] _T_34869; // @[Mux.scala 31:69:@14390.4]
  wire [5:0] _T_34870; // @[Mux.scala 31:69:@14391.4]
  wire [5:0] _T_34871; // @[Mux.scala 31:69:@14392.4]
  wire [5:0] _T_34872; // @[Mux.scala 31:69:@14393.4]
  wire [5:0] _T_34873; // @[Mux.scala 31:69:@14394.4]
  wire [5:0] _T_34874; // @[Mux.scala 31:69:@14395.4]
  wire [5:0] _T_34875; // @[Mux.scala 31:69:@14396.4]
  wire [5:0] _T_34876; // @[Mux.scala 31:69:@14397.4]
  wire [5:0] _T_34877; // @[Mux.scala 31:69:@14398.4]
  wire [5:0] _T_34878; // @[Mux.scala 31:69:@14399.4]
  wire [5:0] _T_34879; // @[Mux.scala 31:69:@14400.4]
  wire [5:0] _T_34880; // @[Mux.scala 31:69:@14401.4]
  wire [5:0] _T_34881; // @[Mux.scala 31:69:@14402.4]
  wire [5:0] _T_34882; // @[Mux.scala 31:69:@14403.4]
  wire [5:0] _T_34883; // @[Mux.scala 31:69:@14404.4]
  wire [5:0] _T_34884; // @[Mux.scala 31:69:@14405.4]
  wire [5:0] _T_34885; // @[Mux.scala 31:69:@14406.4]
  wire [5:0] _T_34886; // @[Mux.scala 31:69:@14407.4]
  wire [5:0] _T_34887; // @[Mux.scala 31:69:@14408.4]
  wire [5:0] _T_34888; // @[Mux.scala 31:69:@14409.4]
  wire [5:0] _T_34889; // @[Mux.scala 31:69:@14410.4]
  wire [5:0] _T_34890; // @[Mux.scala 31:69:@14411.4]
  wire [5:0] _T_34891; // @[Mux.scala 31:69:@14412.4]
  wire [5:0] _T_34892; // @[Mux.scala 31:69:@14413.4]
  wire [5:0] _T_34893; // @[Mux.scala 31:69:@14414.4]
  wire [5:0] _T_34894; // @[Mux.scala 31:69:@14415.4]
  wire [5:0] _T_34895; // @[Mux.scala 31:69:@14416.4]
  wire [5:0] _T_34896; // @[Mux.scala 31:69:@14417.4]
  wire [5:0] _T_34897; // @[Mux.scala 31:69:@14418.4]
  wire [5:0] _T_34898; // @[Mux.scala 31:69:@14419.4]
  wire [5:0] _T_34899; // @[Mux.scala 31:69:@14420.4]
  wire [5:0] _T_34900; // @[Mux.scala 31:69:@14421.4]
  wire [5:0] _T_34901; // @[Mux.scala 31:69:@14422.4]
  wire [5:0] _T_34902; // @[Mux.scala 31:69:@14423.4]
  wire [5:0] _T_34903; // @[Mux.scala 31:69:@14424.4]
  wire [5:0] _T_34904; // @[Mux.scala 31:69:@14425.4]
  wire [5:0] _T_34905; // @[Mux.scala 31:69:@14426.4]
  wire [5:0] _T_34906; // @[Mux.scala 31:69:@14427.4]
  wire [5:0] _T_34907; // @[Mux.scala 31:69:@14428.4]
  wire [5:0] _T_34908; // @[Mux.scala 31:69:@14429.4]
  wire [5:0] _T_34909; // @[Mux.scala 31:69:@14430.4]
  wire [5:0] _T_34910; // @[Mux.scala 31:69:@14431.4]
  wire [5:0] select_44; // @[Mux.scala 31:69:@14432.4]
  wire [47:0] _GEN_2817; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2818; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2819; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2820; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2821; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2822; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2823; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2824; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2825; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2826; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2827; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2828; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2829; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2830; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2831; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2832; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2833; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2834; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2835; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2836; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2837; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2838; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2839; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2840; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2841; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2842; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2843; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2844; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2845; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2846; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2847; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2848; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2849; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2850; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2851; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2852; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2853; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2854; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2855; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2856; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2857; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2858; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2859; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2860; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2861; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2862; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2863; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2864; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2865; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2866; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2867; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2868; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2869; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2870; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2871; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2872; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2873; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2874; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2875; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2876; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2877; // @[Switch.scala 33:19:@14434.4]
  wire [47:0] _GEN_2878; // @[Switch.scala 33:19:@14434.4]
  wire [7:0] _T_34919; // @[Switch.scala 34:32:@14441.4]
  wire [15:0] _T_34927; // @[Switch.scala 34:32:@14449.4]
  wire [7:0] _T_34934; // @[Switch.scala 34:32:@14456.4]
  wire [31:0] _T_34943; // @[Switch.scala 34:32:@14465.4]
  wire [7:0] _T_34950; // @[Switch.scala 34:32:@14472.4]
  wire [15:0] _T_34958; // @[Switch.scala 34:32:@14480.4]
  wire [7:0] _T_34965; // @[Switch.scala 34:32:@14487.4]
  wire [31:0] _T_34974; // @[Switch.scala 34:32:@14496.4]
  wire [63:0] _T_34975; // @[Switch.scala 34:32:@14497.4]
  wire  _T_34979; // @[Switch.scala 30:53:@14500.4]
  wire  valid_45_0; // @[Switch.scala 30:36:@14501.4]
  wire  _T_34982; // @[Switch.scala 30:53:@14503.4]
  wire  valid_45_1; // @[Switch.scala 30:36:@14504.4]
  wire  _T_34985; // @[Switch.scala 30:53:@14506.4]
  wire  valid_45_2; // @[Switch.scala 30:36:@14507.4]
  wire  _T_34988; // @[Switch.scala 30:53:@14509.4]
  wire  valid_45_3; // @[Switch.scala 30:36:@14510.4]
  wire  _T_34991; // @[Switch.scala 30:53:@14512.4]
  wire  valid_45_4; // @[Switch.scala 30:36:@14513.4]
  wire  _T_34994; // @[Switch.scala 30:53:@14515.4]
  wire  valid_45_5; // @[Switch.scala 30:36:@14516.4]
  wire  _T_34997; // @[Switch.scala 30:53:@14518.4]
  wire  valid_45_6; // @[Switch.scala 30:36:@14519.4]
  wire  _T_35000; // @[Switch.scala 30:53:@14521.4]
  wire  valid_45_7; // @[Switch.scala 30:36:@14522.4]
  wire  _T_35003; // @[Switch.scala 30:53:@14524.4]
  wire  valid_45_8; // @[Switch.scala 30:36:@14525.4]
  wire  _T_35006; // @[Switch.scala 30:53:@14527.4]
  wire  valid_45_9; // @[Switch.scala 30:36:@14528.4]
  wire  _T_35009; // @[Switch.scala 30:53:@14530.4]
  wire  valid_45_10; // @[Switch.scala 30:36:@14531.4]
  wire  _T_35012; // @[Switch.scala 30:53:@14533.4]
  wire  valid_45_11; // @[Switch.scala 30:36:@14534.4]
  wire  _T_35015; // @[Switch.scala 30:53:@14536.4]
  wire  valid_45_12; // @[Switch.scala 30:36:@14537.4]
  wire  _T_35018; // @[Switch.scala 30:53:@14539.4]
  wire  valid_45_13; // @[Switch.scala 30:36:@14540.4]
  wire  _T_35021; // @[Switch.scala 30:53:@14542.4]
  wire  valid_45_14; // @[Switch.scala 30:36:@14543.4]
  wire  _T_35024; // @[Switch.scala 30:53:@14545.4]
  wire  valid_45_15; // @[Switch.scala 30:36:@14546.4]
  wire  _T_35027; // @[Switch.scala 30:53:@14548.4]
  wire  valid_45_16; // @[Switch.scala 30:36:@14549.4]
  wire  _T_35030; // @[Switch.scala 30:53:@14551.4]
  wire  valid_45_17; // @[Switch.scala 30:36:@14552.4]
  wire  _T_35033; // @[Switch.scala 30:53:@14554.4]
  wire  valid_45_18; // @[Switch.scala 30:36:@14555.4]
  wire  _T_35036; // @[Switch.scala 30:53:@14557.4]
  wire  valid_45_19; // @[Switch.scala 30:36:@14558.4]
  wire  _T_35039; // @[Switch.scala 30:53:@14560.4]
  wire  valid_45_20; // @[Switch.scala 30:36:@14561.4]
  wire  _T_35042; // @[Switch.scala 30:53:@14563.4]
  wire  valid_45_21; // @[Switch.scala 30:36:@14564.4]
  wire  _T_35045; // @[Switch.scala 30:53:@14566.4]
  wire  valid_45_22; // @[Switch.scala 30:36:@14567.4]
  wire  _T_35048; // @[Switch.scala 30:53:@14569.4]
  wire  valid_45_23; // @[Switch.scala 30:36:@14570.4]
  wire  _T_35051; // @[Switch.scala 30:53:@14572.4]
  wire  valid_45_24; // @[Switch.scala 30:36:@14573.4]
  wire  _T_35054; // @[Switch.scala 30:53:@14575.4]
  wire  valid_45_25; // @[Switch.scala 30:36:@14576.4]
  wire  _T_35057; // @[Switch.scala 30:53:@14578.4]
  wire  valid_45_26; // @[Switch.scala 30:36:@14579.4]
  wire  _T_35060; // @[Switch.scala 30:53:@14581.4]
  wire  valid_45_27; // @[Switch.scala 30:36:@14582.4]
  wire  _T_35063; // @[Switch.scala 30:53:@14584.4]
  wire  valid_45_28; // @[Switch.scala 30:36:@14585.4]
  wire  _T_35066; // @[Switch.scala 30:53:@14587.4]
  wire  valid_45_29; // @[Switch.scala 30:36:@14588.4]
  wire  _T_35069; // @[Switch.scala 30:53:@14590.4]
  wire  valid_45_30; // @[Switch.scala 30:36:@14591.4]
  wire  _T_35072; // @[Switch.scala 30:53:@14593.4]
  wire  valid_45_31; // @[Switch.scala 30:36:@14594.4]
  wire  _T_35075; // @[Switch.scala 30:53:@14596.4]
  wire  valid_45_32; // @[Switch.scala 30:36:@14597.4]
  wire  _T_35078; // @[Switch.scala 30:53:@14599.4]
  wire  valid_45_33; // @[Switch.scala 30:36:@14600.4]
  wire  _T_35081; // @[Switch.scala 30:53:@14602.4]
  wire  valid_45_34; // @[Switch.scala 30:36:@14603.4]
  wire  _T_35084; // @[Switch.scala 30:53:@14605.4]
  wire  valid_45_35; // @[Switch.scala 30:36:@14606.4]
  wire  _T_35087; // @[Switch.scala 30:53:@14608.4]
  wire  valid_45_36; // @[Switch.scala 30:36:@14609.4]
  wire  _T_35090; // @[Switch.scala 30:53:@14611.4]
  wire  valid_45_37; // @[Switch.scala 30:36:@14612.4]
  wire  _T_35093; // @[Switch.scala 30:53:@14614.4]
  wire  valid_45_38; // @[Switch.scala 30:36:@14615.4]
  wire  _T_35096; // @[Switch.scala 30:53:@14617.4]
  wire  valid_45_39; // @[Switch.scala 30:36:@14618.4]
  wire  _T_35099; // @[Switch.scala 30:53:@14620.4]
  wire  valid_45_40; // @[Switch.scala 30:36:@14621.4]
  wire  _T_35102; // @[Switch.scala 30:53:@14623.4]
  wire  valid_45_41; // @[Switch.scala 30:36:@14624.4]
  wire  _T_35105; // @[Switch.scala 30:53:@14626.4]
  wire  valid_45_42; // @[Switch.scala 30:36:@14627.4]
  wire  _T_35108; // @[Switch.scala 30:53:@14629.4]
  wire  valid_45_43; // @[Switch.scala 30:36:@14630.4]
  wire  _T_35111; // @[Switch.scala 30:53:@14632.4]
  wire  valid_45_44; // @[Switch.scala 30:36:@14633.4]
  wire  _T_35114; // @[Switch.scala 30:53:@14635.4]
  wire  valid_45_45; // @[Switch.scala 30:36:@14636.4]
  wire  _T_35117; // @[Switch.scala 30:53:@14638.4]
  wire  valid_45_46; // @[Switch.scala 30:36:@14639.4]
  wire  _T_35120; // @[Switch.scala 30:53:@14641.4]
  wire  valid_45_47; // @[Switch.scala 30:36:@14642.4]
  wire  _T_35123; // @[Switch.scala 30:53:@14644.4]
  wire  valid_45_48; // @[Switch.scala 30:36:@14645.4]
  wire  _T_35126; // @[Switch.scala 30:53:@14647.4]
  wire  valid_45_49; // @[Switch.scala 30:36:@14648.4]
  wire  _T_35129; // @[Switch.scala 30:53:@14650.4]
  wire  valid_45_50; // @[Switch.scala 30:36:@14651.4]
  wire  _T_35132; // @[Switch.scala 30:53:@14653.4]
  wire  valid_45_51; // @[Switch.scala 30:36:@14654.4]
  wire  _T_35135; // @[Switch.scala 30:53:@14656.4]
  wire  valid_45_52; // @[Switch.scala 30:36:@14657.4]
  wire  _T_35138; // @[Switch.scala 30:53:@14659.4]
  wire  valid_45_53; // @[Switch.scala 30:36:@14660.4]
  wire  _T_35141; // @[Switch.scala 30:53:@14662.4]
  wire  valid_45_54; // @[Switch.scala 30:36:@14663.4]
  wire  _T_35144; // @[Switch.scala 30:53:@14665.4]
  wire  valid_45_55; // @[Switch.scala 30:36:@14666.4]
  wire  _T_35147; // @[Switch.scala 30:53:@14668.4]
  wire  valid_45_56; // @[Switch.scala 30:36:@14669.4]
  wire  _T_35150; // @[Switch.scala 30:53:@14671.4]
  wire  valid_45_57; // @[Switch.scala 30:36:@14672.4]
  wire  _T_35153; // @[Switch.scala 30:53:@14674.4]
  wire  valid_45_58; // @[Switch.scala 30:36:@14675.4]
  wire  _T_35156; // @[Switch.scala 30:53:@14677.4]
  wire  valid_45_59; // @[Switch.scala 30:36:@14678.4]
  wire  _T_35159; // @[Switch.scala 30:53:@14680.4]
  wire  valid_45_60; // @[Switch.scala 30:36:@14681.4]
  wire  _T_35162; // @[Switch.scala 30:53:@14683.4]
  wire  valid_45_61; // @[Switch.scala 30:36:@14684.4]
  wire  _T_35165; // @[Switch.scala 30:53:@14686.4]
  wire  valid_45_62; // @[Switch.scala 30:36:@14687.4]
  wire  _T_35168; // @[Switch.scala 30:53:@14689.4]
  wire  valid_45_63; // @[Switch.scala 30:36:@14690.4]
  wire [5:0] _T_35234; // @[Mux.scala 31:69:@14692.4]
  wire [5:0] _T_35235; // @[Mux.scala 31:69:@14693.4]
  wire [5:0] _T_35236; // @[Mux.scala 31:69:@14694.4]
  wire [5:0] _T_35237; // @[Mux.scala 31:69:@14695.4]
  wire [5:0] _T_35238; // @[Mux.scala 31:69:@14696.4]
  wire [5:0] _T_35239; // @[Mux.scala 31:69:@14697.4]
  wire [5:0] _T_35240; // @[Mux.scala 31:69:@14698.4]
  wire [5:0] _T_35241; // @[Mux.scala 31:69:@14699.4]
  wire [5:0] _T_35242; // @[Mux.scala 31:69:@14700.4]
  wire [5:0] _T_35243; // @[Mux.scala 31:69:@14701.4]
  wire [5:0] _T_35244; // @[Mux.scala 31:69:@14702.4]
  wire [5:0] _T_35245; // @[Mux.scala 31:69:@14703.4]
  wire [5:0] _T_35246; // @[Mux.scala 31:69:@14704.4]
  wire [5:0] _T_35247; // @[Mux.scala 31:69:@14705.4]
  wire [5:0] _T_35248; // @[Mux.scala 31:69:@14706.4]
  wire [5:0] _T_35249; // @[Mux.scala 31:69:@14707.4]
  wire [5:0] _T_35250; // @[Mux.scala 31:69:@14708.4]
  wire [5:0] _T_35251; // @[Mux.scala 31:69:@14709.4]
  wire [5:0] _T_35252; // @[Mux.scala 31:69:@14710.4]
  wire [5:0] _T_35253; // @[Mux.scala 31:69:@14711.4]
  wire [5:0] _T_35254; // @[Mux.scala 31:69:@14712.4]
  wire [5:0] _T_35255; // @[Mux.scala 31:69:@14713.4]
  wire [5:0] _T_35256; // @[Mux.scala 31:69:@14714.4]
  wire [5:0] _T_35257; // @[Mux.scala 31:69:@14715.4]
  wire [5:0] _T_35258; // @[Mux.scala 31:69:@14716.4]
  wire [5:0] _T_35259; // @[Mux.scala 31:69:@14717.4]
  wire [5:0] _T_35260; // @[Mux.scala 31:69:@14718.4]
  wire [5:0] _T_35261; // @[Mux.scala 31:69:@14719.4]
  wire [5:0] _T_35262; // @[Mux.scala 31:69:@14720.4]
  wire [5:0] _T_35263; // @[Mux.scala 31:69:@14721.4]
  wire [5:0] _T_35264; // @[Mux.scala 31:69:@14722.4]
  wire [5:0] _T_35265; // @[Mux.scala 31:69:@14723.4]
  wire [5:0] _T_35266; // @[Mux.scala 31:69:@14724.4]
  wire [5:0] _T_35267; // @[Mux.scala 31:69:@14725.4]
  wire [5:0] _T_35268; // @[Mux.scala 31:69:@14726.4]
  wire [5:0] _T_35269; // @[Mux.scala 31:69:@14727.4]
  wire [5:0] _T_35270; // @[Mux.scala 31:69:@14728.4]
  wire [5:0] _T_35271; // @[Mux.scala 31:69:@14729.4]
  wire [5:0] _T_35272; // @[Mux.scala 31:69:@14730.4]
  wire [5:0] _T_35273; // @[Mux.scala 31:69:@14731.4]
  wire [5:0] _T_35274; // @[Mux.scala 31:69:@14732.4]
  wire [5:0] _T_35275; // @[Mux.scala 31:69:@14733.4]
  wire [5:0] _T_35276; // @[Mux.scala 31:69:@14734.4]
  wire [5:0] _T_35277; // @[Mux.scala 31:69:@14735.4]
  wire [5:0] _T_35278; // @[Mux.scala 31:69:@14736.4]
  wire [5:0] _T_35279; // @[Mux.scala 31:69:@14737.4]
  wire [5:0] _T_35280; // @[Mux.scala 31:69:@14738.4]
  wire [5:0] _T_35281; // @[Mux.scala 31:69:@14739.4]
  wire [5:0] _T_35282; // @[Mux.scala 31:69:@14740.4]
  wire [5:0] _T_35283; // @[Mux.scala 31:69:@14741.4]
  wire [5:0] _T_35284; // @[Mux.scala 31:69:@14742.4]
  wire [5:0] _T_35285; // @[Mux.scala 31:69:@14743.4]
  wire [5:0] _T_35286; // @[Mux.scala 31:69:@14744.4]
  wire [5:0] _T_35287; // @[Mux.scala 31:69:@14745.4]
  wire [5:0] _T_35288; // @[Mux.scala 31:69:@14746.4]
  wire [5:0] _T_35289; // @[Mux.scala 31:69:@14747.4]
  wire [5:0] _T_35290; // @[Mux.scala 31:69:@14748.4]
  wire [5:0] _T_35291; // @[Mux.scala 31:69:@14749.4]
  wire [5:0] _T_35292; // @[Mux.scala 31:69:@14750.4]
  wire [5:0] _T_35293; // @[Mux.scala 31:69:@14751.4]
  wire [5:0] _T_35294; // @[Mux.scala 31:69:@14752.4]
  wire [5:0] _T_35295; // @[Mux.scala 31:69:@14753.4]
  wire [5:0] select_45; // @[Mux.scala 31:69:@14754.4]
  wire [47:0] _GEN_2881; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2882; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2883; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2884; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2885; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2886; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2887; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2888; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2889; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2890; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2891; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2892; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2893; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2894; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2895; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2896; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2897; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2898; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2899; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2900; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2901; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2902; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2903; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2904; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2905; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2906; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2907; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2908; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2909; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2910; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2911; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2912; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2913; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2914; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2915; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2916; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2917; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2918; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2919; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2920; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2921; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2922; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2923; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2924; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2925; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2926; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2927; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2928; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2929; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2930; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2931; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2932; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2933; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2934; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2935; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2936; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2937; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2938; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2939; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2940; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2941; // @[Switch.scala 33:19:@14756.4]
  wire [47:0] _GEN_2942; // @[Switch.scala 33:19:@14756.4]
  wire [7:0] _T_35304; // @[Switch.scala 34:32:@14763.4]
  wire [15:0] _T_35312; // @[Switch.scala 34:32:@14771.4]
  wire [7:0] _T_35319; // @[Switch.scala 34:32:@14778.4]
  wire [31:0] _T_35328; // @[Switch.scala 34:32:@14787.4]
  wire [7:0] _T_35335; // @[Switch.scala 34:32:@14794.4]
  wire [15:0] _T_35343; // @[Switch.scala 34:32:@14802.4]
  wire [7:0] _T_35350; // @[Switch.scala 34:32:@14809.4]
  wire [31:0] _T_35359; // @[Switch.scala 34:32:@14818.4]
  wire [63:0] _T_35360; // @[Switch.scala 34:32:@14819.4]
  wire  _T_35364; // @[Switch.scala 30:53:@14822.4]
  wire  valid_46_0; // @[Switch.scala 30:36:@14823.4]
  wire  _T_35367; // @[Switch.scala 30:53:@14825.4]
  wire  valid_46_1; // @[Switch.scala 30:36:@14826.4]
  wire  _T_35370; // @[Switch.scala 30:53:@14828.4]
  wire  valid_46_2; // @[Switch.scala 30:36:@14829.4]
  wire  _T_35373; // @[Switch.scala 30:53:@14831.4]
  wire  valid_46_3; // @[Switch.scala 30:36:@14832.4]
  wire  _T_35376; // @[Switch.scala 30:53:@14834.4]
  wire  valid_46_4; // @[Switch.scala 30:36:@14835.4]
  wire  _T_35379; // @[Switch.scala 30:53:@14837.4]
  wire  valid_46_5; // @[Switch.scala 30:36:@14838.4]
  wire  _T_35382; // @[Switch.scala 30:53:@14840.4]
  wire  valid_46_6; // @[Switch.scala 30:36:@14841.4]
  wire  _T_35385; // @[Switch.scala 30:53:@14843.4]
  wire  valid_46_7; // @[Switch.scala 30:36:@14844.4]
  wire  _T_35388; // @[Switch.scala 30:53:@14846.4]
  wire  valid_46_8; // @[Switch.scala 30:36:@14847.4]
  wire  _T_35391; // @[Switch.scala 30:53:@14849.4]
  wire  valid_46_9; // @[Switch.scala 30:36:@14850.4]
  wire  _T_35394; // @[Switch.scala 30:53:@14852.4]
  wire  valid_46_10; // @[Switch.scala 30:36:@14853.4]
  wire  _T_35397; // @[Switch.scala 30:53:@14855.4]
  wire  valid_46_11; // @[Switch.scala 30:36:@14856.4]
  wire  _T_35400; // @[Switch.scala 30:53:@14858.4]
  wire  valid_46_12; // @[Switch.scala 30:36:@14859.4]
  wire  _T_35403; // @[Switch.scala 30:53:@14861.4]
  wire  valid_46_13; // @[Switch.scala 30:36:@14862.4]
  wire  _T_35406; // @[Switch.scala 30:53:@14864.4]
  wire  valid_46_14; // @[Switch.scala 30:36:@14865.4]
  wire  _T_35409; // @[Switch.scala 30:53:@14867.4]
  wire  valid_46_15; // @[Switch.scala 30:36:@14868.4]
  wire  _T_35412; // @[Switch.scala 30:53:@14870.4]
  wire  valid_46_16; // @[Switch.scala 30:36:@14871.4]
  wire  _T_35415; // @[Switch.scala 30:53:@14873.4]
  wire  valid_46_17; // @[Switch.scala 30:36:@14874.4]
  wire  _T_35418; // @[Switch.scala 30:53:@14876.4]
  wire  valid_46_18; // @[Switch.scala 30:36:@14877.4]
  wire  _T_35421; // @[Switch.scala 30:53:@14879.4]
  wire  valid_46_19; // @[Switch.scala 30:36:@14880.4]
  wire  _T_35424; // @[Switch.scala 30:53:@14882.4]
  wire  valid_46_20; // @[Switch.scala 30:36:@14883.4]
  wire  _T_35427; // @[Switch.scala 30:53:@14885.4]
  wire  valid_46_21; // @[Switch.scala 30:36:@14886.4]
  wire  _T_35430; // @[Switch.scala 30:53:@14888.4]
  wire  valid_46_22; // @[Switch.scala 30:36:@14889.4]
  wire  _T_35433; // @[Switch.scala 30:53:@14891.4]
  wire  valid_46_23; // @[Switch.scala 30:36:@14892.4]
  wire  _T_35436; // @[Switch.scala 30:53:@14894.4]
  wire  valid_46_24; // @[Switch.scala 30:36:@14895.4]
  wire  _T_35439; // @[Switch.scala 30:53:@14897.4]
  wire  valid_46_25; // @[Switch.scala 30:36:@14898.4]
  wire  _T_35442; // @[Switch.scala 30:53:@14900.4]
  wire  valid_46_26; // @[Switch.scala 30:36:@14901.4]
  wire  _T_35445; // @[Switch.scala 30:53:@14903.4]
  wire  valid_46_27; // @[Switch.scala 30:36:@14904.4]
  wire  _T_35448; // @[Switch.scala 30:53:@14906.4]
  wire  valid_46_28; // @[Switch.scala 30:36:@14907.4]
  wire  _T_35451; // @[Switch.scala 30:53:@14909.4]
  wire  valid_46_29; // @[Switch.scala 30:36:@14910.4]
  wire  _T_35454; // @[Switch.scala 30:53:@14912.4]
  wire  valid_46_30; // @[Switch.scala 30:36:@14913.4]
  wire  _T_35457; // @[Switch.scala 30:53:@14915.4]
  wire  valid_46_31; // @[Switch.scala 30:36:@14916.4]
  wire  _T_35460; // @[Switch.scala 30:53:@14918.4]
  wire  valid_46_32; // @[Switch.scala 30:36:@14919.4]
  wire  _T_35463; // @[Switch.scala 30:53:@14921.4]
  wire  valid_46_33; // @[Switch.scala 30:36:@14922.4]
  wire  _T_35466; // @[Switch.scala 30:53:@14924.4]
  wire  valid_46_34; // @[Switch.scala 30:36:@14925.4]
  wire  _T_35469; // @[Switch.scala 30:53:@14927.4]
  wire  valid_46_35; // @[Switch.scala 30:36:@14928.4]
  wire  _T_35472; // @[Switch.scala 30:53:@14930.4]
  wire  valid_46_36; // @[Switch.scala 30:36:@14931.4]
  wire  _T_35475; // @[Switch.scala 30:53:@14933.4]
  wire  valid_46_37; // @[Switch.scala 30:36:@14934.4]
  wire  _T_35478; // @[Switch.scala 30:53:@14936.4]
  wire  valid_46_38; // @[Switch.scala 30:36:@14937.4]
  wire  _T_35481; // @[Switch.scala 30:53:@14939.4]
  wire  valid_46_39; // @[Switch.scala 30:36:@14940.4]
  wire  _T_35484; // @[Switch.scala 30:53:@14942.4]
  wire  valid_46_40; // @[Switch.scala 30:36:@14943.4]
  wire  _T_35487; // @[Switch.scala 30:53:@14945.4]
  wire  valid_46_41; // @[Switch.scala 30:36:@14946.4]
  wire  _T_35490; // @[Switch.scala 30:53:@14948.4]
  wire  valid_46_42; // @[Switch.scala 30:36:@14949.4]
  wire  _T_35493; // @[Switch.scala 30:53:@14951.4]
  wire  valid_46_43; // @[Switch.scala 30:36:@14952.4]
  wire  _T_35496; // @[Switch.scala 30:53:@14954.4]
  wire  valid_46_44; // @[Switch.scala 30:36:@14955.4]
  wire  _T_35499; // @[Switch.scala 30:53:@14957.4]
  wire  valid_46_45; // @[Switch.scala 30:36:@14958.4]
  wire  _T_35502; // @[Switch.scala 30:53:@14960.4]
  wire  valid_46_46; // @[Switch.scala 30:36:@14961.4]
  wire  _T_35505; // @[Switch.scala 30:53:@14963.4]
  wire  valid_46_47; // @[Switch.scala 30:36:@14964.4]
  wire  _T_35508; // @[Switch.scala 30:53:@14966.4]
  wire  valid_46_48; // @[Switch.scala 30:36:@14967.4]
  wire  _T_35511; // @[Switch.scala 30:53:@14969.4]
  wire  valid_46_49; // @[Switch.scala 30:36:@14970.4]
  wire  _T_35514; // @[Switch.scala 30:53:@14972.4]
  wire  valid_46_50; // @[Switch.scala 30:36:@14973.4]
  wire  _T_35517; // @[Switch.scala 30:53:@14975.4]
  wire  valid_46_51; // @[Switch.scala 30:36:@14976.4]
  wire  _T_35520; // @[Switch.scala 30:53:@14978.4]
  wire  valid_46_52; // @[Switch.scala 30:36:@14979.4]
  wire  _T_35523; // @[Switch.scala 30:53:@14981.4]
  wire  valid_46_53; // @[Switch.scala 30:36:@14982.4]
  wire  _T_35526; // @[Switch.scala 30:53:@14984.4]
  wire  valid_46_54; // @[Switch.scala 30:36:@14985.4]
  wire  _T_35529; // @[Switch.scala 30:53:@14987.4]
  wire  valid_46_55; // @[Switch.scala 30:36:@14988.4]
  wire  _T_35532; // @[Switch.scala 30:53:@14990.4]
  wire  valid_46_56; // @[Switch.scala 30:36:@14991.4]
  wire  _T_35535; // @[Switch.scala 30:53:@14993.4]
  wire  valid_46_57; // @[Switch.scala 30:36:@14994.4]
  wire  _T_35538; // @[Switch.scala 30:53:@14996.4]
  wire  valid_46_58; // @[Switch.scala 30:36:@14997.4]
  wire  _T_35541; // @[Switch.scala 30:53:@14999.4]
  wire  valid_46_59; // @[Switch.scala 30:36:@15000.4]
  wire  _T_35544; // @[Switch.scala 30:53:@15002.4]
  wire  valid_46_60; // @[Switch.scala 30:36:@15003.4]
  wire  _T_35547; // @[Switch.scala 30:53:@15005.4]
  wire  valid_46_61; // @[Switch.scala 30:36:@15006.4]
  wire  _T_35550; // @[Switch.scala 30:53:@15008.4]
  wire  valid_46_62; // @[Switch.scala 30:36:@15009.4]
  wire  _T_35553; // @[Switch.scala 30:53:@15011.4]
  wire  valid_46_63; // @[Switch.scala 30:36:@15012.4]
  wire [5:0] _T_35619; // @[Mux.scala 31:69:@15014.4]
  wire [5:0] _T_35620; // @[Mux.scala 31:69:@15015.4]
  wire [5:0] _T_35621; // @[Mux.scala 31:69:@15016.4]
  wire [5:0] _T_35622; // @[Mux.scala 31:69:@15017.4]
  wire [5:0] _T_35623; // @[Mux.scala 31:69:@15018.4]
  wire [5:0] _T_35624; // @[Mux.scala 31:69:@15019.4]
  wire [5:0] _T_35625; // @[Mux.scala 31:69:@15020.4]
  wire [5:0] _T_35626; // @[Mux.scala 31:69:@15021.4]
  wire [5:0] _T_35627; // @[Mux.scala 31:69:@15022.4]
  wire [5:0] _T_35628; // @[Mux.scala 31:69:@15023.4]
  wire [5:0] _T_35629; // @[Mux.scala 31:69:@15024.4]
  wire [5:0] _T_35630; // @[Mux.scala 31:69:@15025.4]
  wire [5:0] _T_35631; // @[Mux.scala 31:69:@15026.4]
  wire [5:0] _T_35632; // @[Mux.scala 31:69:@15027.4]
  wire [5:0] _T_35633; // @[Mux.scala 31:69:@15028.4]
  wire [5:0] _T_35634; // @[Mux.scala 31:69:@15029.4]
  wire [5:0] _T_35635; // @[Mux.scala 31:69:@15030.4]
  wire [5:0] _T_35636; // @[Mux.scala 31:69:@15031.4]
  wire [5:0] _T_35637; // @[Mux.scala 31:69:@15032.4]
  wire [5:0] _T_35638; // @[Mux.scala 31:69:@15033.4]
  wire [5:0] _T_35639; // @[Mux.scala 31:69:@15034.4]
  wire [5:0] _T_35640; // @[Mux.scala 31:69:@15035.4]
  wire [5:0] _T_35641; // @[Mux.scala 31:69:@15036.4]
  wire [5:0] _T_35642; // @[Mux.scala 31:69:@15037.4]
  wire [5:0] _T_35643; // @[Mux.scala 31:69:@15038.4]
  wire [5:0] _T_35644; // @[Mux.scala 31:69:@15039.4]
  wire [5:0] _T_35645; // @[Mux.scala 31:69:@15040.4]
  wire [5:0] _T_35646; // @[Mux.scala 31:69:@15041.4]
  wire [5:0] _T_35647; // @[Mux.scala 31:69:@15042.4]
  wire [5:0] _T_35648; // @[Mux.scala 31:69:@15043.4]
  wire [5:0] _T_35649; // @[Mux.scala 31:69:@15044.4]
  wire [5:0] _T_35650; // @[Mux.scala 31:69:@15045.4]
  wire [5:0] _T_35651; // @[Mux.scala 31:69:@15046.4]
  wire [5:0] _T_35652; // @[Mux.scala 31:69:@15047.4]
  wire [5:0] _T_35653; // @[Mux.scala 31:69:@15048.4]
  wire [5:0] _T_35654; // @[Mux.scala 31:69:@15049.4]
  wire [5:0] _T_35655; // @[Mux.scala 31:69:@15050.4]
  wire [5:0] _T_35656; // @[Mux.scala 31:69:@15051.4]
  wire [5:0] _T_35657; // @[Mux.scala 31:69:@15052.4]
  wire [5:0] _T_35658; // @[Mux.scala 31:69:@15053.4]
  wire [5:0] _T_35659; // @[Mux.scala 31:69:@15054.4]
  wire [5:0] _T_35660; // @[Mux.scala 31:69:@15055.4]
  wire [5:0] _T_35661; // @[Mux.scala 31:69:@15056.4]
  wire [5:0] _T_35662; // @[Mux.scala 31:69:@15057.4]
  wire [5:0] _T_35663; // @[Mux.scala 31:69:@15058.4]
  wire [5:0] _T_35664; // @[Mux.scala 31:69:@15059.4]
  wire [5:0] _T_35665; // @[Mux.scala 31:69:@15060.4]
  wire [5:0] _T_35666; // @[Mux.scala 31:69:@15061.4]
  wire [5:0] _T_35667; // @[Mux.scala 31:69:@15062.4]
  wire [5:0] _T_35668; // @[Mux.scala 31:69:@15063.4]
  wire [5:0] _T_35669; // @[Mux.scala 31:69:@15064.4]
  wire [5:0] _T_35670; // @[Mux.scala 31:69:@15065.4]
  wire [5:0] _T_35671; // @[Mux.scala 31:69:@15066.4]
  wire [5:0] _T_35672; // @[Mux.scala 31:69:@15067.4]
  wire [5:0] _T_35673; // @[Mux.scala 31:69:@15068.4]
  wire [5:0] _T_35674; // @[Mux.scala 31:69:@15069.4]
  wire [5:0] _T_35675; // @[Mux.scala 31:69:@15070.4]
  wire [5:0] _T_35676; // @[Mux.scala 31:69:@15071.4]
  wire [5:0] _T_35677; // @[Mux.scala 31:69:@15072.4]
  wire [5:0] _T_35678; // @[Mux.scala 31:69:@15073.4]
  wire [5:0] _T_35679; // @[Mux.scala 31:69:@15074.4]
  wire [5:0] _T_35680; // @[Mux.scala 31:69:@15075.4]
  wire [5:0] select_46; // @[Mux.scala 31:69:@15076.4]
  wire [47:0] _GEN_2945; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2946; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2947; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2948; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2949; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2950; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2951; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2952; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2953; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2954; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2955; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2956; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2957; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2958; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2959; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2960; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2961; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2962; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2963; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2964; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2965; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2966; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2967; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2968; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2969; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2970; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2971; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2972; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2973; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2974; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2975; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2976; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2977; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2978; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2979; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2980; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2981; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2982; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2983; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2984; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2985; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2986; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2987; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2988; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2989; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2990; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2991; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2992; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2993; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2994; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2995; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2996; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2997; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2998; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_2999; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_3000; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_3001; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_3002; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_3003; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_3004; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_3005; // @[Switch.scala 33:19:@15078.4]
  wire [47:0] _GEN_3006; // @[Switch.scala 33:19:@15078.4]
  wire [7:0] _T_35689; // @[Switch.scala 34:32:@15085.4]
  wire [15:0] _T_35697; // @[Switch.scala 34:32:@15093.4]
  wire [7:0] _T_35704; // @[Switch.scala 34:32:@15100.4]
  wire [31:0] _T_35713; // @[Switch.scala 34:32:@15109.4]
  wire [7:0] _T_35720; // @[Switch.scala 34:32:@15116.4]
  wire [15:0] _T_35728; // @[Switch.scala 34:32:@15124.4]
  wire [7:0] _T_35735; // @[Switch.scala 34:32:@15131.4]
  wire [31:0] _T_35744; // @[Switch.scala 34:32:@15140.4]
  wire [63:0] _T_35745; // @[Switch.scala 34:32:@15141.4]
  wire  _T_35749; // @[Switch.scala 30:53:@15144.4]
  wire  valid_47_0; // @[Switch.scala 30:36:@15145.4]
  wire  _T_35752; // @[Switch.scala 30:53:@15147.4]
  wire  valid_47_1; // @[Switch.scala 30:36:@15148.4]
  wire  _T_35755; // @[Switch.scala 30:53:@15150.4]
  wire  valid_47_2; // @[Switch.scala 30:36:@15151.4]
  wire  _T_35758; // @[Switch.scala 30:53:@15153.4]
  wire  valid_47_3; // @[Switch.scala 30:36:@15154.4]
  wire  _T_35761; // @[Switch.scala 30:53:@15156.4]
  wire  valid_47_4; // @[Switch.scala 30:36:@15157.4]
  wire  _T_35764; // @[Switch.scala 30:53:@15159.4]
  wire  valid_47_5; // @[Switch.scala 30:36:@15160.4]
  wire  _T_35767; // @[Switch.scala 30:53:@15162.4]
  wire  valid_47_6; // @[Switch.scala 30:36:@15163.4]
  wire  _T_35770; // @[Switch.scala 30:53:@15165.4]
  wire  valid_47_7; // @[Switch.scala 30:36:@15166.4]
  wire  _T_35773; // @[Switch.scala 30:53:@15168.4]
  wire  valid_47_8; // @[Switch.scala 30:36:@15169.4]
  wire  _T_35776; // @[Switch.scala 30:53:@15171.4]
  wire  valid_47_9; // @[Switch.scala 30:36:@15172.4]
  wire  _T_35779; // @[Switch.scala 30:53:@15174.4]
  wire  valid_47_10; // @[Switch.scala 30:36:@15175.4]
  wire  _T_35782; // @[Switch.scala 30:53:@15177.4]
  wire  valid_47_11; // @[Switch.scala 30:36:@15178.4]
  wire  _T_35785; // @[Switch.scala 30:53:@15180.4]
  wire  valid_47_12; // @[Switch.scala 30:36:@15181.4]
  wire  _T_35788; // @[Switch.scala 30:53:@15183.4]
  wire  valid_47_13; // @[Switch.scala 30:36:@15184.4]
  wire  _T_35791; // @[Switch.scala 30:53:@15186.4]
  wire  valid_47_14; // @[Switch.scala 30:36:@15187.4]
  wire  _T_35794; // @[Switch.scala 30:53:@15189.4]
  wire  valid_47_15; // @[Switch.scala 30:36:@15190.4]
  wire  _T_35797; // @[Switch.scala 30:53:@15192.4]
  wire  valid_47_16; // @[Switch.scala 30:36:@15193.4]
  wire  _T_35800; // @[Switch.scala 30:53:@15195.4]
  wire  valid_47_17; // @[Switch.scala 30:36:@15196.4]
  wire  _T_35803; // @[Switch.scala 30:53:@15198.4]
  wire  valid_47_18; // @[Switch.scala 30:36:@15199.4]
  wire  _T_35806; // @[Switch.scala 30:53:@15201.4]
  wire  valid_47_19; // @[Switch.scala 30:36:@15202.4]
  wire  _T_35809; // @[Switch.scala 30:53:@15204.4]
  wire  valid_47_20; // @[Switch.scala 30:36:@15205.4]
  wire  _T_35812; // @[Switch.scala 30:53:@15207.4]
  wire  valid_47_21; // @[Switch.scala 30:36:@15208.4]
  wire  _T_35815; // @[Switch.scala 30:53:@15210.4]
  wire  valid_47_22; // @[Switch.scala 30:36:@15211.4]
  wire  _T_35818; // @[Switch.scala 30:53:@15213.4]
  wire  valid_47_23; // @[Switch.scala 30:36:@15214.4]
  wire  _T_35821; // @[Switch.scala 30:53:@15216.4]
  wire  valid_47_24; // @[Switch.scala 30:36:@15217.4]
  wire  _T_35824; // @[Switch.scala 30:53:@15219.4]
  wire  valid_47_25; // @[Switch.scala 30:36:@15220.4]
  wire  _T_35827; // @[Switch.scala 30:53:@15222.4]
  wire  valid_47_26; // @[Switch.scala 30:36:@15223.4]
  wire  _T_35830; // @[Switch.scala 30:53:@15225.4]
  wire  valid_47_27; // @[Switch.scala 30:36:@15226.4]
  wire  _T_35833; // @[Switch.scala 30:53:@15228.4]
  wire  valid_47_28; // @[Switch.scala 30:36:@15229.4]
  wire  _T_35836; // @[Switch.scala 30:53:@15231.4]
  wire  valid_47_29; // @[Switch.scala 30:36:@15232.4]
  wire  _T_35839; // @[Switch.scala 30:53:@15234.4]
  wire  valid_47_30; // @[Switch.scala 30:36:@15235.4]
  wire  _T_35842; // @[Switch.scala 30:53:@15237.4]
  wire  valid_47_31; // @[Switch.scala 30:36:@15238.4]
  wire  _T_35845; // @[Switch.scala 30:53:@15240.4]
  wire  valid_47_32; // @[Switch.scala 30:36:@15241.4]
  wire  _T_35848; // @[Switch.scala 30:53:@15243.4]
  wire  valid_47_33; // @[Switch.scala 30:36:@15244.4]
  wire  _T_35851; // @[Switch.scala 30:53:@15246.4]
  wire  valid_47_34; // @[Switch.scala 30:36:@15247.4]
  wire  _T_35854; // @[Switch.scala 30:53:@15249.4]
  wire  valid_47_35; // @[Switch.scala 30:36:@15250.4]
  wire  _T_35857; // @[Switch.scala 30:53:@15252.4]
  wire  valid_47_36; // @[Switch.scala 30:36:@15253.4]
  wire  _T_35860; // @[Switch.scala 30:53:@15255.4]
  wire  valid_47_37; // @[Switch.scala 30:36:@15256.4]
  wire  _T_35863; // @[Switch.scala 30:53:@15258.4]
  wire  valid_47_38; // @[Switch.scala 30:36:@15259.4]
  wire  _T_35866; // @[Switch.scala 30:53:@15261.4]
  wire  valid_47_39; // @[Switch.scala 30:36:@15262.4]
  wire  _T_35869; // @[Switch.scala 30:53:@15264.4]
  wire  valid_47_40; // @[Switch.scala 30:36:@15265.4]
  wire  _T_35872; // @[Switch.scala 30:53:@15267.4]
  wire  valid_47_41; // @[Switch.scala 30:36:@15268.4]
  wire  _T_35875; // @[Switch.scala 30:53:@15270.4]
  wire  valid_47_42; // @[Switch.scala 30:36:@15271.4]
  wire  _T_35878; // @[Switch.scala 30:53:@15273.4]
  wire  valid_47_43; // @[Switch.scala 30:36:@15274.4]
  wire  _T_35881; // @[Switch.scala 30:53:@15276.4]
  wire  valid_47_44; // @[Switch.scala 30:36:@15277.4]
  wire  _T_35884; // @[Switch.scala 30:53:@15279.4]
  wire  valid_47_45; // @[Switch.scala 30:36:@15280.4]
  wire  _T_35887; // @[Switch.scala 30:53:@15282.4]
  wire  valid_47_46; // @[Switch.scala 30:36:@15283.4]
  wire  _T_35890; // @[Switch.scala 30:53:@15285.4]
  wire  valid_47_47; // @[Switch.scala 30:36:@15286.4]
  wire  _T_35893; // @[Switch.scala 30:53:@15288.4]
  wire  valid_47_48; // @[Switch.scala 30:36:@15289.4]
  wire  _T_35896; // @[Switch.scala 30:53:@15291.4]
  wire  valid_47_49; // @[Switch.scala 30:36:@15292.4]
  wire  _T_35899; // @[Switch.scala 30:53:@15294.4]
  wire  valid_47_50; // @[Switch.scala 30:36:@15295.4]
  wire  _T_35902; // @[Switch.scala 30:53:@15297.4]
  wire  valid_47_51; // @[Switch.scala 30:36:@15298.4]
  wire  _T_35905; // @[Switch.scala 30:53:@15300.4]
  wire  valid_47_52; // @[Switch.scala 30:36:@15301.4]
  wire  _T_35908; // @[Switch.scala 30:53:@15303.4]
  wire  valid_47_53; // @[Switch.scala 30:36:@15304.4]
  wire  _T_35911; // @[Switch.scala 30:53:@15306.4]
  wire  valid_47_54; // @[Switch.scala 30:36:@15307.4]
  wire  _T_35914; // @[Switch.scala 30:53:@15309.4]
  wire  valid_47_55; // @[Switch.scala 30:36:@15310.4]
  wire  _T_35917; // @[Switch.scala 30:53:@15312.4]
  wire  valid_47_56; // @[Switch.scala 30:36:@15313.4]
  wire  _T_35920; // @[Switch.scala 30:53:@15315.4]
  wire  valid_47_57; // @[Switch.scala 30:36:@15316.4]
  wire  _T_35923; // @[Switch.scala 30:53:@15318.4]
  wire  valid_47_58; // @[Switch.scala 30:36:@15319.4]
  wire  _T_35926; // @[Switch.scala 30:53:@15321.4]
  wire  valid_47_59; // @[Switch.scala 30:36:@15322.4]
  wire  _T_35929; // @[Switch.scala 30:53:@15324.4]
  wire  valid_47_60; // @[Switch.scala 30:36:@15325.4]
  wire  _T_35932; // @[Switch.scala 30:53:@15327.4]
  wire  valid_47_61; // @[Switch.scala 30:36:@15328.4]
  wire  _T_35935; // @[Switch.scala 30:53:@15330.4]
  wire  valid_47_62; // @[Switch.scala 30:36:@15331.4]
  wire  _T_35938; // @[Switch.scala 30:53:@15333.4]
  wire  valid_47_63; // @[Switch.scala 30:36:@15334.4]
  wire [5:0] _T_36004; // @[Mux.scala 31:69:@15336.4]
  wire [5:0] _T_36005; // @[Mux.scala 31:69:@15337.4]
  wire [5:0] _T_36006; // @[Mux.scala 31:69:@15338.4]
  wire [5:0] _T_36007; // @[Mux.scala 31:69:@15339.4]
  wire [5:0] _T_36008; // @[Mux.scala 31:69:@15340.4]
  wire [5:0] _T_36009; // @[Mux.scala 31:69:@15341.4]
  wire [5:0] _T_36010; // @[Mux.scala 31:69:@15342.4]
  wire [5:0] _T_36011; // @[Mux.scala 31:69:@15343.4]
  wire [5:0] _T_36012; // @[Mux.scala 31:69:@15344.4]
  wire [5:0] _T_36013; // @[Mux.scala 31:69:@15345.4]
  wire [5:0] _T_36014; // @[Mux.scala 31:69:@15346.4]
  wire [5:0] _T_36015; // @[Mux.scala 31:69:@15347.4]
  wire [5:0] _T_36016; // @[Mux.scala 31:69:@15348.4]
  wire [5:0] _T_36017; // @[Mux.scala 31:69:@15349.4]
  wire [5:0] _T_36018; // @[Mux.scala 31:69:@15350.4]
  wire [5:0] _T_36019; // @[Mux.scala 31:69:@15351.4]
  wire [5:0] _T_36020; // @[Mux.scala 31:69:@15352.4]
  wire [5:0] _T_36021; // @[Mux.scala 31:69:@15353.4]
  wire [5:0] _T_36022; // @[Mux.scala 31:69:@15354.4]
  wire [5:0] _T_36023; // @[Mux.scala 31:69:@15355.4]
  wire [5:0] _T_36024; // @[Mux.scala 31:69:@15356.4]
  wire [5:0] _T_36025; // @[Mux.scala 31:69:@15357.4]
  wire [5:0] _T_36026; // @[Mux.scala 31:69:@15358.4]
  wire [5:0] _T_36027; // @[Mux.scala 31:69:@15359.4]
  wire [5:0] _T_36028; // @[Mux.scala 31:69:@15360.4]
  wire [5:0] _T_36029; // @[Mux.scala 31:69:@15361.4]
  wire [5:0] _T_36030; // @[Mux.scala 31:69:@15362.4]
  wire [5:0] _T_36031; // @[Mux.scala 31:69:@15363.4]
  wire [5:0] _T_36032; // @[Mux.scala 31:69:@15364.4]
  wire [5:0] _T_36033; // @[Mux.scala 31:69:@15365.4]
  wire [5:0] _T_36034; // @[Mux.scala 31:69:@15366.4]
  wire [5:0] _T_36035; // @[Mux.scala 31:69:@15367.4]
  wire [5:0] _T_36036; // @[Mux.scala 31:69:@15368.4]
  wire [5:0] _T_36037; // @[Mux.scala 31:69:@15369.4]
  wire [5:0] _T_36038; // @[Mux.scala 31:69:@15370.4]
  wire [5:0] _T_36039; // @[Mux.scala 31:69:@15371.4]
  wire [5:0] _T_36040; // @[Mux.scala 31:69:@15372.4]
  wire [5:0] _T_36041; // @[Mux.scala 31:69:@15373.4]
  wire [5:0] _T_36042; // @[Mux.scala 31:69:@15374.4]
  wire [5:0] _T_36043; // @[Mux.scala 31:69:@15375.4]
  wire [5:0] _T_36044; // @[Mux.scala 31:69:@15376.4]
  wire [5:0] _T_36045; // @[Mux.scala 31:69:@15377.4]
  wire [5:0] _T_36046; // @[Mux.scala 31:69:@15378.4]
  wire [5:0] _T_36047; // @[Mux.scala 31:69:@15379.4]
  wire [5:0] _T_36048; // @[Mux.scala 31:69:@15380.4]
  wire [5:0] _T_36049; // @[Mux.scala 31:69:@15381.4]
  wire [5:0] _T_36050; // @[Mux.scala 31:69:@15382.4]
  wire [5:0] _T_36051; // @[Mux.scala 31:69:@15383.4]
  wire [5:0] _T_36052; // @[Mux.scala 31:69:@15384.4]
  wire [5:0] _T_36053; // @[Mux.scala 31:69:@15385.4]
  wire [5:0] _T_36054; // @[Mux.scala 31:69:@15386.4]
  wire [5:0] _T_36055; // @[Mux.scala 31:69:@15387.4]
  wire [5:0] _T_36056; // @[Mux.scala 31:69:@15388.4]
  wire [5:0] _T_36057; // @[Mux.scala 31:69:@15389.4]
  wire [5:0] _T_36058; // @[Mux.scala 31:69:@15390.4]
  wire [5:0] _T_36059; // @[Mux.scala 31:69:@15391.4]
  wire [5:0] _T_36060; // @[Mux.scala 31:69:@15392.4]
  wire [5:0] _T_36061; // @[Mux.scala 31:69:@15393.4]
  wire [5:0] _T_36062; // @[Mux.scala 31:69:@15394.4]
  wire [5:0] _T_36063; // @[Mux.scala 31:69:@15395.4]
  wire [5:0] _T_36064; // @[Mux.scala 31:69:@15396.4]
  wire [5:0] _T_36065; // @[Mux.scala 31:69:@15397.4]
  wire [5:0] select_47; // @[Mux.scala 31:69:@15398.4]
  wire [47:0] _GEN_3009; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3010; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3011; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3012; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3013; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3014; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3015; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3016; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3017; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3018; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3019; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3020; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3021; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3022; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3023; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3024; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3025; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3026; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3027; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3028; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3029; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3030; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3031; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3032; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3033; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3034; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3035; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3036; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3037; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3038; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3039; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3040; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3041; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3042; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3043; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3044; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3045; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3046; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3047; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3048; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3049; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3050; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3051; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3052; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3053; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3054; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3055; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3056; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3057; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3058; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3059; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3060; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3061; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3062; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3063; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3064; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3065; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3066; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3067; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3068; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3069; // @[Switch.scala 33:19:@15400.4]
  wire [47:0] _GEN_3070; // @[Switch.scala 33:19:@15400.4]
  wire [7:0] _T_36074; // @[Switch.scala 34:32:@15407.4]
  wire [15:0] _T_36082; // @[Switch.scala 34:32:@15415.4]
  wire [7:0] _T_36089; // @[Switch.scala 34:32:@15422.4]
  wire [31:0] _T_36098; // @[Switch.scala 34:32:@15431.4]
  wire [7:0] _T_36105; // @[Switch.scala 34:32:@15438.4]
  wire [15:0] _T_36113; // @[Switch.scala 34:32:@15446.4]
  wire [7:0] _T_36120; // @[Switch.scala 34:32:@15453.4]
  wire [31:0] _T_36129; // @[Switch.scala 34:32:@15462.4]
  wire [63:0] _T_36130; // @[Switch.scala 34:32:@15463.4]
  wire  _T_36134; // @[Switch.scala 30:53:@15466.4]
  wire  valid_48_0; // @[Switch.scala 30:36:@15467.4]
  wire  _T_36137; // @[Switch.scala 30:53:@15469.4]
  wire  valid_48_1; // @[Switch.scala 30:36:@15470.4]
  wire  _T_36140; // @[Switch.scala 30:53:@15472.4]
  wire  valid_48_2; // @[Switch.scala 30:36:@15473.4]
  wire  _T_36143; // @[Switch.scala 30:53:@15475.4]
  wire  valid_48_3; // @[Switch.scala 30:36:@15476.4]
  wire  _T_36146; // @[Switch.scala 30:53:@15478.4]
  wire  valid_48_4; // @[Switch.scala 30:36:@15479.4]
  wire  _T_36149; // @[Switch.scala 30:53:@15481.4]
  wire  valid_48_5; // @[Switch.scala 30:36:@15482.4]
  wire  _T_36152; // @[Switch.scala 30:53:@15484.4]
  wire  valid_48_6; // @[Switch.scala 30:36:@15485.4]
  wire  _T_36155; // @[Switch.scala 30:53:@15487.4]
  wire  valid_48_7; // @[Switch.scala 30:36:@15488.4]
  wire  _T_36158; // @[Switch.scala 30:53:@15490.4]
  wire  valid_48_8; // @[Switch.scala 30:36:@15491.4]
  wire  _T_36161; // @[Switch.scala 30:53:@15493.4]
  wire  valid_48_9; // @[Switch.scala 30:36:@15494.4]
  wire  _T_36164; // @[Switch.scala 30:53:@15496.4]
  wire  valid_48_10; // @[Switch.scala 30:36:@15497.4]
  wire  _T_36167; // @[Switch.scala 30:53:@15499.4]
  wire  valid_48_11; // @[Switch.scala 30:36:@15500.4]
  wire  _T_36170; // @[Switch.scala 30:53:@15502.4]
  wire  valid_48_12; // @[Switch.scala 30:36:@15503.4]
  wire  _T_36173; // @[Switch.scala 30:53:@15505.4]
  wire  valid_48_13; // @[Switch.scala 30:36:@15506.4]
  wire  _T_36176; // @[Switch.scala 30:53:@15508.4]
  wire  valid_48_14; // @[Switch.scala 30:36:@15509.4]
  wire  _T_36179; // @[Switch.scala 30:53:@15511.4]
  wire  valid_48_15; // @[Switch.scala 30:36:@15512.4]
  wire  _T_36182; // @[Switch.scala 30:53:@15514.4]
  wire  valid_48_16; // @[Switch.scala 30:36:@15515.4]
  wire  _T_36185; // @[Switch.scala 30:53:@15517.4]
  wire  valid_48_17; // @[Switch.scala 30:36:@15518.4]
  wire  _T_36188; // @[Switch.scala 30:53:@15520.4]
  wire  valid_48_18; // @[Switch.scala 30:36:@15521.4]
  wire  _T_36191; // @[Switch.scala 30:53:@15523.4]
  wire  valid_48_19; // @[Switch.scala 30:36:@15524.4]
  wire  _T_36194; // @[Switch.scala 30:53:@15526.4]
  wire  valid_48_20; // @[Switch.scala 30:36:@15527.4]
  wire  _T_36197; // @[Switch.scala 30:53:@15529.4]
  wire  valid_48_21; // @[Switch.scala 30:36:@15530.4]
  wire  _T_36200; // @[Switch.scala 30:53:@15532.4]
  wire  valid_48_22; // @[Switch.scala 30:36:@15533.4]
  wire  _T_36203; // @[Switch.scala 30:53:@15535.4]
  wire  valid_48_23; // @[Switch.scala 30:36:@15536.4]
  wire  _T_36206; // @[Switch.scala 30:53:@15538.4]
  wire  valid_48_24; // @[Switch.scala 30:36:@15539.4]
  wire  _T_36209; // @[Switch.scala 30:53:@15541.4]
  wire  valid_48_25; // @[Switch.scala 30:36:@15542.4]
  wire  _T_36212; // @[Switch.scala 30:53:@15544.4]
  wire  valid_48_26; // @[Switch.scala 30:36:@15545.4]
  wire  _T_36215; // @[Switch.scala 30:53:@15547.4]
  wire  valid_48_27; // @[Switch.scala 30:36:@15548.4]
  wire  _T_36218; // @[Switch.scala 30:53:@15550.4]
  wire  valid_48_28; // @[Switch.scala 30:36:@15551.4]
  wire  _T_36221; // @[Switch.scala 30:53:@15553.4]
  wire  valid_48_29; // @[Switch.scala 30:36:@15554.4]
  wire  _T_36224; // @[Switch.scala 30:53:@15556.4]
  wire  valid_48_30; // @[Switch.scala 30:36:@15557.4]
  wire  _T_36227; // @[Switch.scala 30:53:@15559.4]
  wire  valid_48_31; // @[Switch.scala 30:36:@15560.4]
  wire  _T_36230; // @[Switch.scala 30:53:@15562.4]
  wire  valid_48_32; // @[Switch.scala 30:36:@15563.4]
  wire  _T_36233; // @[Switch.scala 30:53:@15565.4]
  wire  valid_48_33; // @[Switch.scala 30:36:@15566.4]
  wire  _T_36236; // @[Switch.scala 30:53:@15568.4]
  wire  valid_48_34; // @[Switch.scala 30:36:@15569.4]
  wire  _T_36239; // @[Switch.scala 30:53:@15571.4]
  wire  valid_48_35; // @[Switch.scala 30:36:@15572.4]
  wire  _T_36242; // @[Switch.scala 30:53:@15574.4]
  wire  valid_48_36; // @[Switch.scala 30:36:@15575.4]
  wire  _T_36245; // @[Switch.scala 30:53:@15577.4]
  wire  valid_48_37; // @[Switch.scala 30:36:@15578.4]
  wire  _T_36248; // @[Switch.scala 30:53:@15580.4]
  wire  valid_48_38; // @[Switch.scala 30:36:@15581.4]
  wire  _T_36251; // @[Switch.scala 30:53:@15583.4]
  wire  valid_48_39; // @[Switch.scala 30:36:@15584.4]
  wire  _T_36254; // @[Switch.scala 30:53:@15586.4]
  wire  valid_48_40; // @[Switch.scala 30:36:@15587.4]
  wire  _T_36257; // @[Switch.scala 30:53:@15589.4]
  wire  valid_48_41; // @[Switch.scala 30:36:@15590.4]
  wire  _T_36260; // @[Switch.scala 30:53:@15592.4]
  wire  valid_48_42; // @[Switch.scala 30:36:@15593.4]
  wire  _T_36263; // @[Switch.scala 30:53:@15595.4]
  wire  valid_48_43; // @[Switch.scala 30:36:@15596.4]
  wire  _T_36266; // @[Switch.scala 30:53:@15598.4]
  wire  valid_48_44; // @[Switch.scala 30:36:@15599.4]
  wire  _T_36269; // @[Switch.scala 30:53:@15601.4]
  wire  valid_48_45; // @[Switch.scala 30:36:@15602.4]
  wire  _T_36272; // @[Switch.scala 30:53:@15604.4]
  wire  valid_48_46; // @[Switch.scala 30:36:@15605.4]
  wire  _T_36275; // @[Switch.scala 30:53:@15607.4]
  wire  valid_48_47; // @[Switch.scala 30:36:@15608.4]
  wire  _T_36278; // @[Switch.scala 30:53:@15610.4]
  wire  valid_48_48; // @[Switch.scala 30:36:@15611.4]
  wire  _T_36281; // @[Switch.scala 30:53:@15613.4]
  wire  valid_48_49; // @[Switch.scala 30:36:@15614.4]
  wire  _T_36284; // @[Switch.scala 30:53:@15616.4]
  wire  valid_48_50; // @[Switch.scala 30:36:@15617.4]
  wire  _T_36287; // @[Switch.scala 30:53:@15619.4]
  wire  valid_48_51; // @[Switch.scala 30:36:@15620.4]
  wire  _T_36290; // @[Switch.scala 30:53:@15622.4]
  wire  valid_48_52; // @[Switch.scala 30:36:@15623.4]
  wire  _T_36293; // @[Switch.scala 30:53:@15625.4]
  wire  valid_48_53; // @[Switch.scala 30:36:@15626.4]
  wire  _T_36296; // @[Switch.scala 30:53:@15628.4]
  wire  valid_48_54; // @[Switch.scala 30:36:@15629.4]
  wire  _T_36299; // @[Switch.scala 30:53:@15631.4]
  wire  valid_48_55; // @[Switch.scala 30:36:@15632.4]
  wire  _T_36302; // @[Switch.scala 30:53:@15634.4]
  wire  valid_48_56; // @[Switch.scala 30:36:@15635.4]
  wire  _T_36305; // @[Switch.scala 30:53:@15637.4]
  wire  valid_48_57; // @[Switch.scala 30:36:@15638.4]
  wire  _T_36308; // @[Switch.scala 30:53:@15640.4]
  wire  valid_48_58; // @[Switch.scala 30:36:@15641.4]
  wire  _T_36311; // @[Switch.scala 30:53:@15643.4]
  wire  valid_48_59; // @[Switch.scala 30:36:@15644.4]
  wire  _T_36314; // @[Switch.scala 30:53:@15646.4]
  wire  valid_48_60; // @[Switch.scala 30:36:@15647.4]
  wire  _T_36317; // @[Switch.scala 30:53:@15649.4]
  wire  valid_48_61; // @[Switch.scala 30:36:@15650.4]
  wire  _T_36320; // @[Switch.scala 30:53:@15652.4]
  wire  valid_48_62; // @[Switch.scala 30:36:@15653.4]
  wire  _T_36323; // @[Switch.scala 30:53:@15655.4]
  wire  valid_48_63; // @[Switch.scala 30:36:@15656.4]
  wire [5:0] _T_36389; // @[Mux.scala 31:69:@15658.4]
  wire [5:0] _T_36390; // @[Mux.scala 31:69:@15659.4]
  wire [5:0] _T_36391; // @[Mux.scala 31:69:@15660.4]
  wire [5:0] _T_36392; // @[Mux.scala 31:69:@15661.4]
  wire [5:0] _T_36393; // @[Mux.scala 31:69:@15662.4]
  wire [5:0] _T_36394; // @[Mux.scala 31:69:@15663.4]
  wire [5:0] _T_36395; // @[Mux.scala 31:69:@15664.4]
  wire [5:0] _T_36396; // @[Mux.scala 31:69:@15665.4]
  wire [5:0] _T_36397; // @[Mux.scala 31:69:@15666.4]
  wire [5:0] _T_36398; // @[Mux.scala 31:69:@15667.4]
  wire [5:0] _T_36399; // @[Mux.scala 31:69:@15668.4]
  wire [5:0] _T_36400; // @[Mux.scala 31:69:@15669.4]
  wire [5:0] _T_36401; // @[Mux.scala 31:69:@15670.4]
  wire [5:0] _T_36402; // @[Mux.scala 31:69:@15671.4]
  wire [5:0] _T_36403; // @[Mux.scala 31:69:@15672.4]
  wire [5:0] _T_36404; // @[Mux.scala 31:69:@15673.4]
  wire [5:0] _T_36405; // @[Mux.scala 31:69:@15674.4]
  wire [5:0] _T_36406; // @[Mux.scala 31:69:@15675.4]
  wire [5:0] _T_36407; // @[Mux.scala 31:69:@15676.4]
  wire [5:0] _T_36408; // @[Mux.scala 31:69:@15677.4]
  wire [5:0] _T_36409; // @[Mux.scala 31:69:@15678.4]
  wire [5:0] _T_36410; // @[Mux.scala 31:69:@15679.4]
  wire [5:0] _T_36411; // @[Mux.scala 31:69:@15680.4]
  wire [5:0] _T_36412; // @[Mux.scala 31:69:@15681.4]
  wire [5:0] _T_36413; // @[Mux.scala 31:69:@15682.4]
  wire [5:0] _T_36414; // @[Mux.scala 31:69:@15683.4]
  wire [5:0] _T_36415; // @[Mux.scala 31:69:@15684.4]
  wire [5:0] _T_36416; // @[Mux.scala 31:69:@15685.4]
  wire [5:0] _T_36417; // @[Mux.scala 31:69:@15686.4]
  wire [5:0] _T_36418; // @[Mux.scala 31:69:@15687.4]
  wire [5:0] _T_36419; // @[Mux.scala 31:69:@15688.4]
  wire [5:0] _T_36420; // @[Mux.scala 31:69:@15689.4]
  wire [5:0] _T_36421; // @[Mux.scala 31:69:@15690.4]
  wire [5:0] _T_36422; // @[Mux.scala 31:69:@15691.4]
  wire [5:0] _T_36423; // @[Mux.scala 31:69:@15692.4]
  wire [5:0] _T_36424; // @[Mux.scala 31:69:@15693.4]
  wire [5:0] _T_36425; // @[Mux.scala 31:69:@15694.4]
  wire [5:0] _T_36426; // @[Mux.scala 31:69:@15695.4]
  wire [5:0] _T_36427; // @[Mux.scala 31:69:@15696.4]
  wire [5:0] _T_36428; // @[Mux.scala 31:69:@15697.4]
  wire [5:0] _T_36429; // @[Mux.scala 31:69:@15698.4]
  wire [5:0] _T_36430; // @[Mux.scala 31:69:@15699.4]
  wire [5:0] _T_36431; // @[Mux.scala 31:69:@15700.4]
  wire [5:0] _T_36432; // @[Mux.scala 31:69:@15701.4]
  wire [5:0] _T_36433; // @[Mux.scala 31:69:@15702.4]
  wire [5:0] _T_36434; // @[Mux.scala 31:69:@15703.4]
  wire [5:0] _T_36435; // @[Mux.scala 31:69:@15704.4]
  wire [5:0] _T_36436; // @[Mux.scala 31:69:@15705.4]
  wire [5:0] _T_36437; // @[Mux.scala 31:69:@15706.4]
  wire [5:0] _T_36438; // @[Mux.scala 31:69:@15707.4]
  wire [5:0] _T_36439; // @[Mux.scala 31:69:@15708.4]
  wire [5:0] _T_36440; // @[Mux.scala 31:69:@15709.4]
  wire [5:0] _T_36441; // @[Mux.scala 31:69:@15710.4]
  wire [5:0] _T_36442; // @[Mux.scala 31:69:@15711.4]
  wire [5:0] _T_36443; // @[Mux.scala 31:69:@15712.4]
  wire [5:0] _T_36444; // @[Mux.scala 31:69:@15713.4]
  wire [5:0] _T_36445; // @[Mux.scala 31:69:@15714.4]
  wire [5:0] _T_36446; // @[Mux.scala 31:69:@15715.4]
  wire [5:0] _T_36447; // @[Mux.scala 31:69:@15716.4]
  wire [5:0] _T_36448; // @[Mux.scala 31:69:@15717.4]
  wire [5:0] _T_36449; // @[Mux.scala 31:69:@15718.4]
  wire [5:0] _T_36450; // @[Mux.scala 31:69:@15719.4]
  wire [5:0] select_48; // @[Mux.scala 31:69:@15720.4]
  wire [47:0] _GEN_3073; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3074; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3075; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3076; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3077; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3078; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3079; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3080; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3081; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3082; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3083; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3084; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3085; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3086; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3087; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3088; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3089; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3090; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3091; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3092; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3093; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3094; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3095; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3096; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3097; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3098; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3099; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3100; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3101; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3102; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3103; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3104; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3105; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3106; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3107; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3108; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3109; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3110; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3111; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3112; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3113; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3114; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3115; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3116; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3117; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3118; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3119; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3120; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3121; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3122; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3123; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3124; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3125; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3126; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3127; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3128; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3129; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3130; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3131; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3132; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3133; // @[Switch.scala 33:19:@15722.4]
  wire [47:0] _GEN_3134; // @[Switch.scala 33:19:@15722.4]
  wire [7:0] _T_36459; // @[Switch.scala 34:32:@15729.4]
  wire [15:0] _T_36467; // @[Switch.scala 34:32:@15737.4]
  wire [7:0] _T_36474; // @[Switch.scala 34:32:@15744.4]
  wire [31:0] _T_36483; // @[Switch.scala 34:32:@15753.4]
  wire [7:0] _T_36490; // @[Switch.scala 34:32:@15760.4]
  wire [15:0] _T_36498; // @[Switch.scala 34:32:@15768.4]
  wire [7:0] _T_36505; // @[Switch.scala 34:32:@15775.4]
  wire [31:0] _T_36514; // @[Switch.scala 34:32:@15784.4]
  wire [63:0] _T_36515; // @[Switch.scala 34:32:@15785.4]
  wire  _T_36519; // @[Switch.scala 30:53:@15788.4]
  wire  valid_49_0; // @[Switch.scala 30:36:@15789.4]
  wire  _T_36522; // @[Switch.scala 30:53:@15791.4]
  wire  valid_49_1; // @[Switch.scala 30:36:@15792.4]
  wire  _T_36525; // @[Switch.scala 30:53:@15794.4]
  wire  valid_49_2; // @[Switch.scala 30:36:@15795.4]
  wire  _T_36528; // @[Switch.scala 30:53:@15797.4]
  wire  valid_49_3; // @[Switch.scala 30:36:@15798.4]
  wire  _T_36531; // @[Switch.scala 30:53:@15800.4]
  wire  valid_49_4; // @[Switch.scala 30:36:@15801.4]
  wire  _T_36534; // @[Switch.scala 30:53:@15803.4]
  wire  valid_49_5; // @[Switch.scala 30:36:@15804.4]
  wire  _T_36537; // @[Switch.scala 30:53:@15806.4]
  wire  valid_49_6; // @[Switch.scala 30:36:@15807.4]
  wire  _T_36540; // @[Switch.scala 30:53:@15809.4]
  wire  valid_49_7; // @[Switch.scala 30:36:@15810.4]
  wire  _T_36543; // @[Switch.scala 30:53:@15812.4]
  wire  valid_49_8; // @[Switch.scala 30:36:@15813.4]
  wire  _T_36546; // @[Switch.scala 30:53:@15815.4]
  wire  valid_49_9; // @[Switch.scala 30:36:@15816.4]
  wire  _T_36549; // @[Switch.scala 30:53:@15818.4]
  wire  valid_49_10; // @[Switch.scala 30:36:@15819.4]
  wire  _T_36552; // @[Switch.scala 30:53:@15821.4]
  wire  valid_49_11; // @[Switch.scala 30:36:@15822.4]
  wire  _T_36555; // @[Switch.scala 30:53:@15824.4]
  wire  valid_49_12; // @[Switch.scala 30:36:@15825.4]
  wire  _T_36558; // @[Switch.scala 30:53:@15827.4]
  wire  valid_49_13; // @[Switch.scala 30:36:@15828.4]
  wire  _T_36561; // @[Switch.scala 30:53:@15830.4]
  wire  valid_49_14; // @[Switch.scala 30:36:@15831.4]
  wire  _T_36564; // @[Switch.scala 30:53:@15833.4]
  wire  valid_49_15; // @[Switch.scala 30:36:@15834.4]
  wire  _T_36567; // @[Switch.scala 30:53:@15836.4]
  wire  valid_49_16; // @[Switch.scala 30:36:@15837.4]
  wire  _T_36570; // @[Switch.scala 30:53:@15839.4]
  wire  valid_49_17; // @[Switch.scala 30:36:@15840.4]
  wire  _T_36573; // @[Switch.scala 30:53:@15842.4]
  wire  valid_49_18; // @[Switch.scala 30:36:@15843.4]
  wire  _T_36576; // @[Switch.scala 30:53:@15845.4]
  wire  valid_49_19; // @[Switch.scala 30:36:@15846.4]
  wire  _T_36579; // @[Switch.scala 30:53:@15848.4]
  wire  valid_49_20; // @[Switch.scala 30:36:@15849.4]
  wire  _T_36582; // @[Switch.scala 30:53:@15851.4]
  wire  valid_49_21; // @[Switch.scala 30:36:@15852.4]
  wire  _T_36585; // @[Switch.scala 30:53:@15854.4]
  wire  valid_49_22; // @[Switch.scala 30:36:@15855.4]
  wire  _T_36588; // @[Switch.scala 30:53:@15857.4]
  wire  valid_49_23; // @[Switch.scala 30:36:@15858.4]
  wire  _T_36591; // @[Switch.scala 30:53:@15860.4]
  wire  valid_49_24; // @[Switch.scala 30:36:@15861.4]
  wire  _T_36594; // @[Switch.scala 30:53:@15863.4]
  wire  valid_49_25; // @[Switch.scala 30:36:@15864.4]
  wire  _T_36597; // @[Switch.scala 30:53:@15866.4]
  wire  valid_49_26; // @[Switch.scala 30:36:@15867.4]
  wire  _T_36600; // @[Switch.scala 30:53:@15869.4]
  wire  valid_49_27; // @[Switch.scala 30:36:@15870.4]
  wire  _T_36603; // @[Switch.scala 30:53:@15872.4]
  wire  valid_49_28; // @[Switch.scala 30:36:@15873.4]
  wire  _T_36606; // @[Switch.scala 30:53:@15875.4]
  wire  valid_49_29; // @[Switch.scala 30:36:@15876.4]
  wire  _T_36609; // @[Switch.scala 30:53:@15878.4]
  wire  valid_49_30; // @[Switch.scala 30:36:@15879.4]
  wire  _T_36612; // @[Switch.scala 30:53:@15881.4]
  wire  valid_49_31; // @[Switch.scala 30:36:@15882.4]
  wire  _T_36615; // @[Switch.scala 30:53:@15884.4]
  wire  valid_49_32; // @[Switch.scala 30:36:@15885.4]
  wire  _T_36618; // @[Switch.scala 30:53:@15887.4]
  wire  valid_49_33; // @[Switch.scala 30:36:@15888.4]
  wire  _T_36621; // @[Switch.scala 30:53:@15890.4]
  wire  valid_49_34; // @[Switch.scala 30:36:@15891.4]
  wire  _T_36624; // @[Switch.scala 30:53:@15893.4]
  wire  valid_49_35; // @[Switch.scala 30:36:@15894.4]
  wire  _T_36627; // @[Switch.scala 30:53:@15896.4]
  wire  valid_49_36; // @[Switch.scala 30:36:@15897.4]
  wire  _T_36630; // @[Switch.scala 30:53:@15899.4]
  wire  valid_49_37; // @[Switch.scala 30:36:@15900.4]
  wire  _T_36633; // @[Switch.scala 30:53:@15902.4]
  wire  valid_49_38; // @[Switch.scala 30:36:@15903.4]
  wire  _T_36636; // @[Switch.scala 30:53:@15905.4]
  wire  valid_49_39; // @[Switch.scala 30:36:@15906.4]
  wire  _T_36639; // @[Switch.scala 30:53:@15908.4]
  wire  valid_49_40; // @[Switch.scala 30:36:@15909.4]
  wire  _T_36642; // @[Switch.scala 30:53:@15911.4]
  wire  valid_49_41; // @[Switch.scala 30:36:@15912.4]
  wire  _T_36645; // @[Switch.scala 30:53:@15914.4]
  wire  valid_49_42; // @[Switch.scala 30:36:@15915.4]
  wire  _T_36648; // @[Switch.scala 30:53:@15917.4]
  wire  valid_49_43; // @[Switch.scala 30:36:@15918.4]
  wire  _T_36651; // @[Switch.scala 30:53:@15920.4]
  wire  valid_49_44; // @[Switch.scala 30:36:@15921.4]
  wire  _T_36654; // @[Switch.scala 30:53:@15923.4]
  wire  valid_49_45; // @[Switch.scala 30:36:@15924.4]
  wire  _T_36657; // @[Switch.scala 30:53:@15926.4]
  wire  valid_49_46; // @[Switch.scala 30:36:@15927.4]
  wire  _T_36660; // @[Switch.scala 30:53:@15929.4]
  wire  valid_49_47; // @[Switch.scala 30:36:@15930.4]
  wire  _T_36663; // @[Switch.scala 30:53:@15932.4]
  wire  valid_49_48; // @[Switch.scala 30:36:@15933.4]
  wire  _T_36666; // @[Switch.scala 30:53:@15935.4]
  wire  valid_49_49; // @[Switch.scala 30:36:@15936.4]
  wire  _T_36669; // @[Switch.scala 30:53:@15938.4]
  wire  valid_49_50; // @[Switch.scala 30:36:@15939.4]
  wire  _T_36672; // @[Switch.scala 30:53:@15941.4]
  wire  valid_49_51; // @[Switch.scala 30:36:@15942.4]
  wire  _T_36675; // @[Switch.scala 30:53:@15944.4]
  wire  valid_49_52; // @[Switch.scala 30:36:@15945.4]
  wire  _T_36678; // @[Switch.scala 30:53:@15947.4]
  wire  valid_49_53; // @[Switch.scala 30:36:@15948.4]
  wire  _T_36681; // @[Switch.scala 30:53:@15950.4]
  wire  valid_49_54; // @[Switch.scala 30:36:@15951.4]
  wire  _T_36684; // @[Switch.scala 30:53:@15953.4]
  wire  valid_49_55; // @[Switch.scala 30:36:@15954.4]
  wire  _T_36687; // @[Switch.scala 30:53:@15956.4]
  wire  valid_49_56; // @[Switch.scala 30:36:@15957.4]
  wire  _T_36690; // @[Switch.scala 30:53:@15959.4]
  wire  valid_49_57; // @[Switch.scala 30:36:@15960.4]
  wire  _T_36693; // @[Switch.scala 30:53:@15962.4]
  wire  valid_49_58; // @[Switch.scala 30:36:@15963.4]
  wire  _T_36696; // @[Switch.scala 30:53:@15965.4]
  wire  valid_49_59; // @[Switch.scala 30:36:@15966.4]
  wire  _T_36699; // @[Switch.scala 30:53:@15968.4]
  wire  valid_49_60; // @[Switch.scala 30:36:@15969.4]
  wire  _T_36702; // @[Switch.scala 30:53:@15971.4]
  wire  valid_49_61; // @[Switch.scala 30:36:@15972.4]
  wire  _T_36705; // @[Switch.scala 30:53:@15974.4]
  wire  valid_49_62; // @[Switch.scala 30:36:@15975.4]
  wire  _T_36708; // @[Switch.scala 30:53:@15977.4]
  wire  valid_49_63; // @[Switch.scala 30:36:@15978.4]
  wire [5:0] _T_36774; // @[Mux.scala 31:69:@15980.4]
  wire [5:0] _T_36775; // @[Mux.scala 31:69:@15981.4]
  wire [5:0] _T_36776; // @[Mux.scala 31:69:@15982.4]
  wire [5:0] _T_36777; // @[Mux.scala 31:69:@15983.4]
  wire [5:0] _T_36778; // @[Mux.scala 31:69:@15984.4]
  wire [5:0] _T_36779; // @[Mux.scala 31:69:@15985.4]
  wire [5:0] _T_36780; // @[Mux.scala 31:69:@15986.4]
  wire [5:0] _T_36781; // @[Mux.scala 31:69:@15987.4]
  wire [5:0] _T_36782; // @[Mux.scala 31:69:@15988.4]
  wire [5:0] _T_36783; // @[Mux.scala 31:69:@15989.4]
  wire [5:0] _T_36784; // @[Mux.scala 31:69:@15990.4]
  wire [5:0] _T_36785; // @[Mux.scala 31:69:@15991.4]
  wire [5:0] _T_36786; // @[Mux.scala 31:69:@15992.4]
  wire [5:0] _T_36787; // @[Mux.scala 31:69:@15993.4]
  wire [5:0] _T_36788; // @[Mux.scala 31:69:@15994.4]
  wire [5:0] _T_36789; // @[Mux.scala 31:69:@15995.4]
  wire [5:0] _T_36790; // @[Mux.scala 31:69:@15996.4]
  wire [5:0] _T_36791; // @[Mux.scala 31:69:@15997.4]
  wire [5:0] _T_36792; // @[Mux.scala 31:69:@15998.4]
  wire [5:0] _T_36793; // @[Mux.scala 31:69:@15999.4]
  wire [5:0] _T_36794; // @[Mux.scala 31:69:@16000.4]
  wire [5:0] _T_36795; // @[Mux.scala 31:69:@16001.4]
  wire [5:0] _T_36796; // @[Mux.scala 31:69:@16002.4]
  wire [5:0] _T_36797; // @[Mux.scala 31:69:@16003.4]
  wire [5:0] _T_36798; // @[Mux.scala 31:69:@16004.4]
  wire [5:0] _T_36799; // @[Mux.scala 31:69:@16005.4]
  wire [5:0] _T_36800; // @[Mux.scala 31:69:@16006.4]
  wire [5:0] _T_36801; // @[Mux.scala 31:69:@16007.4]
  wire [5:0] _T_36802; // @[Mux.scala 31:69:@16008.4]
  wire [5:0] _T_36803; // @[Mux.scala 31:69:@16009.4]
  wire [5:0] _T_36804; // @[Mux.scala 31:69:@16010.4]
  wire [5:0] _T_36805; // @[Mux.scala 31:69:@16011.4]
  wire [5:0] _T_36806; // @[Mux.scala 31:69:@16012.4]
  wire [5:0] _T_36807; // @[Mux.scala 31:69:@16013.4]
  wire [5:0] _T_36808; // @[Mux.scala 31:69:@16014.4]
  wire [5:0] _T_36809; // @[Mux.scala 31:69:@16015.4]
  wire [5:0] _T_36810; // @[Mux.scala 31:69:@16016.4]
  wire [5:0] _T_36811; // @[Mux.scala 31:69:@16017.4]
  wire [5:0] _T_36812; // @[Mux.scala 31:69:@16018.4]
  wire [5:0] _T_36813; // @[Mux.scala 31:69:@16019.4]
  wire [5:0] _T_36814; // @[Mux.scala 31:69:@16020.4]
  wire [5:0] _T_36815; // @[Mux.scala 31:69:@16021.4]
  wire [5:0] _T_36816; // @[Mux.scala 31:69:@16022.4]
  wire [5:0] _T_36817; // @[Mux.scala 31:69:@16023.4]
  wire [5:0] _T_36818; // @[Mux.scala 31:69:@16024.4]
  wire [5:0] _T_36819; // @[Mux.scala 31:69:@16025.4]
  wire [5:0] _T_36820; // @[Mux.scala 31:69:@16026.4]
  wire [5:0] _T_36821; // @[Mux.scala 31:69:@16027.4]
  wire [5:0] _T_36822; // @[Mux.scala 31:69:@16028.4]
  wire [5:0] _T_36823; // @[Mux.scala 31:69:@16029.4]
  wire [5:0] _T_36824; // @[Mux.scala 31:69:@16030.4]
  wire [5:0] _T_36825; // @[Mux.scala 31:69:@16031.4]
  wire [5:0] _T_36826; // @[Mux.scala 31:69:@16032.4]
  wire [5:0] _T_36827; // @[Mux.scala 31:69:@16033.4]
  wire [5:0] _T_36828; // @[Mux.scala 31:69:@16034.4]
  wire [5:0] _T_36829; // @[Mux.scala 31:69:@16035.4]
  wire [5:0] _T_36830; // @[Mux.scala 31:69:@16036.4]
  wire [5:0] _T_36831; // @[Mux.scala 31:69:@16037.4]
  wire [5:0] _T_36832; // @[Mux.scala 31:69:@16038.4]
  wire [5:0] _T_36833; // @[Mux.scala 31:69:@16039.4]
  wire [5:0] _T_36834; // @[Mux.scala 31:69:@16040.4]
  wire [5:0] _T_36835; // @[Mux.scala 31:69:@16041.4]
  wire [5:0] select_49; // @[Mux.scala 31:69:@16042.4]
  wire [47:0] _GEN_3137; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3138; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3139; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3140; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3141; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3142; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3143; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3144; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3145; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3146; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3147; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3148; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3149; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3150; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3151; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3152; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3153; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3154; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3155; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3156; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3157; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3158; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3159; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3160; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3161; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3162; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3163; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3164; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3165; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3166; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3167; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3168; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3169; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3170; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3171; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3172; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3173; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3174; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3175; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3176; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3177; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3178; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3179; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3180; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3181; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3182; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3183; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3184; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3185; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3186; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3187; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3188; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3189; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3190; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3191; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3192; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3193; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3194; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3195; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3196; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3197; // @[Switch.scala 33:19:@16044.4]
  wire [47:0] _GEN_3198; // @[Switch.scala 33:19:@16044.4]
  wire [7:0] _T_36844; // @[Switch.scala 34:32:@16051.4]
  wire [15:0] _T_36852; // @[Switch.scala 34:32:@16059.4]
  wire [7:0] _T_36859; // @[Switch.scala 34:32:@16066.4]
  wire [31:0] _T_36868; // @[Switch.scala 34:32:@16075.4]
  wire [7:0] _T_36875; // @[Switch.scala 34:32:@16082.4]
  wire [15:0] _T_36883; // @[Switch.scala 34:32:@16090.4]
  wire [7:0] _T_36890; // @[Switch.scala 34:32:@16097.4]
  wire [31:0] _T_36899; // @[Switch.scala 34:32:@16106.4]
  wire [63:0] _T_36900; // @[Switch.scala 34:32:@16107.4]
  wire  _T_36904; // @[Switch.scala 30:53:@16110.4]
  wire  valid_50_0; // @[Switch.scala 30:36:@16111.4]
  wire  _T_36907; // @[Switch.scala 30:53:@16113.4]
  wire  valid_50_1; // @[Switch.scala 30:36:@16114.4]
  wire  _T_36910; // @[Switch.scala 30:53:@16116.4]
  wire  valid_50_2; // @[Switch.scala 30:36:@16117.4]
  wire  _T_36913; // @[Switch.scala 30:53:@16119.4]
  wire  valid_50_3; // @[Switch.scala 30:36:@16120.4]
  wire  _T_36916; // @[Switch.scala 30:53:@16122.4]
  wire  valid_50_4; // @[Switch.scala 30:36:@16123.4]
  wire  _T_36919; // @[Switch.scala 30:53:@16125.4]
  wire  valid_50_5; // @[Switch.scala 30:36:@16126.4]
  wire  _T_36922; // @[Switch.scala 30:53:@16128.4]
  wire  valid_50_6; // @[Switch.scala 30:36:@16129.4]
  wire  _T_36925; // @[Switch.scala 30:53:@16131.4]
  wire  valid_50_7; // @[Switch.scala 30:36:@16132.4]
  wire  _T_36928; // @[Switch.scala 30:53:@16134.4]
  wire  valid_50_8; // @[Switch.scala 30:36:@16135.4]
  wire  _T_36931; // @[Switch.scala 30:53:@16137.4]
  wire  valid_50_9; // @[Switch.scala 30:36:@16138.4]
  wire  _T_36934; // @[Switch.scala 30:53:@16140.4]
  wire  valid_50_10; // @[Switch.scala 30:36:@16141.4]
  wire  _T_36937; // @[Switch.scala 30:53:@16143.4]
  wire  valid_50_11; // @[Switch.scala 30:36:@16144.4]
  wire  _T_36940; // @[Switch.scala 30:53:@16146.4]
  wire  valid_50_12; // @[Switch.scala 30:36:@16147.4]
  wire  _T_36943; // @[Switch.scala 30:53:@16149.4]
  wire  valid_50_13; // @[Switch.scala 30:36:@16150.4]
  wire  _T_36946; // @[Switch.scala 30:53:@16152.4]
  wire  valid_50_14; // @[Switch.scala 30:36:@16153.4]
  wire  _T_36949; // @[Switch.scala 30:53:@16155.4]
  wire  valid_50_15; // @[Switch.scala 30:36:@16156.4]
  wire  _T_36952; // @[Switch.scala 30:53:@16158.4]
  wire  valid_50_16; // @[Switch.scala 30:36:@16159.4]
  wire  _T_36955; // @[Switch.scala 30:53:@16161.4]
  wire  valid_50_17; // @[Switch.scala 30:36:@16162.4]
  wire  _T_36958; // @[Switch.scala 30:53:@16164.4]
  wire  valid_50_18; // @[Switch.scala 30:36:@16165.4]
  wire  _T_36961; // @[Switch.scala 30:53:@16167.4]
  wire  valid_50_19; // @[Switch.scala 30:36:@16168.4]
  wire  _T_36964; // @[Switch.scala 30:53:@16170.4]
  wire  valid_50_20; // @[Switch.scala 30:36:@16171.4]
  wire  _T_36967; // @[Switch.scala 30:53:@16173.4]
  wire  valid_50_21; // @[Switch.scala 30:36:@16174.4]
  wire  _T_36970; // @[Switch.scala 30:53:@16176.4]
  wire  valid_50_22; // @[Switch.scala 30:36:@16177.4]
  wire  _T_36973; // @[Switch.scala 30:53:@16179.4]
  wire  valid_50_23; // @[Switch.scala 30:36:@16180.4]
  wire  _T_36976; // @[Switch.scala 30:53:@16182.4]
  wire  valid_50_24; // @[Switch.scala 30:36:@16183.4]
  wire  _T_36979; // @[Switch.scala 30:53:@16185.4]
  wire  valid_50_25; // @[Switch.scala 30:36:@16186.4]
  wire  _T_36982; // @[Switch.scala 30:53:@16188.4]
  wire  valid_50_26; // @[Switch.scala 30:36:@16189.4]
  wire  _T_36985; // @[Switch.scala 30:53:@16191.4]
  wire  valid_50_27; // @[Switch.scala 30:36:@16192.4]
  wire  _T_36988; // @[Switch.scala 30:53:@16194.4]
  wire  valid_50_28; // @[Switch.scala 30:36:@16195.4]
  wire  _T_36991; // @[Switch.scala 30:53:@16197.4]
  wire  valid_50_29; // @[Switch.scala 30:36:@16198.4]
  wire  _T_36994; // @[Switch.scala 30:53:@16200.4]
  wire  valid_50_30; // @[Switch.scala 30:36:@16201.4]
  wire  _T_36997; // @[Switch.scala 30:53:@16203.4]
  wire  valid_50_31; // @[Switch.scala 30:36:@16204.4]
  wire  _T_37000; // @[Switch.scala 30:53:@16206.4]
  wire  valid_50_32; // @[Switch.scala 30:36:@16207.4]
  wire  _T_37003; // @[Switch.scala 30:53:@16209.4]
  wire  valid_50_33; // @[Switch.scala 30:36:@16210.4]
  wire  _T_37006; // @[Switch.scala 30:53:@16212.4]
  wire  valid_50_34; // @[Switch.scala 30:36:@16213.4]
  wire  _T_37009; // @[Switch.scala 30:53:@16215.4]
  wire  valid_50_35; // @[Switch.scala 30:36:@16216.4]
  wire  _T_37012; // @[Switch.scala 30:53:@16218.4]
  wire  valid_50_36; // @[Switch.scala 30:36:@16219.4]
  wire  _T_37015; // @[Switch.scala 30:53:@16221.4]
  wire  valid_50_37; // @[Switch.scala 30:36:@16222.4]
  wire  _T_37018; // @[Switch.scala 30:53:@16224.4]
  wire  valid_50_38; // @[Switch.scala 30:36:@16225.4]
  wire  _T_37021; // @[Switch.scala 30:53:@16227.4]
  wire  valid_50_39; // @[Switch.scala 30:36:@16228.4]
  wire  _T_37024; // @[Switch.scala 30:53:@16230.4]
  wire  valid_50_40; // @[Switch.scala 30:36:@16231.4]
  wire  _T_37027; // @[Switch.scala 30:53:@16233.4]
  wire  valid_50_41; // @[Switch.scala 30:36:@16234.4]
  wire  _T_37030; // @[Switch.scala 30:53:@16236.4]
  wire  valid_50_42; // @[Switch.scala 30:36:@16237.4]
  wire  _T_37033; // @[Switch.scala 30:53:@16239.4]
  wire  valid_50_43; // @[Switch.scala 30:36:@16240.4]
  wire  _T_37036; // @[Switch.scala 30:53:@16242.4]
  wire  valid_50_44; // @[Switch.scala 30:36:@16243.4]
  wire  _T_37039; // @[Switch.scala 30:53:@16245.4]
  wire  valid_50_45; // @[Switch.scala 30:36:@16246.4]
  wire  _T_37042; // @[Switch.scala 30:53:@16248.4]
  wire  valid_50_46; // @[Switch.scala 30:36:@16249.4]
  wire  _T_37045; // @[Switch.scala 30:53:@16251.4]
  wire  valid_50_47; // @[Switch.scala 30:36:@16252.4]
  wire  _T_37048; // @[Switch.scala 30:53:@16254.4]
  wire  valid_50_48; // @[Switch.scala 30:36:@16255.4]
  wire  _T_37051; // @[Switch.scala 30:53:@16257.4]
  wire  valid_50_49; // @[Switch.scala 30:36:@16258.4]
  wire  _T_37054; // @[Switch.scala 30:53:@16260.4]
  wire  valid_50_50; // @[Switch.scala 30:36:@16261.4]
  wire  _T_37057; // @[Switch.scala 30:53:@16263.4]
  wire  valid_50_51; // @[Switch.scala 30:36:@16264.4]
  wire  _T_37060; // @[Switch.scala 30:53:@16266.4]
  wire  valid_50_52; // @[Switch.scala 30:36:@16267.4]
  wire  _T_37063; // @[Switch.scala 30:53:@16269.4]
  wire  valid_50_53; // @[Switch.scala 30:36:@16270.4]
  wire  _T_37066; // @[Switch.scala 30:53:@16272.4]
  wire  valid_50_54; // @[Switch.scala 30:36:@16273.4]
  wire  _T_37069; // @[Switch.scala 30:53:@16275.4]
  wire  valid_50_55; // @[Switch.scala 30:36:@16276.4]
  wire  _T_37072; // @[Switch.scala 30:53:@16278.4]
  wire  valid_50_56; // @[Switch.scala 30:36:@16279.4]
  wire  _T_37075; // @[Switch.scala 30:53:@16281.4]
  wire  valid_50_57; // @[Switch.scala 30:36:@16282.4]
  wire  _T_37078; // @[Switch.scala 30:53:@16284.4]
  wire  valid_50_58; // @[Switch.scala 30:36:@16285.4]
  wire  _T_37081; // @[Switch.scala 30:53:@16287.4]
  wire  valid_50_59; // @[Switch.scala 30:36:@16288.4]
  wire  _T_37084; // @[Switch.scala 30:53:@16290.4]
  wire  valid_50_60; // @[Switch.scala 30:36:@16291.4]
  wire  _T_37087; // @[Switch.scala 30:53:@16293.4]
  wire  valid_50_61; // @[Switch.scala 30:36:@16294.4]
  wire  _T_37090; // @[Switch.scala 30:53:@16296.4]
  wire  valid_50_62; // @[Switch.scala 30:36:@16297.4]
  wire  _T_37093; // @[Switch.scala 30:53:@16299.4]
  wire  valid_50_63; // @[Switch.scala 30:36:@16300.4]
  wire [5:0] _T_37159; // @[Mux.scala 31:69:@16302.4]
  wire [5:0] _T_37160; // @[Mux.scala 31:69:@16303.4]
  wire [5:0] _T_37161; // @[Mux.scala 31:69:@16304.4]
  wire [5:0] _T_37162; // @[Mux.scala 31:69:@16305.4]
  wire [5:0] _T_37163; // @[Mux.scala 31:69:@16306.4]
  wire [5:0] _T_37164; // @[Mux.scala 31:69:@16307.4]
  wire [5:0] _T_37165; // @[Mux.scala 31:69:@16308.4]
  wire [5:0] _T_37166; // @[Mux.scala 31:69:@16309.4]
  wire [5:0] _T_37167; // @[Mux.scala 31:69:@16310.4]
  wire [5:0] _T_37168; // @[Mux.scala 31:69:@16311.4]
  wire [5:0] _T_37169; // @[Mux.scala 31:69:@16312.4]
  wire [5:0] _T_37170; // @[Mux.scala 31:69:@16313.4]
  wire [5:0] _T_37171; // @[Mux.scala 31:69:@16314.4]
  wire [5:0] _T_37172; // @[Mux.scala 31:69:@16315.4]
  wire [5:0] _T_37173; // @[Mux.scala 31:69:@16316.4]
  wire [5:0] _T_37174; // @[Mux.scala 31:69:@16317.4]
  wire [5:0] _T_37175; // @[Mux.scala 31:69:@16318.4]
  wire [5:0] _T_37176; // @[Mux.scala 31:69:@16319.4]
  wire [5:0] _T_37177; // @[Mux.scala 31:69:@16320.4]
  wire [5:0] _T_37178; // @[Mux.scala 31:69:@16321.4]
  wire [5:0] _T_37179; // @[Mux.scala 31:69:@16322.4]
  wire [5:0] _T_37180; // @[Mux.scala 31:69:@16323.4]
  wire [5:0] _T_37181; // @[Mux.scala 31:69:@16324.4]
  wire [5:0] _T_37182; // @[Mux.scala 31:69:@16325.4]
  wire [5:0] _T_37183; // @[Mux.scala 31:69:@16326.4]
  wire [5:0] _T_37184; // @[Mux.scala 31:69:@16327.4]
  wire [5:0] _T_37185; // @[Mux.scala 31:69:@16328.4]
  wire [5:0] _T_37186; // @[Mux.scala 31:69:@16329.4]
  wire [5:0] _T_37187; // @[Mux.scala 31:69:@16330.4]
  wire [5:0] _T_37188; // @[Mux.scala 31:69:@16331.4]
  wire [5:0] _T_37189; // @[Mux.scala 31:69:@16332.4]
  wire [5:0] _T_37190; // @[Mux.scala 31:69:@16333.4]
  wire [5:0] _T_37191; // @[Mux.scala 31:69:@16334.4]
  wire [5:0] _T_37192; // @[Mux.scala 31:69:@16335.4]
  wire [5:0] _T_37193; // @[Mux.scala 31:69:@16336.4]
  wire [5:0] _T_37194; // @[Mux.scala 31:69:@16337.4]
  wire [5:0] _T_37195; // @[Mux.scala 31:69:@16338.4]
  wire [5:0] _T_37196; // @[Mux.scala 31:69:@16339.4]
  wire [5:0] _T_37197; // @[Mux.scala 31:69:@16340.4]
  wire [5:0] _T_37198; // @[Mux.scala 31:69:@16341.4]
  wire [5:0] _T_37199; // @[Mux.scala 31:69:@16342.4]
  wire [5:0] _T_37200; // @[Mux.scala 31:69:@16343.4]
  wire [5:0] _T_37201; // @[Mux.scala 31:69:@16344.4]
  wire [5:0] _T_37202; // @[Mux.scala 31:69:@16345.4]
  wire [5:0] _T_37203; // @[Mux.scala 31:69:@16346.4]
  wire [5:0] _T_37204; // @[Mux.scala 31:69:@16347.4]
  wire [5:0] _T_37205; // @[Mux.scala 31:69:@16348.4]
  wire [5:0] _T_37206; // @[Mux.scala 31:69:@16349.4]
  wire [5:0] _T_37207; // @[Mux.scala 31:69:@16350.4]
  wire [5:0] _T_37208; // @[Mux.scala 31:69:@16351.4]
  wire [5:0] _T_37209; // @[Mux.scala 31:69:@16352.4]
  wire [5:0] _T_37210; // @[Mux.scala 31:69:@16353.4]
  wire [5:0] _T_37211; // @[Mux.scala 31:69:@16354.4]
  wire [5:0] _T_37212; // @[Mux.scala 31:69:@16355.4]
  wire [5:0] _T_37213; // @[Mux.scala 31:69:@16356.4]
  wire [5:0] _T_37214; // @[Mux.scala 31:69:@16357.4]
  wire [5:0] _T_37215; // @[Mux.scala 31:69:@16358.4]
  wire [5:0] _T_37216; // @[Mux.scala 31:69:@16359.4]
  wire [5:0] _T_37217; // @[Mux.scala 31:69:@16360.4]
  wire [5:0] _T_37218; // @[Mux.scala 31:69:@16361.4]
  wire [5:0] _T_37219; // @[Mux.scala 31:69:@16362.4]
  wire [5:0] _T_37220; // @[Mux.scala 31:69:@16363.4]
  wire [5:0] select_50; // @[Mux.scala 31:69:@16364.4]
  wire [47:0] _GEN_3201; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3202; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3203; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3204; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3205; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3206; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3207; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3208; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3209; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3210; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3211; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3212; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3213; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3214; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3215; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3216; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3217; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3218; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3219; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3220; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3221; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3222; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3223; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3224; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3225; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3226; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3227; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3228; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3229; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3230; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3231; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3232; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3233; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3234; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3235; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3236; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3237; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3238; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3239; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3240; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3241; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3242; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3243; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3244; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3245; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3246; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3247; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3248; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3249; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3250; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3251; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3252; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3253; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3254; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3255; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3256; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3257; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3258; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3259; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3260; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3261; // @[Switch.scala 33:19:@16366.4]
  wire [47:0] _GEN_3262; // @[Switch.scala 33:19:@16366.4]
  wire [7:0] _T_37229; // @[Switch.scala 34:32:@16373.4]
  wire [15:0] _T_37237; // @[Switch.scala 34:32:@16381.4]
  wire [7:0] _T_37244; // @[Switch.scala 34:32:@16388.4]
  wire [31:0] _T_37253; // @[Switch.scala 34:32:@16397.4]
  wire [7:0] _T_37260; // @[Switch.scala 34:32:@16404.4]
  wire [15:0] _T_37268; // @[Switch.scala 34:32:@16412.4]
  wire [7:0] _T_37275; // @[Switch.scala 34:32:@16419.4]
  wire [31:0] _T_37284; // @[Switch.scala 34:32:@16428.4]
  wire [63:0] _T_37285; // @[Switch.scala 34:32:@16429.4]
  wire  _T_37289; // @[Switch.scala 30:53:@16432.4]
  wire  valid_51_0; // @[Switch.scala 30:36:@16433.4]
  wire  _T_37292; // @[Switch.scala 30:53:@16435.4]
  wire  valid_51_1; // @[Switch.scala 30:36:@16436.4]
  wire  _T_37295; // @[Switch.scala 30:53:@16438.4]
  wire  valid_51_2; // @[Switch.scala 30:36:@16439.4]
  wire  _T_37298; // @[Switch.scala 30:53:@16441.4]
  wire  valid_51_3; // @[Switch.scala 30:36:@16442.4]
  wire  _T_37301; // @[Switch.scala 30:53:@16444.4]
  wire  valid_51_4; // @[Switch.scala 30:36:@16445.4]
  wire  _T_37304; // @[Switch.scala 30:53:@16447.4]
  wire  valid_51_5; // @[Switch.scala 30:36:@16448.4]
  wire  _T_37307; // @[Switch.scala 30:53:@16450.4]
  wire  valid_51_6; // @[Switch.scala 30:36:@16451.4]
  wire  _T_37310; // @[Switch.scala 30:53:@16453.4]
  wire  valid_51_7; // @[Switch.scala 30:36:@16454.4]
  wire  _T_37313; // @[Switch.scala 30:53:@16456.4]
  wire  valid_51_8; // @[Switch.scala 30:36:@16457.4]
  wire  _T_37316; // @[Switch.scala 30:53:@16459.4]
  wire  valid_51_9; // @[Switch.scala 30:36:@16460.4]
  wire  _T_37319; // @[Switch.scala 30:53:@16462.4]
  wire  valid_51_10; // @[Switch.scala 30:36:@16463.4]
  wire  _T_37322; // @[Switch.scala 30:53:@16465.4]
  wire  valid_51_11; // @[Switch.scala 30:36:@16466.4]
  wire  _T_37325; // @[Switch.scala 30:53:@16468.4]
  wire  valid_51_12; // @[Switch.scala 30:36:@16469.4]
  wire  _T_37328; // @[Switch.scala 30:53:@16471.4]
  wire  valid_51_13; // @[Switch.scala 30:36:@16472.4]
  wire  _T_37331; // @[Switch.scala 30:53:@16474.4]
  wire  valid_51_14; // @[Switch.scala 30:36:@16475.4]
  wire  _T_37334; // @[Switch.scala 30:53:@16477.4]
  wire  valid_51_15; // @[Switch.scala 30:36:@16478.4]
  wire  _T_37337; // @[Switch.scala 30:53:@16480.4]
  wire  valid_51_16; // @[Switch.scala 30:36:@16481.4]
  wire  _T_37340; // @[Switch.scala 30:53:@16483.4]
  wire  valid_51_17; // @[Switch.scala 30:36:@16484.4]
  wire  _T_37343; // @[Switch.scala 30:53:@16486.4]
  wire  valid_51_18; // @[Switch.scala 30:36:@16487.4]
  wire  _T_37346; // @[Switch.scala 30:53:@16489.4]
  wire  valid_51_19; // @[Switch.scala 30:36:@16490.4]
  wire  _T_37349; // @[Switch.scala 30:53:@16492.4]
  wire  valid_51_20; // @[Switch.scala 30:36:@16493.4]
  wire  _T_37352; // @[Switch.scala 30:53:@16495.4]
  wire  valid_51_21; // @[Switch.scala 30:36:@16496.4]
  wire  _T_37355; // @[Switch.scala 30:53:@16498.4]
  wire  valid_51_22; // @[Switch.scala 30:36:@16499.4]
  wire  _T_37358; // @[Switch.scala 30:53:@16501.4]
  wire  valid_51_23; // @[Switch.scala 30:36:@16502.4]
  wire  _T_37361; // @[Switch.scala 30:53:@16504.4]
  wire  valid_51_24; // @[Switch.scala 30:36:@16505.4]
  wire  _T_37364; // @[Switch.scala 30:53:@16507.4]
  wire  valid_51_25; // @[Switch.scala 30:36:@16508.4]
  wire  _T_37367; // @[Switch.scala 30:53:@16510.4]
  wire  valid_51_26; // @[Switch.scala 30:36:@16511.4]
  wire  _T_37370; // @[Switch.scala 30:53:@16513.4]
  wire  valid_51_27; // @[Switch.scala 30:36:@16514.4]
  wire  _T_37373; // @[Switch.scala 30:53:@16516.4]
  wire  valid_51_28; // @[Switch.scala 30:36:@16517.4]
  wire  _T_37376; // @[Switch.scala 30:53:@16519.4]
  wire  valid_51_29; // @[Switch.scala 30:36:@16520.4]
  wire  _T_37379; // @[Switch.scala 30:53:@16522.4]
  wire  valid_51_30; // @[Switch.scala 30:36:@16523.4]
  wire  _T_37382; // @[Switch.scala 30:53:@16525.4]
  wire  valid_51_31; // @[Switch.scala 30:36:@16526.4]
  wire  _T_37385; // @[Switch.scala 30:53:@16528.4]
  wire  valid_51_32; // @[Switch.scala 30:36:@16529.4]
  wire  _T_37388; // @[Switch.scala 30:53:@16531.4]
  wire  valid_51_33; // @[Switch.scala 30:36:@16532.4]
  wire  _T_37391; // @[Switch.scala 30:53:@16534.4]
  wire  valid_51_34; // @[Switch.scala 30:36:@16535.4]
  wire  _T_37394; // @[Switch.scala 30:53:@16537.4]
  wire  valid_51_35; // @[Switch.scala 30:36:@16538.4]
  wire  _T_37397; // @[Switch.scala 30:53:@16540.4]
  wire  valid_51_36; // @[Switch.scala 30:36:@16541.4]
  wire  _T_37400; // @[Switch.scala 30:53:@16543.4]
  wire  valid_51_37; // @[Switch.scala 30:36:@16544.4]
  wire  _T_37403; // @[Switch.scala 30:53:@16546.4]
  wire  valid_51_38; // @[Switch.scala 30:36:@16547.4]
  wire  _T_37406; // @[Switch.scala 30:53:@16549.4]
  wire  valid_51_39; // @[Switch.scala 30:36:@16550.4]
  wire  _T_37409; // @[Switch.scala 30:53:@16552.4]
  wire  valid_51_40; // @[Switch.scala 30:36:@16553.4]
  wire  _T_37412; // @[Switch.scala 30:53:@16555.4]
  wire  valid_51_41; // @[Switch.scala 30:36:@16556.4]
  wire  _T_37415; // @[Switch.scala 30:53:@16558.4]
  wire  valid_51_42; // @[Switch.scala 30:36:@16559.4]
  wire  _T_37418; // @[Switch.scala 30:53:@16561.4]
  wire  valid_51_43; // @[Switch.scala 30:36:@16562.4]
  wire  _T_37421; // @[Switch.scala 30:53:@16564.4]
  wire  valid_51_44; // @[Switch.scala 30:36:@16565.4]
  wire  _T_37424; // @[Switch.scala 30:53:@16567.4]
  wire  valid_51_45; // @[Switch.scala 30:36:@16568.4]
  wire  _T_37427; // @[Switch.scala 30:53:@16570.4]
  wire  valid_51_46; // @[Switch.scala 30:36:@16571.4]
  wire  _T_37430; // @[Switch.scala 30:53:@16573.4]
  wire  valid_51_47; // @[Switch.scala 30:36:@16574.4]
  wire  _T_37433; // @[Switch.scala 30:53:@16576.4]
  wire  valid_51_48; // @[Switch.scala 30:36:@16577.4]
  wire  _T_37436; // @[Switch.scala 30:53:@16579.4]
  wire  valid_51_49; // @[Switch.scala 30:36:@16580.4]
  wire  _T_37439; // @[Switch.scala 30:53:@16582.4]
  wire  valid_51_50; // @[Switch.scala 30:36:@16583.4]
  wire  _T_37442; // @[Switch.scala 30:53:@16585.4]
  wire  valid_51_51; // @[Switch.scala 30:36:@16586.4]
  wire  _T_37445; // @[Switch.scala 30:53:@16588.4]
  wire  valid_51_52; // @[Switch.scala 30:36:@16589.4]
  wire  _T_37448; // @[Switch.scala 30:53:@16591.4]
  wire  valid_51_53; // @[Switch.scala 30:36:@16592.4]
  wire  _T_37451; // @[Switch.scala 30:53:@16594.4]
  wire  valid_51_54; // @[Switch.scala 30:36:@16595.4]
  wire  _T_37454; // @[Switch.scala 30:53:@16597.4]
  wire  valid_51_55; // @[Switch.scala 30:36:@16598.4]
  wire  _T_37457; // @[Switch.scala 30:53:@16600.4]
  wire  valid_51_56; // @[Switch.scala 30:36:@16601.4]
  wire  _T_37460; // @[Switch.scala 30:53:@16603.4]
  wire  valid_51_57; // @[Switch.scala 30:36:@16604.4]
  wire  _T_37463; // @[Switch.scala 30:53:@16606.4]
  wire  valid_51_58; // @[Switch.scala 30:36:@16607.4]
  wire  _T_37466; // @[Switch.scala 30:53:@16609.4]
  wire  valid_51_59; // @[Switch.scala 30:36:@16610.4]
  wire  _T_37469; // @[Switch.scala 30:53:@16612.4]
  wire  valid_51_60; // @[Switch.scala 30:36:@16613.4]
  wire  _T_37472; // @[Switch.scala 30:53:@16615.4]
  wire  valid_51_61; // @[Switch.scala 30:36:@16616.4]
  wire  _T_37475; // @[Switch.scala 30:53:@16618.4]
  wire  valid_51_62; // @[Switch.scala 30:36:@16619.4]
  wire  _T_37478; // @[Switch.scala 30:53:@16621.4]
  wire  valid_51_63; // @[Switch.scala 30:36:@16622.4]
  wire [5:0] _T_37544; // @[Mux.scala 31:69:@16624.4]
  wire [5:0] _T_37545; // @[Mux.scala 31:69:@16625.4]
  wire [5:0] _T_37546; // @[Mux.scala 31:69:@16626.4]
  wire [5:0] _T_37547; // @[Mux.scala 31:69:@16627.4]
  wire [5:0] _T_37548; // @[Mux.scala 31:69:@16628.4]
  wire [5:0] _T_37549; // @[Mux.scala 31:69:@16629.4]
  wire [5:0] _T_37550; // @[Mux.scala 31:69:@16630.4]
  wire [5:0] _T_37551; // @[Mux.scala 31:69:@16631.4]
  wire [5:0] _T_37552; // @[Mux.scala 31:69:@16632.4]
  wire [5:0] _T_37553; // @[Mux.scala 31:69:@16633.4]
  wire [5:0] _T_37554; // @[Mux.scala 31:69:@16634.4]
  wire [5:0] _T_37555; // @[Mux.scala 31:69:@16635.4]
  wire [5:0] _T_37556; // @[Mux.scala 31:69:@16636.4]
  wire [5:0] _T_37557; // @[Mux.scala 31:69:@16637.4]
  wire [5:0] _T_37558; // @[Mux.scala 31:69:@16638.4]
  wire [5:0] _T_37559; // @[Mux.scala 31:69:@16639.4]
  wire [5:0] _T_37560; // @[Mux.scala 31:69:@16640.4]
  wire [5:0] _T_37561; // @[Mux.scala 31:69:@16641.4]
  wire [5:0] _T_37562; // @[Mux.scala 31:69:@16642.4]
  wire [5:0] _T_37563; // @[Mux.scala 31:69:@16643.4]
  wire [5:0] _T_37564; // @[Mux.scala 31:69:@16644.4]
  wire [5:0] _T_37565; // @[Mux.scala 31:69:@16645.4]
  wire [5:0] _T_37566; // @[Mux.scala 31:69:@16646.4]
  wire [5:0] _T_37567; // @[Mux.scala 31:69:@16647.4]
  wire [5:0] _T_37568; // @[Mux.scala 31:69:@16648.4]
  wire [5:0] _T_37569; // @[Mux.scala 31:69:@16649.4]
  wire [5:0] _T_37570; // @[Mux.scala 31:69:@16650.4]
  wire [5:0] _T_37571; // @[Mux.scala 31:69:@16651.4]
  wire [5:0] _T_37572; // @[Mux.scala 31:69:@16652.4]
  wire [5:0] _T_37573; // @[Mux.scala 31:69:@16653.4]
  wire [5:0] _T_37574; // @[Mux.scala 31:69:@16654.4]
  wire [5:0] _T_37575; // @[Mux.scala 31:69:@16655.4]
  wire [5:0] _T_37576; // @[Mux.scala 31:69:@16656.4]
  wire [5:0] _T_37577; // @[Mux.scala 31:69:@16657.4]
  wire [5:0] _T_37578; // @[Mux.scala 31:69:@16658.4]
  wire [5:0] _T_37579; // @[Mux.scala 31:69:@16659.4]
  wire [5:0] _T_37580; // @[Mux.scala 31:69:@16660.4]
  wire [5:0] _T_37581; // @[Mux.scala 31:69:@16661.4]
  wire [5:0] _T_37582; // @[Mux.scala 31:69:@16662.4]
  wire [5:0] _T_37583; // @[Mux.scala 31:69:@16663.4]
  wire [5:0] _T_37584; // @[Mux.scala 31:69:@16664.4]
  wire [5:0] _T_37585; // @[Mux.scala 31:69:@16665.4]
  wire [5:0] _T_37586; // @[Mux.scala 31:69:@16666.4]
  wire [5:0] _T_37587; // @[Mux.scala 31:69:@16667.4]
  wire [5:0] _T_37588; // @[Mux.scala 31:69:@16668.4]
  wire [5:0] _T_37589; // @[Mux.scala 31:69:@16669.4]
  wire [5:0] _T_37590; // @[Mux.scala 31:69:@16670.4]
  wire [5:0] _T_37591; // @[Mux.scala 31:69:@16671.4]
  wire [5:0] _T_37592; // @[Mux.scala 31:69:@16672.4]
  wire [5:0] _T_37593; // @[Mux.scala 31:69:@16673.4]
  wire [5:0] _T_37594; // @[Mux.scala 31:69:@16674.4]
  wire [5:0] _T_37595; // @[Mux.scala 31:69:@16675.4]
  wire [5:0] _T_37596; // @[Mux.scala 31:69:@16676.4]
  wire [5:0] _T_37597; // @[Mux.scala 31:69:@16677.4]
  wire [5:0] _T_37598; // @[Mux.scala 31:69:@16678.4]
  wire [5:0] _T_37599; // @[Mux.scala 31:69:@16679.4]
  wire [5:0] _T_37600; // @[Mux.scala 31:69:@16680.4]
  wire [5:0] _T_37601; // @[Mux.scala 31:69:@16681.4]
  wire [5:0] _T_37602; // @[Mux.scala 31:69:@16682.4]
  wire [5:0] _T_37603; // @[Mux.scala 31:69:@16683.4]
  wire [5:0] _T_37604; // @[Mux.scala 31:69:@16684.4]
  wire [5:0] _T_37605; // @[Mux.scala 31:69:@16685.4]
  wire [5:0] select_51; // @[Mux.scala 31:69:@16686.4]
  wire [47:0] _GEN_3265; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3266; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3267; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3268; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3269; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3270; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3271; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3272; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3273; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3274; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3275; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3276; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3277; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3278; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3279; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3280; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3281; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3282; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3283; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3284; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3285; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3286; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3287; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3288; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3289; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3290; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3291; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3292; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3293; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3294; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3295; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3296; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3297; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3298; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3299; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3300; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3301; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3302; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3303; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3304; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3305; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3306; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3307; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3308; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3309; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3310; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3311; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3312; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3313; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3314; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3315; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3316; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3317; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3318; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3319; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3320; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3321; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3322; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3323; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3324; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3325; // @[Switch.scala 33:19:@16688.4]
  wire [47:0] _GEN_3326; // @[Switch.scala 33:19:@16688.4]
  wire [7:0] _T_37614; // @[Switch.scala 34:32:@16695.4]
  wire [15:0] _T_37622; // @[Switch.scala 34:32:@16703.4]
  wire [7:0] _T_37629; // @[Switch.scala 34:32:@16710.4]
  wire [31:0] _T_37638; // @[Switch.scala 34:32:@16719.4]
  wire [7:0] _T_37645; // @[Switch.scala 34:32:@16726.4]
  wire [15:0] _T_37653; // @[Switch.scala 34:32:@16734.4]
  wire [7:0] _T_37660; // @[Switch.scala 34:32:@16741.4]
  wire [31:0] _T_37669; // @[Switch.scala 34:32:@16750.4]
  wire [63:0] _T_37670; // @[Switch.scala 34:32:@16751.4]
  wire  _T_37674; // @[Switch.scala 30:53:@16754.4]
  wire  valid_52_0; // @[Switch.scala 30:36:@16755.4]
  wire  _T_37677; // @[Switch.scala 30:53:@16757.4]
  wire  valid_52_1; // @[Switch.scala 30:36:@16758.4]
  wire  _T_37680; // @[Switch.scala 30:53:@16760.4]
  wire  valid_52_2; // @[Switch.scala 30:36:@16761.4]
  wire  _T_37683; // @[Switch.scala 30:53:@16763.4]
  wire  valid_52_3; // @[Switch.scala 30:36:@16764.4]
  wire  _T_37686; // @[Switch.scala 30:53:@16766.4]
  wire  valid_52_4; // @[Switch.scala 30:36:@16767.4]
  wire  _T_37689; // @[Switch.scala 30:53:@16769.4]
  wire  valid_52_5; // @[Switch.scala 30:36:@16770.4]
  wire  _T_37692; // @[Switch.scala 30:53:@16772.4]
  wire  valid_52_6; // @[Switch.scala 30:36:@16773.4]
  wire  _T_37695; // @[Switch.scala 30:53:@16775.4]
  wire  valid_52_7; // @[Switch.scala 30:36:@16776.4]
  wire  _T_37698; // @[Switch.scala 30:53:@16778.4]
  wire  valid_52_8; // @[Switch.scala 30:36:@16779.4]
  wire  _T_37701; // @[Switch.scala 30:53:@16781.4]
  wire  valid_52_9; // @[Switch.scala 30:36:@16782.4]
  wire  _T_37704; // @[Switch.scala 30:53:@16784.4]
  wire  valid_52_10; // @[Switch.scala 30:36:@16785.4]
  wire  _T_37707; // @[Switch.scala 30:53:@16787.4]
  wire  valid_52_11; // @[Switch.scala 30:36:@16788.4]
  wire  _T_37710; // @[Switch.scala 30:53:@16790.4]
  wire  valid_52_12; // @[Switch.scala 30:36:@16791.4]
  wire  _T_37713; // @[Switch.scala 30:53:@16793.4]
  wire  valid_52_13; // @[Switch.scala 30:36:@16794.4]
  wire  _T_37716; // @[Switch.scala 30:53:@16796.4]
  wire  valid_52_14; // @[Switch.scala 30:36:@16797.4]
  wire  _T_37719; // @[Switch.scala 30:53:@16799.4]
  wire  valid_52_15; // @[Switch.scala 30:36:@16800.4]
  wire  _T_37722; // @[Switch.scala 30:53:@16802.4]
  wire  valid_52_16; // @[Switch.scala 30:36:@16803.4]
  wire  _T_37725; // @[Switch.scala 30:53:@16805.4]
  wire  valid_52_17; // @[Switch.scala 30:36:@16806.4]
  wire  _T_37728; // @[Switch.scala 30:53:@16808.4]
  wire  valid_52_18; // @[Switch.scala 30:36:@16809.4]
  wire  _T_37731; // @[Switch.scala 30:53:@16811.4]
  wire  valid_52_19; // @[Switch.scala 30:36:@16812.4]
  wire  _T_37734; // @[Switch.scala 30:53:@16814.4]
  wire  valid_52_20; // @[Switch.scala 30:36:@16815.4]
  wire  _T_37737; // @[Switch.scala 30:53:@16817.4]
  wire  valid_52_21; // @[Switch.scala 30:36:@16818.4]
  wire  _T_37740; // @[Switch.scala 30:53:@16820.4]
  wire  valid_52_22; // @[Switch.scala 30:36:@16821.4]
  wire  _T_37743; // @[Switch.scala 30:53:@16823.4]
  wire  valid_52_23; // @[Switch.scala 30:36:@16824.4]
  wire  _T_37746; // @[Switch.scala 30:53:@16826.4]
  wire  valid_52_24; // @[Switch.scala 30:36:@16827.4]
  wire  _T_37749; // @[Switch.scala 30:53:@16829.4]
  wire  valid_52_25; // @[Switch.scala 30:36:@16830.4]
  wire  _T_37752; // @[Switch.scala 30:53:@16832.4]
  wire  valid_52_26; // @[Switch.scala 30:36:@16833.4]
  wire  _T_37755; // @[Switch.scala 30:53:@16835.4]
  wire  valid_52_27; // @[Switch.scala 30:36:@16836.4]
  wire  _T_37758; // @[Switch.scala 30:53:@16838.4]
  wire  valid_52_28; // @[Switch.scala 30:36:@16839.4]
  wire  _T_37761; // @[Switch.scala 30:53:@16841.4]
  wire  valid_52_29; // @[Switch.scala 30:36:@16842.4]
  wire  _T_37764; // @[Switch.scala 30:53:@16844.4]
  wire  valid_52_30; // @[Switch.scala 30:36:@16845.4]
  wire  _T_37767; // @[Switch.scala 30:53:@16847.4]
  wire  valid_52_31; // @[Switch.scala 30:36:@16848.4]
  wire  _T_37770; // @[Switch.scala 30:53:@16850.4]
  wire  valid_52_32; // @[Switch.scala 30:36:@16851.4]
  wire  _T_37773; // @[Switch.scala 30:53:@16853.4]
  wire  valid_52_33; // @[Switch.scala 30:36:@16854.4]
  wire  _T_37776; // @[Switch.scala 30:53:@16856.4]
  wire  valid_52_34; // @[Switch.scala 30:36:@16857.4]
  wire  _T_37779; // @[Switch.scala 30:53:@16859.4]
  wire  valid_52_35; // @[Switch.scala 30:36:@16860.4]
  wire  _T_37782; // @[Switch.scala 30:53:@16862.4]
  wire  valid_52_36; // @[Switch.scala 30:36:@16863.4]
  wire  _T_37785; // @[Switch.scala 30:53:@16865.4]
  wire  valid_52_37; // @[Switch.scala 30:36:@16866.4]
  wire  _T_37788; // @[Switch.scala 30:53:@16868.4]
  wire  valid_52_38; // @[Switch.scala 30:36:@16869.4]
  wire  _T_37791; // @[Switch.scala 30:53:@16871.4]
  wire  valid_52_39; // @[Switch.scala 30:36:@16872.4]
  wire  _T_37794; // @[Switch.scala 30:53:@16874.4]
  wire  valid_52_40; // @[Switch.scala 30:36:@16875.4]
  wire  _T_37797; // @[Switch.scala 30:53:@16877.4]
  wire  valid_52_41; // @[Switch.scala 30:36:@16878.4]
  wire  _T_37800; // @[Switch.scala 30:53:@16880.4]
  wire  valid_52_42; // @[Switch.scala 30:36:@16881.4]
  wire  _T_37803; // @[Switch.scala 30:53:@16883.4]
  wire  valid_52_43; // @[Switch.scala 30:36:@16884.4]
  wire  _T_37806; // @[Switch.scala 30:53:@16886.4]
  wire  valid_52_44; // @[Switch.scala 30:36:@16887.4]
  wire  _T_37809; // @[Switch.scala 30:53:@16889.4]
  wire  valid_52_45; // @[Switch.scala 30:36:@16890.4]
  wire  _T_37812; // @[Switch.scala 30:53:@16892.4]
  wire  valid_52_46; // @[Switch.scala 30:36:@16893.4]
  wire  _T_37815; // @[Switch.scala 30:53:@16895.4]
  wire  valid_52_47; // @[Switch.scala 30:36:@16896.4]
  wire  _T_37818; // @[Switch.scala 30:53:@16898.4]
  wire  valid_52_48; // @[Switch.scala 30:36:@16899.4]
  wire  _T_37821; // @[Switch.scala 30:53:@16901.4]
  wire  valid_52_49; // @[Switch.scala 30:36:@16902.4]
  wire  _T_37824; // @[Switch.scala 30:53:@16904.4]
  wire  valid_52_50; // @[Switch.scala 30:36:@16905.4]
  wire  _T_37827; // @[Switch.scala 30:53:@16907.4]
  wire  valid_52_51; // @[Switch.scala 30:36:@16908.4]
  wire  _T_37830; // @[Switch.scala 30:53:@16910.4]
  wire  valid_52_52; // @[Switch.scala 30:36:@16911.4]
  wire  _T_37833; // @[Switch.scala 30:53:@16913.4]
  wire  valid_52_53; // @[Switch.scala 30:36:@16914.4]
  wire  _T_37836; // @[Switch.scala 30:53:@16916.4]
  wire  valid_52_54; // @[Switch.scala 30:36:@16917.4]
  wire  _T_37839; // @[Switch.scala 30:53:@16919.4]
  wire  valid_52_55; // @[Switch.scala 30:36:@16920.4]
  wire  _T_37842; // @[Switch.scala 30:53:@16922.4]
  wire  valid_52_56; // @[Switch.scala 30:36:@16923.4]
  wire  _T_37845; // @[Switch.scala 30:53:@16925.4]
  wire  valid_52_57; // @[Switch.scala 30:36:@16926.4]
  wire  _T_37848; // @[Switch.scala 30:53:@16928.4]
  wire  valid_52_58; // @[Switch.scala 30:36:@16929.4]
  wire  _T_37851; // @[Switch.scala 30:53:@16931.4]
  wire  valid_52_59; // @[Switch.scala 30:36:@16932.4]
  wire  _T_37854; // @[Switch.scala 30:53:@16934.4]
  wire  valid_52_60; // @[Switch.scala 30:36:@16935.4]
  wire  _T_37857; // @[Switch.scala 30:53:@16937.4]
  wire  valid_52_61; // @[Switch.scala 30:36:@16938.4]
  wire  _T_37860; // @[Switch.scala 30:53:@16940.4]
  wire  valid_52_62; // @[Switch.scala 30:36:@16941.4]
  wire  _T_37863; // @[Switch.scala 30:53:@16943.4]
  wire  valid_52_63; // @[Switch.scala 30:36:@16944.4]
  wire [5:0] _T_37929; // @[Mux.scala 31:69:@16946.4]
  wire [5:0] _T_37930; // @[Mux.scala 31:69:@16947.4]
  wire [5:0] _T_37931; // @[Mux.scala 31:69:@16948.4]
  wire [5:0] _T_37932; // @[Mux.scala 31:69:@16949.4]
  wire [5:0] _T_37933; // @[Mux.scala 31:69:@16950.4]
  wire [5:0] _T_37934; // @[Mux.scala 31:69:@16951.4]
  wire [5:0] _T_37935; // @[Mux.scala 31:69:@16952.4]
  wire [5:0] _T_37936; // @[Mux.scala 31:69:@16953.4]
  wire [5:0] _T_37937; // @[Mux.scala 31:69:@16954.4]
  wire [5:0] _T_37938; // @[Mux.scala 31:69:@16955.4]
  wire [5:0] _T_37939; // @[Mux.scala 31:69:@16956.4]
  wire [5:0] _T_37940; // @[Mux.scala 31:69:@16957.4]
  wire [5:0] _T_37941; // @[Mux.scala 31:69:@16958.4]
  wire [5:0] _T_37942; // @[Mux.scala 31:69:@16959.4]
  wire [5:0] _T_37943; // @[Mux.scala 31:69:@16960.4]
  wire [5:0] _T_37944; // @[Mux.scala 31:69:@16961.4]
  wire [5:0] _T_37945; // @[Mux.scala 31:69:@16962.4]
  wire [5:0] _T_37946; // @[Mux.scala 31:69:@16963.4]
  wire [5:0] _T_37947; // @[Mux.scala 31:69:@16964.4]
  wire [5:0] _T_37948; // @[Mux.scala 31:69:@16965.4]
  wire [5:0] _T_37949; // @[Mux.scala 31:69:@16966.4]
  wire [5:0] _T_37950; // @[Mux.scala 31:69:@16967.4]
  wire [5:0] _T_37951; // @[Mux.scala 31:69:@16968.4]
  wire [5:0] _T_37952; // @[Mux.scala 31:69:@16969.4]
  wire [5:0] _T_37953; // @[Mux.scala 31:69:@16970.4]
  wire [5:0] _T_37954; // @[Mux.scala 31:69:@16971.4]
  wire [5:0] _T_37955; // @[Mux.scala 31:69:@16972.4]
  wire [5:0] _T_37956; // @[Mux.scala 31:69:@16973.4]
  wire [5:0] _T_37957; // @[Mux.scala 31:69:@16974.4]
  wire [5:0] _T_37958; // @[Mux.scala 31:69:@16975.4]
  wire [5:0] _T_37959; // @[Mux.scala 31:69:@16976.4]
  wire [5:0] _T_37960; // @[Mux.scala 31:69:@16977.4]
  wire [5:0] _T_37961; // @[Mux.scala 31:69:@16978.4]
  wire [5:0] _T_37962; // @[Mux.scala 31:69:@16979.4]
  wire [5:0] _T_37963; // @[Mux.scala 31:69:@16980.4]
  wire [5:0] _T_37964; // @[Mux.scala 31:69:@16981.4]
  wire [5:0] _T_37965; // @[Mux.scala 31:69:@16982.4]
  wire [5:0] _T_37966; // @[Mux.scala 31:69:@16983.4]
  wire [5:0] _T_37967; // @[Mux.scala 31:69:@16984.4]
  wire [5:0] _T_37968; // @[Mux.scala 31:69:@16985.4]
  wire [5:0] _T_37969; // @[Mux.scala 31:69:@16986.4]
  wire [5:0] _T_37970; // @[Mux.scala 31:69:@16987.4]
  wire [5:0] _T_37971; // @[Mux.scala 31:69:@16988.4]
  wire [5:0] _T_37972; // @[Mux.scala 31:69:@16989.4]
  wire [5:0] _T_37973; // @[Mux.scala 31:69:@16990.4]
  wire [5:0] _T_37974; // @[Mux.scala 31:69:@16991.4]
  wire [5:0] _T_37975; // @[Mux.scala 31:69:@16992.4]
  wire [5:0] _T_37976; // @[Mux.scala 31:69:@16993.4]
  wire [5:0] _T_37977; // @[Mux.scala 31:69:@16994.4]
  wire [5:0] _T_37978; // @[Mux.scala 31:69:@16995.4]
  wire [5:0] _T_37979; // @[Mux.scala 31:69:@16996.4]
  wire [5:0] _T_37980; // @[Mux.scala 31:69:@16997.4]
  wire [5:0] _T_37981; // @[Mux.scala 31:69:@16998.4]
  wire [5:0] _T_37982; // @[Mux.scala 31:69:@16999.4]
  wire [5:0] _T_37983; // @[Mux.scala 31:69:@17000.4]
  wire [5:0] _T_37984; // @[Mux.scala 31:69:@17001.4]
  wire [5:0] _T_37985; // @[Mux.scala 31:69:@17002.4]
  wire [5:0] _T_37986; // @[Mux.scala 31:69:@17003.4]
  wire [5:0] _T_37987; // @[Mux.scala 31:69:@17004.4]
  wire [5:0] _T_37988; // @[Mux.scala 31:69:@17005.4]
  wire [5:0] _T_37989; // @[Mux.scala 31:69:@17006.4]
  wire [5:0] _T_37990; // @[Mux.scala 31:69:@17007.4]
  wire [5:0] select_52; // @[Mux.scala 31:69:@17008.4]
  wire [47:0] _GEN_3329; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3330; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3331; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3332; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3333; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3334; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3335; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3336; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3337; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3338; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3339; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3340; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3341; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3342; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3343; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3344; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3345; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3346; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3347; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3348; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3349; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3350; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3351; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3352; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3353; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3354; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3355; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3356; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3357; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3358; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3359; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3360; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3361; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3362; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3363; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3364; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3365; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3366; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3367; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3368; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3369; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3370; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3371; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3372; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3373; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3374; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3375; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3376; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3377; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3378; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3379; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3380; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3381; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3382; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3383; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3384; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3385; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3386; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3387; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3388; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3389; // @[Switch.scala 33:19:@17010.4]
  wire [47:0] _GEN_3390; // @[Switch.scala 33:19:@17010.4]
  wire [7:0] _T_37999; // @[Switch.scala 34:32:@17017.4]
  wire [15:0] _T_38007; // @[Switch.scala 34:32:@17025.4]
  wire [7:0] _T_38014; // @[Switch.scala 34:32:@17032.4]
  wire [31:0] _T_38023; // @[Switch.scala 34:32:@17041.4]
  wire [7:0] _T_38030; // @[Switch.scala 34:32:@17048.4]
  wire [15:0] _T_38038; // @[Switch.scala 34:32:@17056.4]
  wire [7:0] _T_38045; // @[Switch.scala 34:32:@17063.4]
  wire [31:0] _T_38054; // @[Switch.scala 34:32:@17072.4]
  wire [63:0] _T_38055; // @[Switch.scala 34:32:@17073.4]
  wire  _T_38059; // @[Switch.scala 30:53:@17076.4]
  wire  valid_53_0; // @[Switch.scala 30:36:@17077.4]
  wire  _T_38062; // @[Switch.scala 30:53:@17079.4]
  wire  valid_53_1; // @[Switch.scala 30:36:@17080.4]
  wire  _T_38065; // @[Switch.scala 30:53:@17082.4]
  wire  valid_53_2; // @[Switch.scala 30:36:@17083.4]
  wire  _T_38068; // @[Switch.scala 30:53:@17085.4]
  wire  valid_53_3; // @[Switch.scala 30:36:@17086.4]
  wire  _T_38071; // @[Switch.scala 30:53:@17088.4]
  wire  valid_53_4; // @[Switch.scala 30:36:@17089.4]
  wire  _T_38074; // @[Switch.scala 30:53:@17091.4]
  wire  valid_53_5; // @[Switch.scala 30:36:@17092.4]
  wire  _T_38077; // @[Switch.scala 30:53:@17094.4]
  wire  valid_53_6; // @[Switch.scala 30:36:@17095.4]
  wire  _T_38080; // @[Switch.scala 30:53:@17097.4]
  wire  valid_53_7; // @[Switch.scala 30:36:@17098.4]
  wire  _T_38083; // @[Switch.scala 30:53:@17100.4]
  wire  valid_53_8; // @[Switch.scala 30:36:@17101.4]
  wire  _T_38086; // @[Switch.scala 30:53:@17103.4]
  wire  valid_53_9; // @[Switch.scala 30:36:@17104.4]
  wire  _T_38089; // @[Switch.scala 30:53:@17106.4]
  wire  valid_53_10; // @[Switch.scala 30:36:@17107.4]
  wire  _T_38092; // @[Switch.scala 30:53:@17109.4]
  wire  valid_53_11; // @[Switch.scala 30:36:@17110.4]
  wire  _T_38095; // @[Switch.scala 30:53:@17112.4]
  wire  valid_53_12; // @[Switch.scala 30:36:@17113.4]
  wire  _T_38098; // @[Switch.scala 30:53:@17115.4]
  wire  valid_53_13; // @[Switch.scala 30:36:@17116.4]
  wire  _T_38101; // @[Switch.scala 30:53:@17118.4]
  wire  valid_53_14; // @[Switch.scala 30:36:@17119.4]
  wire  _T_38104; // @[Switch.scala 30:53:@17121.4]
  wire  valid_53_15; // @[Switch.scala 30:36:@17122.4]
  wire  _T_38107; // @[Switch.scala 30:53:@17124.4]
  wire  valid_53_16; // @[Switch.scala 30:36:@17125.4]
  wire  _T_38110; // @[Switch.scala 30:53:@17127.4]
  wire  valid_53_17; // @[Switch.scala 30:36:@17128.4]
  wire  _T_38113; // @[Switch.scala 30:53:@17130.4]
  wire  valid_53_18; // @[Switch.scala 30:36:@17131.4]
  wire  _T_38116; // @[Switch.scala 30:53:@17133.4]
  wire  valid_53_19; // @[Switch.scala 30:36:@17134.4]
  wire  _T_38119; // @[Switch.scala 30:53:@17136.4]
  wire  valid_53_20; // @[Switch.scala 30:36:@17137.4]
  wire  _T_38122; // @[Switch.scala 30:53:@17139.4]
  wire  valid_53_21; // @[Switch.scala 30:36:@17140.4]
  wire  _T_38125; // @[Switch.scala 30:53:@17142.4]
  wire  valid_53_22; // @[Switch.scala 30:36:@17143.4]
  wire  _T_38128; // @[Switch.scala 30:53:@17145.4]
  wire  valid_53_23; // @[Switch.scala 30:36:@17146.4]
  wire  _T_38131; // @[Switch.scala 30:53:@17148.4]
  wire  valid_53_24; // @[Switch.scala 30:36:@17149.4]
  wire  _T_38134; // @[Switch.scala 30:53:@17151.4]
  wire  valid_53_25; // @[Switch.scala 30:36:@17152.4]
  wire  _T_38137; // @[Switch.scala 30:53:@17154.4]
  wire  valid_53_26; // @[Switch.scala 30:36:@17155.4]
  wire  _T_38140; // @[Switch.scala 30:53:@17157.4]
  wire  valid_53_27; // @[Switch.scala 30:36:@17158.4]
  wire  _T_38143; // @[Switch.scala 30:53:@17160.4]
  wire  valid_53_28; // @[Switch.scala 30:36:@17161.4]
  wire  _T_38146; // @[Switch.scala 30:53:@17163.4]
  wire  valid_53_29; // @[Switch.scala 30:36:@17164.4]
  wire  _T_38149; // @[Switch.scala 30:53:@17166.4]
  wire  valid_53_30; // @[Switch.scala 30:36:@17167.4]
  wire  _T_38152; // @[Switch.scala 30:53:@17169.4]
  wire  valid_53_31; // @[Switch.scala 30:36:@17170.4]
  wire  _T_38155; // @[Switch.scala 30:53:@17172.4]
  wire  valid_53_32; // @[Switch.scala 30:36:@17173.4]
  wire  _T_38158; // @[Switch.scala 30:53:@17175.4]
  wire  valid_53_33; // @[Switch.scala 30:36:@17176.4]
  wire  _T_38161; // @[Switch.scala 30:53:@17178.4]
  wire  valid_53_34; // @[Switch.scala 30:36:@17179.4]
  wire  _T_38164; // @[Switch.scala 30:53:@17181.4]
  wire  valid_53_35; // @[Switch.scala 30:36:@17182.4]
  wire  _T_38167; // @[Switch.scala 30:53:@17184.4]
  wire  valid_53_36; // @[Switch.scala 30:36:@17185.4]
  wire  _T_38170; // @[Switch.scala 30:53:@17187.4]
  wire  valid_53_37; // @[Switch.scala 30:36:@17188.4]
  wire  _T_38173; // @[Switch.scala 30:53:@17190.4]
  wire  valid_53_38; // @[Switch.scala 30:36:@17191.4]
  wire  _T_38176; // @[Switch.scala 30:53:@17193.4]
  wire  valid_53_39; // @[Switch.scala 30:36:@17194.4]
  wire  _T_38179; // @[Switch.scala 30:53:@17196.4]
  wire  valid_53_40; // @[Switch.scala 30:36:@17197.4]
  wire  _T_38182; // @[Switch.scala 30:53:@17199.4]
  wire  valid_53_41; // @[Switch.scala 30:36:@17200.4]
  wire  _T_38185; // @[Switch.scala 30:53:@17202.4]
  wire  valid_53_42; // @[Switch.scala 30:36:@17203.4]
  wire  _T_38188; // @[Switch.scala 30:53:@17205.4]
  wire  valid_53_43; // @[Switch.scala 30:36:@17206.4]
  wire  _T_38191; // @[Switch.scala 30:53:@17208.4]
  wire  valid_53_44; // @[Switch.scala 30:36:@17209.4]
  wire  _T_38194; // @[Switch.scala 30:53:@17211.4]
  wire  valid_53_45; // @[Switch.scala 30:36:@17212.4]
  wire  _T_38197; // @[Switch.scala 30:53:@17214.4]
  wire  valid_53_46; // @[Switch.scala 30:36:@17215.4]
  wire  _T_38200; // @[Switch.scala 30:53:@17217.4]
  wire  valid_53_47; // @[Switch.scala 30:36:@17218.4]
  wire  _T_38203; // @[Switch.scala 30:53:@17220.4]
  wire  valid_53_48; // @[Switch.scala 30:36:@17221.4]
  wire  _T_38206; // @[Switch.scala 30:53:@17223.4]
  wire  valid_53_49; // @[Switch.scala 30:36:@17224.4]
  wire  _T_38209; // @[Switch.scala 30:53:@17226.4]
  wire  valid_53_50; // @[Switch.scala 30:36:@17227.4]
  wire  _T_38212; // @[Switch.scala 30:53:@17229.4]
  wire  valid_53_51; // @[Switch.scala 30:36:@17230.4]
  wire  _T_38215; // @[Switch.scala 30:53:@17232.4]
  wire  valid_53_52; // @[Switch.scala 30:36:@17233.4]
  wire  _T_38218; // @[Switch.scala 30:53:@17235.4]
  wire  valid_53_53; // @[Switch.scala 30:36:@17236.4]
  wire  _T_38221; // @[Switch.scala 30:53:@17238.4]
  wire  valid_53_54; // @[Switch.scala 30:36:@17239.4]
  wire  _T_38224; // @[Switch.scala 30:53:@17241.4]
  wire  valid_53_55; // @[Switch.scala 30:36:@17242.4]
  wire  _T_38227; // @[Switch.scala 30:53:@17244.4]
  wire  valid_53_56; // @[Switch.scala 30:36:@17245.4]
  wire  _T_38230; // @[Switch.scala 30:53:@17247.4]
  wire  valid_53_57; // @[Switch.scala 30:36:@17248.4]
  wire  _T_38233; // @[Switch.scala 30:53:@17250.4]
  wire  valid_53_58; // @[Switch.scala 30:36:@17251.4]
  wire  _T_38236; // @[Switch.scala 30:53:@17253.4]
  wire  valid_53_59; // @[Switch.scala 30:36:@17254.4]
  wire  _T_38239; // @[Switch.scala 30:53:@17256.4]
  wire  valid_53_60; // @[Switch.scala 30:36:@17257.4]
  wire  _T_38242; // @[Switch.scala 30:53:@17259.4]
  wire  valid_53_61; // @[Switch.scala 30:36:@17260.4]
  wire  _T_38245; // @[Switch.scala 30:53:@17262.4]
  wire  valid_53_62; // @[Switch.scala 30:36:@17263.4]
  wire  _T_38248; // @[Switch.scala 30:53:@17265.4]
  wire  valid_53_63; // @[Switch.scala 30:36:@17266.4]
  wire [5:0] _T_38314; // @[Mux.scala 31:69:@17268.4]
  wire [5:0] _T_38315; // @[Mux.scala 31:69:@17269.4]
  wire [5:0] _T_38316; // @[Mux.scala 31:69:@17270.4]
  wire [5:0] _T_38317; // @[Mux.scala 31:69:@17271.4]
  wire [5:0] _T_38318; // @[Mux.scala 31:69:@17272.4]
  wire [5:0] _T_38319; // @[Mux.scala 31:69:@17273.4]
  wire [5:0] _T_38320; // @[Mux.scala 31:69:@17274.4]
  wire [5:0] _T_38321; // @[Mux.scala 31:69:@17275.4]
  wire [5:0] _T_38322; // @[Mux.scala 31:69:@17276.4]
  wire [5:0] _T_38323; // @[Mux.scala 31:69:@17277.4]
  wire [5:0] _T_38324; // @[Mux.scala 31:69:@17278.4]
  wire [5:0] _T_38325; // @[Mux.scala 31:69:@17279.4]
  wire [5:0] _T_38326; // @[Mux.scala 31:69:@17280.4]
  wire [5:0] _T_38327; // @[Mux.scala 31:69:@17281.4]
  wire [5:0] _T_38328; // @[Mux.scala 31:69:@17282.4]
  wire [5:0] _T_38329; // @[Mux.scala 31:69:@17283.4]
  wire [5:0] _T_38330; // @[Mux.scala 31:69:@17284.4]
  wire [5:0] _T_38331; // @[Mux.scala 31:69:@17285.4]
  wire [5:0] _T_38332; // @[Mux.scala 31:69:@17286.4]
  wire [5:0] _T_38333; // @[Mux.scala 31:69:@17287.4]
  wire [5:0] _T_38334; // @[Mux.scala 31:69:@17288.4]
  wire [5:0] _T_38335; // @[Mux.scala 31:69:@17289.4]
  wire [5:0] _T_38336; // @[Mux.scala 31:69:@17290.4]
  wire [5:0] _T_38337; // @[Mux.scala 31:69:@17291.4]
  wire [5:0] _T_38338; // @[Mux.scala 31:69:@17292.4]
  wire [5:0] _T_38339; // @[Mux.scala 31:69:@17293.4]
  wire [5:0] _T_38340; // @[Mux.scala 31:69:@17294.4]
  wire [5:0] _T_38341; // @[Mux.scala 31:69:@17295.4]
  wire [5:0] _T_38342; // @[Mux.scala 31:69:@17296.4]
  wire [5:0] _T_38343; // @[Mux.scala 31:69:@17297.4]
  wire [5:0] _T_38344; // @[Mux.scala 31:69:@17298.4]
  wire [5:0] _T_38345; // @[Mux.scala 31:69:@17299.4]
  wire [5:0] _T_38346; // @[Mux.scala 31:69:@17300.4]
  wire [5:0] _T_38347; // @[Mux.scala 31:69:@17301.4]
  wire [5:0] _T_38348; // @[Mux.scala 31:69:@17302.4]
  wire [5:0] _T_38349; // @[Mux.scala 31:69:@17303.4]
  wire [5:0] _T_38350; // @[Mux.scala 31:69:@17304.4]
  wire [5:0] _T_38351; // @[Mux.scala 31:69:@17305.4]
  wire [5:0] _T_38352; // @[Mux.scala 31:69:@17306.4]
  wire [5:0] _T_38353; // @[Mux.scala 31:69:@17307.4]
  wire [5:0] _T_38354; // @[Mux.scala 31:69:@17308.4]
  wire [5:0] _T_38355; // @[Mux.scala 31:69:@17309.4]
  wire [5:0] _T_38356; // @[Mux.scala 31:69:@17310.4]
  wire [5:0] _T_38357; // @[Mux.scala 31:69:@17311.4]
  wire [5:0] _T_38358; // @[Mux.scala 31:69:@17312.4]
  wire [5:0] _T_38359; // @[Mux.scala 31:69:@17313.4]
  wire [5:0] _T_38360; // @[Mux.scala 31:69:@17314.4]
  wire [5:0] _T_38361; // @[Mux.scala 31:69:@17315.4]
  wire [5:0] _T_38362; // @[Mux.scala 31:69:@17316.4]
  wire [5:0] _T_38363; // @[Mux.scala 31:69:@17317.4]
  wire [5:0] _T_38364; // @[Mux.scala 31:69:@17318.4]
  wire [5:0] _T_38365; // @[Mux.scala 31:69:@17319.4]
  wire [5:0] _T_38366; // @[Mux.scala 31:69:@17320.4]
  wire [5:0] _T_38367; // @[Mux.scala 31:69:@17321.4]
  wire [5:0] _T_38368; // @[Mux.scala 31:69:@17322.4]
  wire [5:0] _T_38369; // @[Mux.scala 31:69:@17323.4]
  wire [5:0] _T_38370; // @[Mux.scala 31:69:@17324.4]
  wire [5:0] _T_38371; // @[Mux.scala 31:69:@17325.4]
  wire [5:0] _T_38372; // @[Mux.scala 31:69:@17326.4]
  wire [5:0] _T_38373; // @[Mux.scala 31:69:@17327.4]
  wire [5:0] _T_38374; // @[Mux.scala 31:69:@17328.4]
  wire [5:0] _T_38375; // @[Mux.scala 31:69:@17329.4]
  wire [5:0] select_53; // @[Mux.scala 31:69:@17330.4]
  wire [47:0] _GEN_3393; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3394; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3395; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3396; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3397; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3398; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3399; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3400; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3401; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3402; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3403; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3404; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3405; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3406; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3407; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3408; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3409; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3410; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3411; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3412; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3413; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3414; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3415; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3416; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3417; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3418; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3419; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3420; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3421; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3422; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3423; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3424; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3425; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3426; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3427; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3428; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3429; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3430; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3431; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3432; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3433; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3434; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3435; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3436; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3437; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3438; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3439; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3440; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3441; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3442; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3443; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3444; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3445; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3446; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3447; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3448; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3449; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3450; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3451; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3452; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3453; // @[Switch.scala 33:19:@17332.4]
  wire [47:0] _GEN_3454; // @[Switch.scala 33:19:@17332.4]
  wire [7:0] _T_38384; // @[Switch.scala 34:32:@17339.4]
  wire [15:0] _T_38392; // @[Switch.scala 34:32:@17347.4]
  wire [7:0] _T_38399; // @[Switch.scala 34:32:@17354.4]
  wire [31:0] _T_38408; // @[Switch.scala 34:32:@17363.4]
  wire [7:0] _T_38415; // @[Switch.scala 34:32:@17370.4]
  wire [15:0] _T_38423; // @[Switch.scala 34:32:@17378.4]
  wire [7:0] _T_38430; // @[Switch.scala 34:32:@17385.4]
  wire [31:0] _T_38439; // @[Switch.scala 34:32:@17394.4]
  wire [63:0] _T_38440; // @[Switch.scala 34:32:@17395.4]
  wire  _T_38444; // @[Switch.scala 30:53:@17398.4]
  wire  valid_54_0; // @[Switch.scala 30:36:@17399.4]
  wire  _T_38447; // @[Switch.scala 30:53:@17401.4]
  wire  valid_54_1; // @[Switch.scala 30:36:@17402.4]
  wire  _T_38450; // @[Switch.scala 30:53:@17404.4]
  wire  valid_54_2; // @[Switch.scala 30:36:@17405.4]
  wire  _T_38453; // @[Switch.scala 30:53:@17407.4]
  wire  valid_54_3; // @[Switch.scala 30:36:@17408.4]
  wire  _T_38456; // @[Switch.scala 30:53:@17410.4]
  wire  valid_54_4; // @[Switch.scala 30:36:@17411.4]
  wire  _T_38459; // @[Switch.scala 30:53:@17413.4]
  wire  valid_54_5; // @[Switch.scala 30:36:@17414.4]
  wire  _T_38462; // @[Switch.scala 30:53:@17416.4]
  wire  valid_54_6; // @[Switch.scala 30:36:@17417.4]
  wire  _T_38465; // @[Switch.scala 30:53:@17419.4]
  wire  valid_54_7; // @[Switch.scala 30:36:@17420.4]
  wire  _T_38468; // @[Switch.scala 30:53:@17422.4]
  wire  valid_54_8; // @[Switch.scala 30:36:@17423.4]
  wire  _T_38471; // @[Switch.scala 30:53:@17425.4]
  wire  valid_54_9; // @[Switch.scala 30:36:@17426.4]
  wire  _T_38474; // @[Switch.scala 30:53:@17428.4]
  wire  valid_54_10; // @[Switch.scala 30:36:@17429.4]
  wire  _T_38477; // @[Switch.scala 30:53:@17431.4]
  wire  valid_54_11; // @[Switch.scala 30:36:@17432.4]
  wire  _T_38480; // @[Switch.scala 30:53:@17434.4]
  wire  valid_54_12; // @[Switch.scala 30:36:@17435.4]
  wire  _T_38483; // @[Switch.scala 30:53:@17437.4]
  wire  valid_54_13; // @[Switch.scala 30:36:@17438.4]
  wire  _T_38486; // @[Switch.scala 30:53:@17440.4]
  wire  valid_54_14; // @[Switch.scala 30:36:@17441.4]
  wire  _T_38489; // @[Switch.scala 30:53:@17443.4]
  wire  valid_54_15; // @[Switch.scala 30:36:@17444.4]
  wire  _T_38492; // @[Switch.scala 30:53:@17446.4]
  wire  valid_54_16; // @[Switch.scala 30:36:@17447.4]
  wire  _T_38495; // @[Switch.scala 30:53:@17449.4]
  wire  valid_54_17; // @[Switch.scala 30:36:@17450.4]
  wire  _T_38498; // @[Switch.scala 30:53:@17452.4]
  wire  valid_54_18; // @[Switch.scala 30:36:@17453.4]
  wire  _T_38501; // @[Switch.scala 30:53:@17455.4]
  wire  valid_54_19; // @[Switch.scala 30:36:@17456.4]
  wire  _T_38504; // @[Switch.scala 30:53:@17458.4]
  wire  valid_54_20; // @[Switch.scala 30:36:@17459.4]
  wire  _T_38507; // @[Switch.scala 30:53:@17461.4]
  wire  valid_54_21; // @[Switch.scala 30:36:@17462.4]
  wire  _T_38510; // @[Switch.scala 30:53:@17464.4]
  wire  valid_54_22; // @[Switch.scala 30:36:@17465.4]
  wire  _T_38513; // @[Switch.scala 30:53:@17467.4]
  wire  valid_54_23; // @[Switch.scala 30:36:@17468.4]
  wire  _T_38516; // @[Switch.scala 30:53:@17470.4]
  wire  valid_54_24; // @[Switch.scala 30:36:@17471.4]
  wire  _T_38519; // @[Switch.scala 30:53:@17473.4]
  wire  valid_54_25; // @[Switch.scala 30:36:@17474.4]
  wire  _T_38522; // @[Switch.scala 30:53:@17476.4]
  wire  valid_54_26; // @[Switch.scala 30:36:@17477.4]
  wire  _T_38525; // @[Switch.scala 30:53:@17479.4]
  wire  valid_54_27; // @[Switch.scala 30:36:@17480.4]
  wire  _T_38528; // @[Switch.scala 30:53:@17482.4]
  wire  valid_54_28; // @[Switch.scala 30:36:@17483.4]
  wire  _T_38531; // @[Switch.scala 30:53:@17485.4]
  wire  valid_54_29; // @[Switch.scala 30:36:@17486.4]
  wire  _T_38534; // @[Switch.scala 30:53:@17488.4]
  wire  valid_54_30; // @[Switch.scala 30:36:@17489.4]
  wire  _T_38537; // @[Switch.scala 30:53:@17491.4]
  wire  valid_54_31; // @[Switch.scala 30:36:@17492.4]
  wire  _T_38540; // @[Switch.scala 30:53:@17494.4]
  wire  valid_54_32; // @[Switch.scala 30:36:@17495.4]
  wire  _T_38543; // @[Switch.scala 30:53:@17497.4]
  wire  valid_54_33; // @[Switch.scala 30:36:@17498.4]
  wire  _T_38546; // @[Switch.scala 30:53:@17500.4]
  wire  valid_54_34; // @[Switch.scala 30:36:@17501.4]
  wire  _T_38549; // @[Switch.scala 30:53:@17503.4]
  wire  valid_54_35; // @[Switch.scala 30:36:@17504.4]
  wire  _T_38552; // @[Switch.scala 30:53:@17506.4]
  wire  valid_54_36; // @[Switch.scala 30:36:@17507.4]
  wire  _T_38555; // @[Switch.scala 30:53:@17509.4]
  wire  valid_54_37; // @[Switch.scala 30:36:@17510.4]
  wire  _T_38558; // @[Switch.scala 30:53:@17512.4]
  wire  valid_54_38; // @[Switch.scala 30:36:@17513.4]
  wire  _T_38561; // @[Switch.scala 30:53:@17515.4]
  wire  valid_54_39; // @[Switch.scala 30:36:@17516.4]
  wire  _T_38564; // @[Switch.scala 30:53:@17518.4]
  wire  valid_54_40; // @[Switch.scala 30:36:@17519.4]
  wire  _T_38567; // @[Switch.scala 30:53:@17521.4]
  wire  valid_54_41; // @[Switch.scala 30:36:@17522.4]
  wire  _T_38570; // @[Switch.scala 30:53:@17524.4]
  wire  valid_54_42; // @[Switch.scala 30:36:@17525.4]
  wire  _T_38573; // @[Switch.scala 30:53:@17527.4]
  wire  valid_54_43; // @[Switch.scala 30:36:@17528.4]
  wire  _T_38576; // @[Switch.scala 30:53:@17530.4]
  wire  valid_54_44; // @[Switch.scala 30:36:@17531.4]
  wire  _T_38579; // @[Switch.scala 30:53:@17533.4]
  wire  valid_54_45; // @[Switch.scala 30:36:@17534.4]
  wire  _T_38582; // @[Switch.scala 30:53:@17536.4]
  wire  valid_54_46; // @[Switch.scala 30:36:@17537.4]
  wire  _T_38585; // @[Switch.scala 30:53:@17539.4]
  wire  valid_54_47; // @[Switch.scala 30:36:@17540.4]
  wire  _T_38588; // @[Switch.scala 30:53:@17542.4]
  wire  valid_54_48; // @[Switch.scala 30:36:@17543.4]
  wire  _T_38591; // @[Switch.scala 30:53:@17545.4]
  wire  valid_54_49; // @[Switch.scala 30:36:@17546.4]
  wire  _T_38594; // @[Switch.scala 30:53:@17548.4]
  wire  valid_54_50; // @[Switch.scala 30:36:@17549.4]
  wire  _T_38597; // @[Switch.scala 30:53:@17551.4]
  wire  valid_54_51; // @[Switch.scala 30:36:@17552.4]
  wire  _T_38600; // @[Switch.scala 30:53:@17554.4]
  wire  valid_54_52; // @[Switch.scala 30:36:@17555.4]
  wire  _T_38603; // @[Switch.scala 30:53:@17557.4]
  wire  valid_54_53; // @[Switch.scala 30:36:@17558.4]
  wire  _T_38606; // @[Switch.scala 30:53:@17560.4]
  wire  valid_54_54; // @[Switch.scala 30:36:@17561.4]
  wire  _T_38609; // @[Switch.scala 30:53:@17563.4]
  wire  valid_54_55; // @[Switch.scala 30:36:@17564.4]
  wire  _T_38612; // @[Switch.scala 30:53:@17566.4]
  wire  valid_54_56; // @[Switch.scala 30:36:@17567.4]
  wire  _T_38615; // @[Switch.scala 30:53:@17569.4]
  wire  valid_54_57; // @[Switch.scala 30:36:@17570.4]
  wire  _T_38618; // @[Switch.scala 30:53:@17572.4]
  wire  valid_54_58; // @[Switch.scala 30:36:@17573.4]
  wire  _T_38621; // @[Switch.scala 30:53:@17575.4]
  wire  valid_54_59; // @[Switch.scala 30:36:@17576.4]
  wire  _T_38624; // @[Switch.scala 30:53:@17578.4]
  wire  valid_54_60; // @[Switch.scala 30:36:@17579.4]
  wire  _T_38627; // @[Switch.scala 30:53:@17581.4]
  wire  valid_54_61; // @[Switch.scala 30:36:@17582.4]
  wire  _T_38630; // @[Switch.scala 30:53:@17584.4]
  wire  valid_54_62; // @[Switch.scala 30:36:@17585.4]
  wire  _T_38633; // @[Switch.scala 30:53:@17587.4]
  wire  valid_54_63; // @[Switch.scala 30:36:@17588.4]
  wire [5:0] _T_38699; // @[Mux.scala 31:69:@17590.4]
  wire [5:0] _T_38700; // @[Mux.scala 31:69:@17591.4]
  wire [5:0] _T_38701; // @[Mux.scala 31:69:@17592.4]
  wire [5:0] _T_38702; // @[Mux.scala 31:69:@17593.4]
  wire [5:0] _T_38703; // @[Mux.scala 31:69:@17594.4]
  wire [5:0] _T_38704; // @[Mux.scala 31:69:@17595.4]
  wire [5:0] _T_38705; // @[Mux.scala 31:69:@17596.4]
  wire [5:0] _T_38706; // @[Mux.scala 31:69:@17597.4]
  wire [5:0] _T_38707; // @[Mux.scala 31:69:@17598.4]
  wire [5:0] _T_38708; // @[Mux.scala 31:69:@17599.4]
  wire [5:0] _T_38709; // @[Mux.scala 31:69:@17600.4]
  wire [5:0] _T_38710; // @[Mux.scala 31:69:@17601.4]
  wire [5:0] _T_38711; // @[Mux.scala 31:69:@17602.4]
  wire [5:0] _T_38712; // @[Mux.scala 31:69:@17603.4]
  wire [5:0] _T_38713; // @[Mux.scala 31:69:@17604.4]
  wire [5:0] _T_38714; // @[Mux.scala 31:69:@17605.4]
  wire [5:0] _T_38715; // @[Mux.scala 31:69:@17606.4]
  wire [5:0] _T_38716; // @[Mux.scala 31:69:@17607.4]
  wire [5:0] _T_38717; // @[Mux.scala 31:69:@17608.4]
  wire [5:0] _T_38718; // @[Mux.scala 31:69:@17609.4]
  wire [5:0] _T_38719; // @[Mux.scala 31:69:@17610.4]
  wire [5:0] _T_38720; // @[Mux.scala 31:69:@17611.4]
  wire [5:0] _T_38721; // @[Mux.scala 31:69:@17612.4]
  wire [5:0] _T_38722; // @[Mux.scala 31:69:@17613.4]
  wire [5:0] _T_38723; // @[Mux.scala 31:69:@17614.4]
  wire [5:0] _T_38724; // @[Mux.scala 31:69:@17615.4]
  wire [5:0] _T_38725; // @[Mux.scala 31:69:@17616.4]
  wire [5:0] _T_38726; // @[Mux.scala 31:69:@17617.4]
  wire [5:0] _T_38727; // @[Mux.scala 31:69:@17618.4]
  wire [5:0] _T_38728; // @[Mux.scala 31:69:@17619.4]
  wire [5:0] _T_38729; // @[Mux.scala 31:69:@17620.4]
  wire [5:0] _T_38730; // @[Mux.scala 31:69:@17621.4]
  wire [5:0] _T_38731; // @[Mux.scala 31:69:@17622.4]
  wire [5:0] _T_38732; // @[Mux.scala 31:69:@17623.4]
  wire [5:0] _T_38733; // @[Mux.scala 31:69:@17624.4]
  wire [5:0] _T_38734; // @[Mux.scala 31:69:@17625.4]
  wire [5:0] _T_38735; // @[Mux.scala 31:69:@17626.4]
  wire [5:0] _T_38736; // @[Mux.scala 31:69:@17627.4]
  wire [5:0] _T_38737; // @[Mux.scala 31:69:@17628.4]
  wire [5:0] _T_38738; // @[Mux.scala 31:69:@17629.4]
  wire [5:0] _T_38739; // @[Mux.scala 31:69:@17630.4]
  wire [5:0] _T_38740; // @[Mux.scala 31:69:@17631.4]
  wire [5:0] _T_38741; // @[Mux.scala 31:69:@17632.4]
  wire [5:0] _T_38742; // @[Mux.scala 31:69:@17633.4]
  wire [5:0] _T_38743; // @[Mux.scala 31:69:@17634.4]
  wire [5:0] _T_38744; // @[Mux.scala 31:69:@17635.4]
  wire [5:0] _T_38745; // @[Mux.scala 31:69:@17636.4]
  wire [5:0] _T_38746; // @[Mux.scala 31:69:@17637.4]
  wire [5:0] _T_38747; // @[Mux.scala 31:69:@17638.4]
  wire [5:0] _T_38748; // @[Mux.scala 31:69:@17639.4]
  wire [5:0] _T_38749; // @[Mux.scala 31:69:@17640.4]
  wire [5:0] _T_38750; // @[Mux.scala 31:69:@17641.4]
  wire [5:0] _T_38751; // @[Mux.scala 31:69:@17642.4]
  wire [5:0] _T_38752; // @[Mux.scala 31:69:@17643.4]
  wire [5:0] _T_38753; // @[Mux.scala 31:69:@17644.4]
  wire [5:0] _T_38754; // @[Mux.scala 31:69:@17645.4]
  wire [5:0] _T_38755; // @[Mux.scala 31:69:@17646.4]
  wire [5:0] _T_38756; // @[Mux.scala 31:69:@17647.4]
  wire [5:0] _T_38757; // @[Mux.scala 31:69:@17648.4]
  wire [5:0] _T_38758; // @[Mux.scala 31:69:@17649.4]
  wire [5:0] _T_38759; // @[Mux.scala 31:69:@17650.4]
  wire [5:0] _T_38760; // @[Mux.scala 31:69:@17651.4]
  wire [5:0] select_54; // @[Mux.scala 31:69:@17652.4]
  wire [47:0] _GEN_3457; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3458; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3459; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3460; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3461; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3462; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3463; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3464; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3465; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3466; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3467; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3468; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3469; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3470; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3471; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3472; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3473; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3474; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3475; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3476; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3477; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3478; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3479; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3480; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3481; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3482; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3483; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3484; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3485; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3486; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3487; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3488; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3489; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3490; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3491; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3492; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3493; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3494; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3495; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3496; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3497; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3498; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3499; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3500; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3501; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3502; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3503; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3504; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3505; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3506; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3507; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3508; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3509; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3510; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3511; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3512; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3513; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3514; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3515; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3516; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3517; // @[Switch.scala 33:19:@17654.4]
  wire [47:0] _GEN_3518; // @[Switch.scala 33:19:@17654.4]
  wire [7:0] _T_38769; // @[Switch.scala 34:32:@17661.4]
  wire [15:0] _T_38777; // @[Switch.scala 34:32:@17669.4]
  wire [7:0] _T_38784; // @[Switch.scala 34:32:@17676.4]
  wire [31:0] _T_38793; // @[Switch.scala 34:32:@17685.4]
  wire [7:0] _T_38800; // @[Switch.scala 34:32:@17692.4]
  wire [15:0] _T_38808; // @[Switch.scala 34:32:@17700.4]
  wire [7:0] _T_38815; // @[Switch.scala 34:32:@17707.4]
  wire [31:0] _T_38824; // @[Switch.scala 34:32:@17716.4]
  wire [63:0] _T_38825; // @[Switch.scala 34:32:@17717.4]
  wire  _T_38829; // @[Switch.scala 30:53:@17720.4]
  wire  valid_55_0; // @[Switch.scala 30:36:@17721.4]
  wire  _T_38832; // @[Switch.scala 30:53:@17723.4]
  wire  valid_55_1; // @[Switch.scala 30:36:@17724.4]
  wire  _T_38835; // @[Switch.scala 30:53:@17726.4]
  wire  valid_55_2; // @[Switch.scala 30:36:@17727.4]
  wire  _T_38838; // @[Switch.scala 30:53:@17729.4]
  wire  valid_55_3; // @[Switch.scala 30:36:@17730.4]
  wire  _T_38841; // @[Switch.scala 30:53:@17732.4]
  wire  valid_55_4; // @[Switch.scala 30:36:@17733.4]
  wire  _T_38844; // @[Switch.scala 30:53:@17735.4]
  wire  valid_55_5; // @[Switch.scala 30:36:@17736.4]
  wire  _T_38847; // @[Switch.scala 30:53:@17738.4]
  wire  valid_55_6; // @[Switch.scala 30:36:@17739.4]
  wire  _T_38850; // @[Switch.scala 30:53:@17741.4]
  wire  valid_55_7; // @[Switch.scala 30:36:@17742.4]
  wire  _T_38853; // @[Switch.scala 30:53:@17744.4]
  wire  valid_55_8; // @[Switch.scala 30:36:@17745.4]
  wire  _T_38856; // @[Switch.scala 30:53:@17747.4]
  wire  valid_55_9; // @[Switch.scala 30:36:@17748.4]
  wire  _T_38859; // @[Switch.scala 30:53:@17750.4]
  wire  valid_55_10; // @[Switch.scala 30:36:@17751.4]
  wire  _T_38862; // @[Switch.scala 30:53:@17753.4]
  wire  valid_55_11; // @[Switch.scala 30:36:@17754.4]
  wire  _T_38865; // @[Switch.scala 30:53:@17756.4]
  wire  valid_55_12; // @[Switch.scala 30:36:@17757.4]
  wire  _T_38868; // @[Switch.scala 30:53:@17759.4]
  wire  valid_55_13; // @[Switch.scala 30:36:@17760.4]
  wire  _T_38871; // @[Switch.scala 30:53:@17762.4]
  wire  valid_55_14; // @[Switch.scala 30:36:@17763.4]
  wire  _T_38874; // @[Switch.scala 30:53:@17765.4]
  wire  valid_55_15; // @[Switch.scala 30:36:@17766.4]
  wire  _T_38877; // @[Switch.scala 30:53:@17768.4]
  wire  valid_55_16; // @[Switch.scala 30:36:@17769.4]
  wire  _T_38880; // @[Switch.scala 30:53:@17771.4]
  wire  valid_55_17; // @[Switch.scala 30:36:@17772.4]
  wire  _T_38883; // @[Switch.scala 30:53:@17774.4]
  wire  valid_55_18; // @[Switch.scala 30:36:@17775.4]
  wire  _T_38886; // @[Switch.scala 30:53:@17777.4]
  wire  valid_55_19; // @[Switch.scala 30:36:@17778.4]
  wire  _T_38889; // @[Switch.scala 30:53:@17780.4]
  wire  valid_55_20; // @[Switch.scala 30:36:@17781.4]
  wire  _T_38892; // @[Switch.scala 30:53:@17783.4]
  wire  valid_55_21; // @[Switch.scala 30:36:@17784.4]
  wire  _T_38895; // @[Switch.scala 30:53:@17786.4]
  wire  valid_55_22; // @[Switch.scala 30:36:@17787.4]
  wire  _T_38898; // @[Switch.scala 30:53:@17789.4]
  wire  valid_55_23; // @[Switch.scala 30:36:@17790.4]
  wire  _T_38901; // @[Switch.scala 30:53:@17792.4]
  wire  valid_55_24; // @[Switch.scala 30:36:@17793.4]
  wire  _T_38904; // @[Switch.scala 30:53:@17795.4]
  wire  valid_55_25; // @[Switch.scala 30:36:@17796.4]
  wire  _T_38907; // @[Switch.scala 30:53:@17798.4]
  wire  valid_55_26; // @[Switch.scala 30:36:@17799.4]
  wire  _T_38910; // @[Switch.scala 30:53:@17801.4]
  wire  valid_55_27; // @[Switch.scala 30:36:@17802.4]
  wire  _T_38913; // @[Switch.scala 30:53:@17804.4]
  wire  valid_55_28; // @[Switch.scala 30:36:@17805.4]
  wire  _T_38916; // @[Switch.scala 30:53:@17807.4]
  wire  valid_55_29; // @[Switch.scala 30:36:@17808.4]
  wire  _T_38919; // @[Switch.scala 30:53:@17810.4]
  wire  valid_55_30; // @[Switch.scala 30:36:@17811.4]
  wire  _T_38922; // @[Switch.scala 30:53:@17813.4]
  wire  valid_55_31; // @[Switch.scala 30:36:@17814.4]
  wire  _T_38925; // @[Switch.scala 30:53:@17816.4]
  wire  valid_55_32; // @[Switch.scala 30:36:@17817.4]
  wire  _T_38928; // @[Switch.scala 30:53:@17819.4]
  wire  valid_55_33; // @[Switch.scala 30:36:@17820.4]
  wire  _T_38931; // @[Switch.scala 30:53:@17822.4]
  wire  valid_55_34; // @[Switch.scala 30:36:@17823.4]
  wire  _T_38934; // @[Switch.scala 30:53:@17825.4]
  wire  valid_55_35; // @[Switch.scala 30:36:@17826.4]
  wire  _T_38937; // @[Switch.scala 30:53:@17828.4]
  wire  valid_55_36; // @[Switch.scala 30:36:@17829.4]
  wire  _T_38940; // @[Switch.scala 30:53:@17831.4]
  wire  valid_55_37; // @[Switch.scala 30:36:@17832.4]
  wire  _T_38943; // @[Switch.scala 30:53:@17834.4]
  wire  valid_55_38; // @[Switch.scala 30:36:@17835.4]
  wire  _T_38946; // @[Switch.scala 30:53:@17837.4]
  wire  valid_55_39; // @[Switch.scala 30:36:@17838.4]
  wire  _T_38949; // @[Switch.scala 30:53:@17840.4]
  wire  valid_55_40; // @[Switch.scala 30:36:@17841.4]
  wire  _T_38952; // @[Switch.scala 30:53:@17843.4]
  wire  valid_55_41; // @[Switch.scala 30:36:@17844.4]
  wire  _T_38955; // @[Switch.scala 30:53:@17846.4]
  wire  valid_55_42; // @[Switch.scala 30:36:@17847.4]
  wire  _T_38958; // @[Switch.scala 30:53:@17849.4]
  wire  valid_55_43; // @[Switch.scala 30:36:@17850.4]
  wire  _T_38961; // @[Switch.scala 30:53:@17852.4]
  wire  valid_55_44; // @[Switch.scala 30:36:@17853.4]
  wire  _T_38964; // @[Switch.scala 30:53:@17855.4]
  wire  valid_55_45; // @[Switch.scala 30:36:@17856.4]
  wire  _T_38967; // @[Switch.scala 30:53:@17858.4]
  wire  valid_55_46; // @[Switch.scala 30:36:@17859.4]
  wire  _T_38970; // @[Switch.scala 30:53:@17861.4]
  wire  valid_55_47; // @[Switch.scala 30:36:@17862.4]
  wire  _T_38973; // @[Switch.scala 30:53:@17864.4]
  wire  valid_55_48; // @[Switch.scala 30:36:@17865.4]
  wire  _T_38976; // @[Switch.scala 30:53:@17867.4]
  wire  valid_55_49; // @[Switch.scala 30:36:@17868.4]
  wire  _T_38979; // @[Switch.scala 30:53:@17870.4]
  wire  valid_55_50; // @[Switch.scala 30:36:@17871.4]
  wire  _T_38982; // @[Switch.scala 30:53:@17873.4]
  wire  valid_55_51; // @[Switch.scala 30:36:@17874.4]
  wire  _T_38985; // @[Switch.scala 30:53:@17876.4]
  wire  valid_55_52; // @[Switch.scala 30:36:@17877.4]
  wire  _T_38988; // @[Switch.scala 30:53:@17879.4]
  wire  valid_55_53; // @[Switch.scala 30:36:@17880.4]
  wire  _T_38991; // @[Switch.scala 30:53:@17882.4]
  wire  valid_55_54; // @[Switch.scala 30:36:@17883.4]
  wire  _T_38994; // @[Switch.scala 30:53:@17885.4]
  wire  valid_55_55; // @[Switch.scala 30:36:@17886.4]
  wire  _T_38997; // @[Switch.scala 30:53:@17888.4]
  wire  valid_55_56; // @[Switch.scala 30:36:@17889.4]
  wire  _T_39000; // @[Switch.scala 30:53:@17891.4]
  wire  valid_55_57; // @[Switch.scala 30:36:@17892.4]
  wire  _T_39003; // @[Switch.scala 30:53:@17894.4]
  wire  valid_55_58; // @[Switch.scala 30:36:@17895.4]
  wire  _T_39006; // @[Switch.scala 30:53:@17897.4]
  wire  valid_55_59; // @[Switch.scala 30:36:@17898.4]
  wire  _T_39009; // @[Switch.scala 30:53:@17900.4]
  wire  valid_55_60; // @[Switch.scala 30:36:@17901.4]
  wire  _T_39012; // @[Switch.scala 30:53:@17903.4]
  wire  valid_55_61; // @[Switch.scala 30:36:@17904.4]
  wire  _T_39015; // @[Switch.scala 30:53:@17906.4]
  wire  valid_55_62; // @[Switch.scala 30:36:@17907.4]
  wire  _T_39018; // @[Switch.scala 30:53:@17909.4]
  wire  valid_55_63; // @[Switch.scala 30:36:@17910.4]
  wire [5:0] _T_39084; // @[Mux.scala 31:69:@17912.4]
  wire [5:0] _T_39085; // @[Mux.scala 31:69:@17913.4]
  wire [5:0] _T_39086; // @[Mux.scala 31:69:@17914.4]
  wire [5:0] _T_39087; // @[Mux.scala 31:69:@17915.4]
  wire [5:0] _T_39088; // @[Mux.scala 31:69:@17916.4]
  wire [5:0] _T_39089; // @[Mux.scala 31:69:@17917.4]
  wire [5:0] _T_39090; // @[Mux.scala 31:69:@17918.4]
  wire [5:0] _T_39091; // @[Mux.scala 31:69:@17919.4]
  wire [5:0] _T_39092; // @[Mux.scala 31:69:@17920.4]
  wire [5:0] _T_39093; // @[Mux.scala 31:69:@17921.4]
  wire [5:0] _T_39094; // @[Mux.scala 31:69:@17922.4]
  wire [5:0] _T_39095; // @[Mux.scala 31:69:@17923.4]
  wire [5:0] _T_39096; // @[Mux.scala 31:69:@17924.4]
  wire [5:0] _T_39097; // @[Mux.scala 31:69:@17925.4]
  wire [5:0] _T_39098; // @[Mux.scala 31:69:@17926.4]
  wire [5:0] _T_39099; // @[Mux.scala 31:69:@17927.4]
  wire [5:0] _T_39100; // @[Mux.scala 31:69:@17928.4]
  wire [5:0] _T_39101; // @[Mux.scala 31:69:@17929.4]
  wire [5:0] _T_39102; // @[Mux.scala 31:69:@17930.4]
  wire [5:0] _T_39103; // @[Mux.scala 31:69:@17931.4]
  wire [5:0] _T_39104; // @[Mux.scala 31:69:@17932.4]
  wire [5:0] _T_39105; // @[Mux.scala 31:69:@17933.4]
  wire [5:0] _T_39106; // @[Mux.scala 31:69:@17934.4]
  wire [5:0] _T_39107; // @[Mux.scala 31:69:@17935.4]
  wire [5:0] _T_39108; // @[Mux.scala 31:69:@17936.4]
  wire [5:0] _T_39109; // @[Mux.scala 31:69:@17937.4]
  wire [5:0] _T_39110; // @[Mux.scala 31:69:@17938.4]
  wire [5:0] _T_39111; // @[Mux.scala 31:69:@17939.4]
  wire [5:0] _T_39112; // @[Mux.scala 31:69:@17940.4]
  wire [5:0] _T_39113; // @[Mux.scala 31:69:@17941.4]
  wire [5:0] _T_39114; // @[Mux.scala 31:69:@17942.4]
  wire [5:0] _T_39115; // @[Mux.scala 31:69:@17943.4]
  wire [5:0] _T_39116; // @[Mux.scala 31:69:@17944.4]
  wire [5:0] _T_39117; // @[Mux.scala 31:69:@17945.4]
  wire [5:0] _T_39118; // @[Mux.scala 31:69:@17946.4]
  wire [5:0] _T_39119; // @[Mux.scala 31:69:@17947.4]
  wire [5:0] _T_39120; // @[Mux.scala 31:69:@17948.4]
  wire [5:0] _T_39121; // @[Mux.scala 31:69:@17949.4]
  wire [5:0] _T_39122; // @[Mux.scala 31:69:@17950.4]
  wire [5:0] _T_39123; // @[Mux.scala 31:69:@17951.4]
  wire [5:0] _T_39124; // @[Mux.scala 31:69:@17952.4]
  wire [5:0] _T_39125; // @[Mux.scala 31:69:@17953.4]
  wire [5:0] _T_39126; // @[Mux.scala 31:69:@17954.4]
  wire [5:0] _T_39127; // @[Mux.scala 31:69:@17955.4]
  wire [5:0] _T_39128; // @[Mux.scala 31:69:@17956.4]
  wire [5:0] _T_39129; // @[Mux.scala 31:69:@17957.4]
  wire [5:0] _T_39130; // @[Mux.scala 31:69:@17958.4]
  wire [5:0] _T_39131; // @[Mux.scala 31:69:@17959.4]
  wire [5:0] _T_39132; // @[Mux.scala 31:69:@17960.4]
  wire [5:0] _T_39133; // @[Mux.scala 31:69:@17961.4]
  wire [5:0] _T_39134; // @[Mux.scala 31:69:@17962.4]
  wire [5:0] _T_39135; // @[Mux.scala 31:69:@17963.4]
  wire [5:0] _T_39136; // @[Mux.scala 31:69:@17964.4]
  wire [5:0] _T_39137; // @[Mux.scala 31:69:@17965.4]
  wire [5:0] _T_39138; // @[Mux.scala 31:69:@17966.4]
  wire [5:0] _T_39139; // @[Mux.scala 31:69:@17967.4]
  wire [5:0] _T_39140; // @[Mux.scala 31:69:@17968.4]
  wire [5:0] _T_39141; // @[Mux.scala 31:69:@17969.4]
  wire [5:0] _T_39142; // @[Mux.scala 31:69:@17970.4]
  wire [5:0] _T_39143; // @[Mux.scala 31:69:@17971.4]
  wire [5:0] _T_39144; // @[Mux.scala 31:69:@17972.4]
  wire [5:0] _T_39145; // @[Mux.scala 31:69:@17973.4]
  wire [5:0] select_55; // @[Mux.scala 31:69:@17974.4]
  wire [47:0] _GEN_3521; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3522; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3523; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3524; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3525; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3526; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3527; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3528; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3529; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3530; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3531; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3532; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3533; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3534; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3535; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3536; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3537; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3538; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3539; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3540; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3541; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3542; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3543; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3544; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3545; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3546; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3547; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3548; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3549; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3550; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3551; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3552; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3553; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3554; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3555; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3556; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3557; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3558; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3559; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3560; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3561; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3562; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3563; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3564; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3565; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3566; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3567; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3568; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3569; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3570; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3571; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3572; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3573; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3574; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3575; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3576; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3577; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3578; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3579; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3580; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3581; // @[Switch.scala 33:19:@17976.4]
  wire [47:0] _GEN_3582; // @[Switch.scala 33:19:@17976.4]
  wire [7:0] _T_39154; // @[Switch.scala 34:32:@17983.4]
  wire [15:0] _T_39162; // @[Switch.scala 34:32:@17991.4]
  wire [7:0] _T_39169; // @[Switch.scala 34:32:@17998.4]
  wire [31:0] _T_39178; // @[Switch.scala 34:32:@18007.4]
  wire [7:0] _T_39185; // @[Switch.scala 34:32:@18014.4]
  wire [15:0] _T_39193; // @[Switch.scala 34:32:@18022.4]
  wire [7:0] _T_39200; // @[Switch.scala 34:32:@18029.4]
  wire [31:0] _T_39209; // @[Switch.scala 34:32:@18038.4]
  wire [63:0] _T_39210; // @[Switch.scala 34:32:@18039.4]
  wire  _T_39214; // @[Switch.scala 30:53:@18042.4]
  wire  valid_56_0; // @[Switch.scala 30:36:@18043.4]
  wire  _T_39217; // @[Switch.scala 30:53:@18045.4]
  wire  valid_56_1; // @[Switch.scala 30:36:@18046.4]
  wire  _T_39220; // @[Switch.scala 30:53:@18048.4]
  wire  valid_56_2; // @[Switch.scala 30:36:@18049.4]
  wire  _T_39223; // @[Switch.scala 30:53:@18051.4]
  wire  valid_56_3; // @[Switch.scala 30:36:@18052.4]
  wire  _T_39226; // @[Switch.scala 30:53:@18054.4]
  wire  valid_56_4; // @[Switch.scala 30:36:@18055.4]
  wire  _T_39229; // @[Switch.scala 30:53:@18057.4]
  wire  valid_56_5; // @[Switch.scala 30:36:@18058.4]
  wire  _T_39232; // @[Switch.scala 30:53:@18060.4]
  wire  valid_56_6; // @[Switch.scala 30:36:@18061.4]
  wire  _T_39235; // @[Switch.scala 30:53:@18063.4]
  wire  valid_56_7; // @[Switch.scala 30:36:@18064.4]
  wire  _T_39238; // @[Switch.scala 30:53:@18066.4]
  wire  valid_56_8; // @[Switch.scala 30:36:@18067.4]
  wire  _T_39241; // @[Switch.scala 30:53:@18069.4]
  wire  valid_56_9; // @[Switch.scala 30:36:@18070.4]
  wire  _T_39244; // @[Switch.scala 30:53:@18072.4]
  wire  valid_56_10; // @[Switch.scala 30:36:@18073.4]
  wire  _T_39247; // @[Switch.scala 30:53:@18075.4]
  wire  valid_56_11; // @[Switch.scala 30:36:@18076.4]
  wire  _T_39250; // @[Switch.scala 30:53:@18078.4]
  wire  valid_56_12; // @[Switch.scala 30:36:@18079.4]
  wire  _T_39253; // @[Switch.scala 30:53:@18081.4]
  wire  valid_56_13; // @[Switch.scala 30:36:@18082.4]
  wire  _T_39256; // @[Switch.scala 30:53:@18084.4]
  wire  valid_56_14; // @[Switch.scala 30:36:@18085.4]
  wire  _T_39259; // @[Switch.scala 30:53:@18087.4]
  wire  valid_56_15; // @[Switch.scala 30:36:@18088.4]
  wire  _T_39262; // @[Switch.scala 30:53:@18090.4]
  wire  valid_56_16; // @[Switch.scala 30:36:@18091.4]
  wire  _T_39265; // @[Switch.scala 30:53:@18093.4]
  wire  valid_56_17; // @[Switch.scala 30:36:@18094.4]
  wire  _T_39268; // @[Switch.scala 30:53:@18096.4]
  wire  valid_56_18; // @[Switch.scala 30:36:@18097.4]
  wire  _T_39271; // @[Switch.scala 30:53:@18099.4]
  wire  valid_56_19; // @[Switch.scala 30:36:@18100.4]
  wire  _T_39274; // @[Switch.scala 30:53:@18102.4]
  wire  valid_56_20; // @[Switch.scala 30:36:@18103.4]
  wire  _T_39277; // @[Switch.scala 30:53:@18105.4]
  wire  valid_56_21; // @[Switch.scala 30:36:@18106.4]
  wire  _T_39280; // @[Switch.scala 30:53:@18108.4]
  wire  valid_56_22; // @[Switch.scala 30:36:@18109.4]
  wire  _T_39283; // @[Switch.scala 30:53:@18111.4]
  wire  valid_56_23; // @[Switch.scala 30:36:@18112.4]
  wire  _T_39286; // @[Switch.scala 30:53:@18114.4]
  wire  valid_56_24; // @[Switch.scala 30:36:@18115.4]
  wire  _T_39289; // @[Switch.scala 30:53:@18117.4]
  wire  valid_56_25; // @[Switch.scala 30:36:@18118.4]
  wire  _T_39292; // @[Switch.scala 30:53:@18120.4]
  wire  valid_56_26; // @[Switch.scala 30:36:@18121.4]
  wire  _T_39295; // @[Switch.scala 30:53:@18123.4]
  wire  valid_56_27; // @[Switch.scala 30:36:@18124.4]
  wire  _T_39298; // @[Switch.scala 30:53:@18126.4]
  wire  valid_56_28; // @[Switch.scala 30:36:@18127.4]
  wire  _T_39301; // @[Switch.scala 30:53:@18129.4]
  wire  valid_56_29; // @[Switch.scala 30:36:@18130.4]
  wire  _T_39304; // @[Switch.scala 30:53:@18132.4]
  wire  valid_56_30; // @[Switch.scala 30:36:@18133.4]
  wire  _T_39307; // @[Switch.scala 30:53:@18135.4]
  wire  valid_56_31; // @[Switch.scala 30:36:@18136.4]
  wire  _T_39310; // @[Switch.scala 30:53:@18138.4]
  wire  valid_56_32; // @[Switch.scala 30:36:@18139.4]
  wire  _T_39313; // @[Switch.scala 30:53:@18141.4]
  wire  valid_56_33; // @[Switch.scala 30:36:@18142.4]
  wire  _T_39316; // @[Switch.scala 30:53:@18144.4]
  wire  valid_56_34; // @[Switch.scala 30:36:@18145.4]
  wire  _T_39319; // @[Switch.scala 30:53:@18147.4]
  wire  valid_56_35; // @[Switch.scala 30:36:@18148.4]
  wire  _T_39322; // @[Switch.scala 30:53:@18150.4]
  wire  valid_56_36; // @[Switch.scala 30:36:@18151.4]
  wire  _T_39325; // @[Switch.scala 30:53:@18153.4]
  wire  valid_56_37; // @[Switch.scala 30:36:@18154.4]
  wire  _T_39328; // @[Switch.scala 30:53:@18156.4]
  wire  valid_56_38; // @[Switch.scala 30:36:@18157.4]
  wire  _T_39331; // @[Switch.scala 30:53:@18159.4]
  wire  valid_56_39; // @[Switch.scala 30:36:@18160.4]
  wire  _T_39334; // @[Switch.scala 30:53:@18162.4]
  wire  valid_56_40; // @[Switch.scala 30:36:@18163.4]
  wire  _T_39337; // @[Switch.scala 30:53:@18165.4]
  wire  valid_56_41; // @[Switch.scala 30:36:@18166.4]
  wire  _T_39340; // @[Switch.scala 30:53:@18168.4]
  wire  valid_56_42; // @[Switch.scala 30:36:@18169.4]
  wire  _T_39343; // @[Switch.scala 30:53:@18171.4]
  wire  valid_56_43; // @[Switch.scala 30:36:@18172.4]
  wire  _T_39346; // @[Switch.scala 30:53:@18174.4]
  wire  valid_56_44; // @[Switch.scala 30:36:@18175.4]
  wire  _T_39349; // @[Switch.scala 30:53:@18177.4]
  wire  valid_56_45; // @[Switch.scala 30:36:@18178.4]
  wire  _T_39352; // @[Switch.scala 30:53:@18180.4]
  wire  valid_56_46; // @[Switch.scala 30:36:@18181.4]
  wire  _T_39355; // @[Switch.scala 30:53:@18183.4]
  wire  valid_56_47; // @[Switch.scala 30:36:@18184.4]
  wire  _T_39358; // @[Switch.scala 30:53:@18186.4]
  wire  valid_56_48; // @[Switch.scala 30:36:@18187.4]
  wire  _T_39361; // @[Switch.scala 30:53:@18189.4]
  wire  valid_56_49; // @[Switch.scala 30:36:@18190.4]
  wire  _T_39364; // @[Switch.scala 30:53:@18192.4]
  wire  valid_56_50; // @[Switch.scala 30:36:@18193.4]
  wire  _T_39367; // @[Switch.scala 30:53:@18195.4]
  wire  valid_56_51; // @[Switch.scala 30:36:@18196.4]
  wire  _T_39370; // @[Switch.scala 30:53:@18198.4]
  wire  valid_56_52; // @[Switch.scala 30:36:@18199.4]
  wire  _T_39373; // @[Switch.scala 30:53:@18201.4]
  wire  valid_56_53; // @[Switch.scala 30:36:@18202.4]
  wire  _T_39376; // @[Switch.scala 30:53:@18204.4]
  wire  valid_56_54; // @[Switch.scala 30:36:@18205.4]
  wire  _T_39379; // @[Switch.scala 30:53:@18207.4]
  wire  valid_56_55; // @[Switch.scala 30:36:@18208.4]
  wire  _T_39382; // @[Switch.scala 30:53:@18210.4]
  wire  valid_56_56; // @[Switch.scala 30:36:@18211.4]
  wire  _T_39385; // @[Switch.scala 30:53:@18213.4]
  wire  valid_56_57; // @[Switch.scala 30:36:@18214.4]
  wire  _T_39388; // @[Switch.scala 30:53:@18216.4]
  wire  valid_56_58; // @[Switch.scala 30:36:@18217.4]
  wire  _T_39391; // @[Switch.scala 30:53:@18219.4]
  wire  valid_56_59; // @[Switch.scala 30:36:@18220.4]
  wire  _T_39394; // @[Switch.scala 30:53:@18222.4]
  wire  valid_56_60; // @[Switch.scala 30:36:@18223.4]
  wire  _T_39397; // @[Switch.scala 30:53:@18225.4]
  wire  valid_56_61; // @[Switch.scala 30:36:@18226.4]
  wire  _T_39400; // @[Switch.scala 30:53:@18228.4]
  wire  valid_56_62; // @[Switch.scala 30:36:@18229.4]
  wire  _T_39403; // @[Switch.scala 30:53:@18231.4]
  wire  valid_56_63; // @[Switch.scala 30:36:@18232.4]
  wire [5:0] _T_39469; // @[Mux.scala 31:69:@18234.4]
  wire [5:0] _T_39470; // @[Mux.scala 31:69:@18235.4]
  wire [5:0] _T_39471; // @[Mux.scala 31:69:@18236.4]
  wire [5:0] _T_39472; // @[Mux.scala 31:69:@18237.4]
  wire [5:0] _T_39473; // @[Mux.scala 31:69:@18238.4]
  wire [5:0] _T_39474; // @[Mux.scala 31:69:@18239.4]
  wire [5:0] _T_39475; // @[Mux.scala 31:69:@18240.4]
  wire [5:0] _T_39476; // @[Mux.scala 31:69:@18241.4]
  wire [5:0] _T_39477; // @[Mux.scala 31:69:@18242.4]
  wire [5:0] _T_39478; // @[Mux.scala 31:69:@18243.4]
  wire [5:0] _T_39479; // @[Mux.scala 31:69:@18244.4]
  wire [5:0] _T_39480; // @[Mux.scala 31:69:@18245.4]
  wire [5:0] _T_39481; // @[Mux.scala 31:69:@18246.4]
  wire [5:0] _T_39482; // @[Mux.scala 31:69:@18247.4]
  wire [5:0] _T_39483; // @[Mux.scala 31:69:@18248.4]
  wire [5:0] _T_39484; // @[Mux.scala 31:69:@18249.4]
  wire [5:0] _T_39485; // @[Mux.scala 31:69:@18250.4]
  wire [5:0] _T_39486; // @[Mux.scala 31:69:@18251.4]
  wire [5:0] _T_39487; // @[Mux.scala 31:69:@18252.4]
  wire [5:0] _T_39488; // @[Mux.scala 31:69:@18253.4]
  wire [5:0] _T_39489; // @[Mux.scala 31:69:@18254.4]
  wire [5:0] _T_39490; // @[Mux.scala 31:69:@18255.4]
  wire [5:0] _T_39491; // @[Mux.scala 31:69:@18256.4]
  wire [5:0] _T_39492; // @[Mux.scala 31:69:@18257.4]
  wire [5:0] _T_39493; // @[Mux.scala 31:69:@18258.4]
  wire [5:0] _T_39494; // @[Mux.scala 31:69:@18259.4]
  wire [5:0] _T_39495; // @[Mux.scala 31:69:@18260.4]
  wire [5:0] _T_39496; // @[Mux.scala 31:69:@18261.4]
  wire [5:0] _T_39497; // @[Mux.scala 31:69:@18262.4]
  wire [5:0] _T_39498; // @[Mux.scala 31:69:@18263.4]
  wire [5:0] _T_39499; // @[Mux.scala 31:69:@18264.4]
  wire [5:0] _T_39500; // @[Mux.scala 31:69:@18265.4]
  wire [5:0] _T_39501; // @[Mux.scala 31:69:@18266.4]
  wire [5:0] _T_39502; // @[Mux.scala 31:69:@18267.4]
  wire [5:0] _T_39503; // @[Mux.scala 31:69:@18268.4]
  wire [5:0] _T_39504; // @[Mux.scala 31:69:@18269.4]
  wire [5:0] _T_39505; // @[Mux.scala 31:69:@18270.4]
  wire [5:0] _T_39506; // @[Mux.scala 31:69:@18271.4]
  wire [5:0] _T_39507; // @[Mux.scala 31:69:@18272.4]
  wire [5:0] _T_39508; // @[Mux.scala 31:69:@18273.4]
  wire [5:0] _T_39509; // @[Mux.scala 31:69:@18274.4]
  wire [5:0] _T_39510; // @[Mux.scala 31:69:@18275.4]
  wire [5:0] _T_39511; // @[Mux.scala 31:69:@18276.4]
  wire [5:0] _T_39512; // @[Mux.scala 31:69:@18277.4]
  wire [5:0] _T_39513; // @[Mux.scala 31:69:@18278.4]
  wire [5:0] _T_39514; // @[Mux.scala 31:69:@18279.4]
  wire [5:0] _T_39515; // @[Mux.scala 31:69:@18280.4]
  wire [5:0] _T_39516; // @[Mux.scala 31:69:@18281.4]
  wire [5:0] _T_39517; // @[Mux.scala 31:69:@18282.4]
  wire [5:0] _T_39518; // @[Mux.scala 31:69:@18283.4]
  wire [5:0] _T_39519; // @[Mux.scala 31:69:@18284.4]
  wire [5:0] _T_39520; // @[Mux.scala 31:69:@18285.4]
  wire [5:0] _T_39521; // @[Mux.scala 31:69:@18286.4]
  wire [5:0] _T_39522; // @[Mux.scala 31:69:@18287.4]
  wire [5:0] _T_39523; // @[Mux.scala 31:69:@18288.4]
  wire [5:0] _T_39524; // @[Mux.scala 31:69:@18289.4]
  wire [5:0] _T_39525; // @[Mux.scala 31:69:@18290.4]
  wire [5:0] _T_39526; // @[Mux.scala 31:69:@18291.4]
  wire [5:0] _T_39527; // @[Mux.scala 31:69:@18292.4]
  wire [5:0] _T_39528; // @[Mux.scala 31:69:@18293.4]
  wire [5:0] _T_39529; // @[Mux.scala 31:69:@18294.4]
  wire [5:0] _T_39530; // @[Mux.scala 31:69:@18295.4]
  wire [5:0] select_56; // @[Mux.scala 31:69:@18296.4]
  wire [47:0] _GEN_3585; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3586; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3587; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3588; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3589; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3590; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3591; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3592; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3593; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3594; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3595; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3596; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3597; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3598; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3599; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3600; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3601; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3602; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3603; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3604; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3605; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3606; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3607; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3608; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3609; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3610; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3611; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3612; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3613; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3614; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3615; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3616; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3617; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3618; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3619; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3620; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3621; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3622; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3623; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3624; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3625; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3626; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3627; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3628; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3629; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3630; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3631; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3632; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3633; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3634; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3635; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3636; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3637; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3638; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3639; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3640; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3641; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3642; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3643; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3644; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3645; // @[Switch.scala 33:19:@18298.4]
  wire [47:0] _GEN_3646; // @[Switch.scala 33:19:@18298.4]
  wire [7:0] _T_39539; // @[Switch.scala 34:32:@18305.4]
  wire [15:0] _T_39547; // @[Switch.scala 34:32:@18313.4]
  wire [7:0] _T_39554; // @[Switch.scala 34:32:@18320.4]
  wire [31:0] _T_39563; // @[Switch.scala 34:32:@18329.4]
  wire [7:0] _T_39570; // @[Switch.scala 34:32:@18336.4]
  wire [15:0] _T_39578; // @[Switch.scala 34:32:@18344.4]
  wire [7:0] _T_39585; // @[Switch.scala 34:32:@18351.4]
  wire [31:0] _T_39594; // @[Switch.scala 34:32:@18360.4]
  wire [63:0] _T_39595; // @[Switch.scala 34:32:@18361.4]
  wire  _T_39599; // @[Switch.scala 30:53:@18364.4]
  wire  valid_57_0; // @[Switch.scala 30:36:@18365.4]
  wire  _T_39602; // @[Switch.scala 30:53:@18367.4]
  wire  valid_57_1; // @[Switch.scala 30:36:@18368.4]
  wire  _T_39605; // @[Switch.scala 30:53:@18370.4]
  wire  valid_57_2; // @[Switch.scala 30:36:@18371.4]
  wire  _T_39608; // @[Switch.scala 30:53:@18373.4]
  wire  valid_57_3; // @[Switch.scala 30:36:@18374.4]
  wire  _T_39611; // @[Switch.scala 30:53:@18376.4]
  wire  valid_57_4; // @[Switch.scala 30:36:@18377.4]
  wire  _T_39614; // @[Switch.scala 30:53:@18379.4]
  wire  valid_57_5; // @[Switch.scala 30:36:@18380.4]
  wire  _T_39617; // @[Switch.scala 30:53:@18382.4]
  wire  valid_57_6; // @[Switch.scala 30:36:@18383.4]
  wire  _T_39620; // @[Switch.scala 30:53:@18385.4]
  wire  valid_57_7; // @[Switch.scala 30:36:@18386.4]
  wire  _T_39623; // @[Switch.scala 30:53:@18388.4]
  wire  valid_57_8; // @[Switch.scala 30:36:@18389.4]
  wire  _T_39626; // @[Switch.scala 30:53:@18391.4]
  wire  valid_57_9; // @[Switch.scala 30:36:@18392.4]
  wire  _T_39629; // @[Switch.scala 30:53:@18394.4]
  wire  valid_57_10; // @[Switch.scala 30:36:@18395.4]
  wire  _T_39632; // @[Switch.scala 30:53:@18397.4]
  wire  valid_57_11; // @[Switch.scala 30:36:@18398.4]
  wire  _T_39635; // @[Switch.scala 30:53:@18400.4]
  wire  valid_57_12; // @[Switch.scala 30:36:@18401.4]
  wire  _T_39638; // @[Switch.scala 30:53:@18403.4]
  wire  valid_57_13; // @[Switch.scala 30:36:@18404.4]
  wire  _T_39641; // @[Switch.scala 30:53:@18406.4]
  wire  valid_57_14; // @[Switch.scala 30:36:@18407.4]
  wire  _T_39644; // @[Switch.scala 30:53:@18409.4]
  wire  valid_57_15; // @[Switch.scala 30:36:@18410.4]
  wire  _T_39647; // @[Switch.scala 30:53:@18412.4]
  wire  valid_57_16; // @[Switch.scala 30:36:@18413.4]
  wire  _T_39650; // @[Switch.scala 30:53:@18415.4]
  wire  valid_57_17; // @[Switch.scala 30:36:@18416.4]
  wire  _T_39653; // @[Switch.scala 30:53:@18418.4]
  wire  valid_57_18; // @[Switch.scala 30:36:@18419.4]
  wire  _T_39656; // @[Switch.scala 30:53:@18421.4]
  wire  valid_57_19; // @[Switch.scala 30:36:@18422.4]
  wire  _T_39659; // @[Switch.scala 30:53:@18424.4]
  wire  valid_57_20; // @[Switch.scala 30:36:@18425.4]
  wire  _T_39662; // @[Switch.scala 30:53:@18427.4]
  wire  valid_57_21; // @[Switch.scala 30:36:@18428.4]
  wire  _T_39665; // @[Switch.scala 30:53:@18430.4]
  wire  valid_57_22; // @[Switch.scala 30:36:@18431.4]
  wire  _T_39668; // @[Switch.scala 30:53:@18433.4]
  wire  valid_57_23; // @[Switch.scala 30:36:@18434.4]
  wire  _T_39671; // @[Switch.scala 30:53:@18436.4]
  wire  valid_57_24; // @[Switch.scala 30:36:@18437.4]
  wire  _T_39674; // @[Switch.scala 30:53:@18439.4]
  wire  valid_57_25; // @[Switch.scala 30:36:@18440.4]
  wire  _T_39677; // @[Switch.scala 30:53:@18442.4]
  wire  valid_57_26; // @[Switch.scala 30:36:@18443.4]
  wire  _T_39680; // @[Switch.scala 30:53:@18445.4]
  wire  valid_57_27; // @[Switch.scala 30:36:@18446.4]
  wire  _T_39683; // @[Switch.scala 30:53:@18448.4]
  wire  valid_57_28; // @[Switch.scala 30:36:@18449.4]
  wire  _T_39686; // @[Switch.scala 30:53:@18451.4]
  wire  valid_57_29; // @[Switch.scala 30:36:@18452.4]
  wire  _T_39689; // @[Switch.scala 30:53:@18454.4]
  wire  valid_57_30; // @[Switch.scala 30:36:@18455.4]
  wire  _T_39692; // @[Switch.scala 30:53:@18457.4]
  wire  valid_57_31; // @[Switch.scala 30:36:@18458.4]
  wire  _T_39695; // @[Switch.scala 30:53:@18460.4]
  wire  valid_57_32; // @[Switch.scala 30:36:@18461.4]
  wire  _T_39698; // @[Switch.scala 30:53:@18463.4]
  wire  valid_57_33; // @[Switch.scala 30:36:@18464.4]
  wire  _T_39701; // @[Switch.scala 30:53:@18466.4]
  wire  valid_57_34; // @[Switch.scala 30:36:@18467.4]
  wire  _T_39704; // @[Switch.scala 30:53:@18469.4]
  wire  valid_57_35; // @[Switch.scala 30:36:@18470.4]
  wire  _T_39707; // @[Switch.scala 30:53:@18472.4]
  wire  valid_57_36; // @[Switch.scala 30:36:@18473.4]
  wire  _T_39710; // @[Switch.scala 30:53:@18475.4]
  wire  valid_57_37; // @[Switch.scala 30:36:@18476.4]
  wire  _T_39713; // @[Switch.scala 30:53:@18478.4]
  wire  valid_57_38; // @[Switch.scala 30:36:@18479.4]
  wire  _T_39716; // @[Switch.scala 30:53:@18481.4]
  wire  valid_57_39; // @[Switch.scala 30:36:@18482.4]
  wire  _T_39719; // @[Switch.scala 30:53:@18484.4]
  wire  valid_57_40; // @[Switch.scala 30:36:@18485.4]
  wire  _T_39722; // @[Switch.scala 30:53:@18487.4]
  wire  valid_57_41; // @[Switch.scala 30:36:@18488.4]
  wire  _T_39725; // @[Switch.scala 30:53:@18490.4]
  wire  valid_57_42; // @[Switch.scala 30:36:@18491.4]
  wire  _T_39728; // @[Switch.scala 30:53:@18493.4]
  wire  valid_57_43; // @[Switch.scala 30:36:@18494.4]
  wire  _T_39731; // @[Switch.scala 30:53:@18496.4]
  wire  valid_57_44; // @[Switch.scala 30:36:@18497.4]
  wire  _T_39734; // @[Switch.scala 30:53:@18499.4]
  wire  valid_57_45; // @[Switch.scala 30:36:@18500.4]
  wire  _T_39737; // @[Switch.scala 30:53:@18502.4]
  wire  valid_57_46; // @[Switch.scala 30:36:@18503.4]
  wire  _T_39740; // @[Switch.scala 30:53:@18505.4]
  wire  valid_57_47; // @[Switch.scala 30:36:@18506.4]
  wire  _T_39743; // @[Switch.scala 30:53:@18508.4]
  wire  valid_57_48; // @[Switch.scala 30:36:@18509.4]
  wire  _T_39746; // @[Switch.scala 30:53:@18511.4]
  wire  valid_57_49; // @[Switch.scala 30:36:@18512.4]
  wire  _T_39749; // @[Switch.scala 30:53:@18514.4]
  wire  valid_57_50; // @[Switch.scala 30:36:@18515.4]
  wire  _T_39752; // @[Switch.scala 30:53:@18517.4]
  wire  valid_57_51; // @[Switch.scala 30:36:@18518.4]
  wire  _T_39755; // @[Switch.scala 30:53:@18520.4]
  wire  valid_57_52; // @[Switch.scala 30:36:@18521.4]
  wire  _T_39758; // @[Switch.scala 30:53:@18523.4]
  wire  valid_57_53; // @[Switch.scala 30:36:@18524.4]
  wire  _T_39761; // @[Switch.scala 30:53:@18526.4]
  wire  valid_57_54; // @[Switch.scala 30:36:@18527.4]
  wire  _T_39764; // @[Switch.scala 30:53:@18529.4]
  wire  valid_57_55; // @[Switch.scala 30:36:@18530.4]
  wire  _T_39767; // @[Switch.scala 30:53:@18532.4]
  wire  valid_57_56; // @[Switch.scala 30:36:@18533.4]
  wire  _T_39770; // @[Switch.scala 30:53:@18535.4]
  wire  valid_57_57; // @[Switch.scala 30:36:@18536.4]
  wire  _T_39773; // @[Switch.scala 30:53:@18538.4]
  wire  valid_57_58; // @[Switch.scala 30:36:@18539.4]
  wire  _T_39776; // @[Switch.scala 30:53:@18541.4]
  wire  valid_57_59; // @[Switch.scala 30:36:@18542.4]
  wire  _T_39779; // @[Switch.scala 30:53:@18544.4]
  wire  valid_57_60; // @[Switch.scala 30:36:@18545.4]
  wire  _T_39782; // @[Switch.scala 30:53:@18547.4]
  wire  valid_57_61; // @[Switch.scala 30:36:@18548.4]
  wire  _T_39785; // @[Switch.scala 30:53:@18550.4]
  wire  valid_57_62; // @[Switch.scala 30:36:@18551.4]
  wire  _T_39788; // @[Switch.scala 30:53:@18553.4]
  wire  valid_57_63; // @[Switch.scala 30:36:@18554.4]
  wire [5:0] _T_39854; // @[Mux.scala 31:69:@18556.4]
  wire [5:0] _T_39855; // @[Mux.scala 31:69:@18557.4]
  wire [5:0] _T_39856; // @[Mux.scala 31:69:@18558.4]
  wire [5:0] _T_39857; // @[Mux.scala 31:69:@18559.4]
  wire [5:0] _T_39858; // @[Mux.scala 31:69:@18560.4]
  wire [5:0] _T_39859; // @[Mux.scala 31:69:@18561.4]
  wire [5:0] _T_39860; // @[Mux.scala 31:69:@18562.4]
  wire [5:0] _T_39861; // @[Mux.scala 31:69:@18563.4]
  wire [5:0] _T_39862; // @[Mux.scala 31:69:@18564.4]
  wire [5:0] _T_39863; // @[Mux.scala 31:69:@18565.4]
  wire [5:0] _T_39864; // @[Mux.scala 31:69:@18566.4]
  wire [5:0] _T_39865; // @[Mux.scala 31:69:@18567.4]
  wire [5:0] _T_39866; // @[Mux.scala 31:69:@18568.4]
  wire [5:0] _T_39867; // @[Mux.scala 31:69:@18569.4]
  wire [5:0] _T_39868; // @[Mux.scala 31:69:@18570.4]
  wire [5:0] _T_39869; // @[Mux.scala 31:69:@18571.4]
  wire [5:0] _T_39870; // @[Mux.scala 31:69:@18572.4]
  wire [5:0] _T_39871; // @[Mux.scala 31:69:@18573.4]
  wire [5:0] _T_39872; // @[Mux.scala 31:69:@18574.4]
  wire [5:0] _T_39873; // @[Mux.scala 31:69:@18575.4]
  wire [5:0] _T_39874; // @[Mux.scala 31:69:@18576.4]
  wire [5:0] _T_39875; // @[Mux.scala 31:69:@18577.4]
  wire [5:0] _T_39876; // @[Mux.scala 31:69:@18578.4]
  wire [5:0] _T_39877; // @[Mux.scala 31:69:@18579.4]
  wire [5:0] _T_39878; // @[Mux.scala 31:69:@18580.4]
  wire [5:0] _T_39879; // @[Mux.scala 31:69:@18581.4]
  wire [5:0] _T_39880; // @[Mux.scala 31:69:@18582.4]
  wire [5:0] _T_39881; // @[Mux.scala 31:69:@18583.4]
  wire [5:0] _T_39882; // @[Mux.scala 31:69:@18584.4]
  wire [5:0] _T_39883; // @[Mux.scala 31:69:@18585.4]
  wire [5:0] _T_39884; // @[Mux.scala 31:69:@18586.4]
  wire [5:0] _T_39885; // @[Mux.scala 31:69:@18587.4]
  wire [5:0] _T_39886; // @[Mux.scala 31:69:@18588.4]
  wire [5:0] _T_39887; // @[Mux.scala 31:69:@18589.4]
  wire [5:0] _T_39888; // @[Mux.scala 31:69:@18590.4]
  wire [5:0] _T_39889; // @[Mux.scala 31:69:@18591.4]
  wire [5:0] _T_39890; // @[Mux.scala 31:69:@18592.4]
  wire [5:0] _T_39891; // @[Mux.scala 31:69:@18593.4]
  wire [5:0] _T_39892; // @[Mux.scala 31:69:@18594.4]
  wire [5:0] _T_39893; // @[Mux.scala 31:69:@18595.4]
  wire [5:0] _T_39894; // @[Mux.scala 31:69:@18596.4]
  wire [5:0] _T_39895; // @[Mux.scala 31:69:@18597.4]
  wire [5:0] _T_39896; // @[Mux.scala 31:69:@18598.4]
  wire [5:0] _T_39897; // @[Mux.scala 31:69:@18599.4]
  wire [5:0] _T_39898; // @[Mux.scala 31:69:@18600.4]
  wire [5:0] _T_39899; // @[Mux.scala 31:69:@18601.4]
  wire [5:0] _T_39900; // @[Mux.scala 31:69:@18602.4]
  wire [5:0] _T_39901; // @[Mux.scala 31:69:@18603.4]
  wire [5:0] _T_39902; // @[Mux.scala 31:69:@18604.4]
  wire [5:0] _T_39903; // @[Mux.scala 31:69:@18605.4]
  wire [5:0] _T_39904; // @[Mux.scala 31:69:@18606.4]
  wire [5:0] _T_39905; // @[Mux.scala 31:69:@18607.4]
  wire [5:0] _T_39906; // @[Mux.scala 31:69:@18608.4]
  wire [5:0] _T_39907; // @[Mux.scala 31:69:@18609.4]
  wire [5:0] _T_39908; // @[Mux.scala 31:69:@18610.4]
  wire [5:0] _T_39909; // @[Mux.scala 31:69:@18611.4]
  wire [5:0] _T_39910; // @[Mux.scala 31:69:@18612.4]
  wire [5:0] _T_39911; // @[Mux.scala 31:69:@18613.4]
  wire [5:0] _T_39912; // @[Mux.scala 31:69:@18614.4]
  wire [5:0] _T_39913; // @[Mux.scala 31:69:@18615.4]
  wire [5:0] _T_39914; // @[Mux.scala 31:69:@18616.4]
  wire [5:0] _T_39915; // @[Mux.scala 31:69:@18617.4]
  wire [5:0] select_57; // @[Mux.scala 31:69:@18618.4]
  wire [47:0] _GEN_3649; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3650; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3651; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3652; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3653; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3654; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3655; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3656; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3657; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3658; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3659; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3660; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3661; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3662; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3663; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3664; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3665; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3666; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3667; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3668; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3669; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3670; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3671; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3672; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3673; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3674; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3675; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3676; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3677; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3678; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3679; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3680; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3681; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3682; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3683; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3684; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3685; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3686; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3687; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3688; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3689; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3690; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3691; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3692; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3693; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3694; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3695; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3696; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3697; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3698; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3699; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3700; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3701; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3702; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3703; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3704; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3705; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3706; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3707; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3708; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3709; // @[Switch.scala 33:19:@18620.4]
  wire [47:0] _GEN_3710; // @[Switch.scala 33:19:@18620.4]
  wire [7:0] _T_39924; // @[Switch.scala 34:32:@18627.4]
  wire [15:0] _T_39932; // @[Switch.scala 34:32:@18635.4]
  wire [7:0] _T_39939; // @[Switch.scala 34:32:@18642.4]
  wire [31:0] _T_39948; // @[Switch.scala 34:32:@18651.4]
  wire [7:0] _T_39955; // @[Switch.scala 34:32:@18658.4]
  wire [15:0] _T_39963; // @[Switch.scala 34:32:@18666.4]
  wire [7:0] _T_39970; // @[Switch.scala 34:32:@18673.4]
  wire [31:0] _T_39979; // @[Switch.scala 34:32:@18682.4]
  wire [63:0] _T_39980; // @[Switch.scala 34:32:@18683.4]
  wire  _T_39984; // @[Switch.scala 30:53:@18686.4]
  wire  valid_58_0; // @[Switch.scala 30:36:@18687.4]
  wire  _T_39987; // @[Switch.scala 30:53:@18689.4]
  wire  valid_58_1; // @[Switch.scala 30:36:@18690.4]
  wire  _T_39990; // @[Switch.scala 30:53:@18692.4]
  wire  valid_58_2; // @[Switch.scala 30:36:@18693.4]
  wire  _T_39993; // @[Switch.scala 30:53:@18695.4]
  wire  valid_58_3; // @[Switch.scala 30:36:@18696.4]
  wire  _T_39996; // @[Switch.scala 30:53:@18698.4]
  wire  valid_58_4; // @[Switch.scala 30:36:@18699.4]
  wire  _T_39999; // @[Switch.scala 30:53:@18701.4]
  wire  valid_58_5; // @[Switch.scala 30:36:@18702.4]
  wire  _T_40002; // @[Switch.scala 30:53:@18704.4]
  wire  valid_58_6; // @[Switch.scala 30:36:@18705.4]
  wire  _T_40005; // @[Switch.scala 30:53:@18707.4]
  wire  valid_58_7; // @[Switch.scala 30:36:@18708.4]
  wire  _T_40008; // @[Switch.scala 30:53:@18710.4]
  wire  valid_58_8; // @[Switch.scala 30:36:@18711.4]
  wire  _T_40011; // @[Switch.scala 30:53:@18713.4]
  wire  valid_58_9; // @[Switch.scala 30:36:@18714.4]
  wire  _T_40014; // @[Switch.scala 30:53:@18716.4]
  wire  valid_58_10; // @[Switch.scala 30:36:@18717.4]
  wire  _T_40017; // @[Switch.scala 30:53:@18719.4]
  wire  valid_58_11; // @[Switch.scala 30:36:@18720.4]
  wire  _T_40020; // @[Switch.scala 30:53:@18722.4]
  wire  valid_58_12; // @[Switch.scala 30:36:@18723.4]
  wire  _T_40023; // @[Switch.scala 30:53:@18725.4]
  wire  valid_58_13; // @[Switch.scala 30:36:@18726.4]
  wire  _T_40026; // @[Switch.scala 30:53:@18728.4]
  wire  valid_58_14; // @[Switch.scala 30:36:@18729.4]
  wire  _T_40029; // @[Switch.scala 30:53:@18731.4]
  wire  valid_58_15; // @[Switch.scala 30:36:@18732.4]
  wire  _T_40032; // @[Switch.scala 30:53:@18734.4]
  wire  valid_58_16; // @[Switch.scala 30:36:@18735.4]
  wire  _T_40035; // @[Switch.scala 30:53:@18737.4]
  wire  valid_58_17; // @[Switch.scala 30:36:@18738.4]
  wire  _T_40038; // @[Switch.scala 30:53:@18740.4]
  wire  valid_58_18; // @[Switch.scala 30:36:@18741.4]
  wire  _T_40041; // @[Switch.scala 30:53:@18743.4]
  wire  valid_58_19; // @[Switch.scala 30:36:@18744.4]
  wire  _T_40044; // @[Switch.scala 30:53:@18746.4]
  wire  valid_58_20; // @[Switch.scala 30:36:@18747.4]
  wire  _T_40047; // @[Switch.scala 30:53:@18749.4]
  wire  valid_58_21; // @[Switch.scala 30:36:@18750.4]
  wire  _T_40050; // @[Switch.scala 30:53:@18752.4]
  wire  valid_58_22; // @[Switch.scala 30:36:@18753.4]
  wire  _T_40053; // @[Switch.scala 30:53:@18755.4]
  wire  valid_58_23; // @[Switch.scala 30:36:@18756.4]
  wire  _T_40056; // @[Switch.scala 30:53:@18758.4]
  wire  valid_58_24; // @[Switch.scala 30:36:@18759.4]
  wire  _T_40059; // @[Switch.scala 30:53:@18761.4]
  wire  valid_58_25; // @[Switch.scala 30:36:@18762.4]
  wire  _T_40062; // @[Switch.scala 30:53:@18764.4]
  wire  valid_58_26; // @[Switch.scala 30:36:@18765.4]
  wire  _T_40065; // @[Switch.scala 30:53:@18767.4]
  wire  valid_58_27; // @[Switch.scala 30:36:@18768.4]
  wire  _T_40068; // @[Switch.scala 30:53:@18770.4]
  wire  valid_58_28; // @[Switch.scala 30:36:@18771.4]
  wire  _T_40071; // @[Switch.scala 30:53:@18773.4]
  wire  valid_58_29; // @[Switch.scala 30:36:@18774.4]
  wire  _T_40074; // @[Switch.scala 30:53:@18776.4]
  wire  valid_58_30; // @[Switch.scala 30:36:@18777.4]
  wire  _T_40077; // @[Switch.scala 30:53:@18779.4]
  wire  valid_58_31; // @[Switch.scala 30:36:@18780.4]
  wire  _T_40080; // @[Switch.scala 30:53:@18782.4]
  wire  valid_58_32; // @[Switch.scala 30:36:@18783.4]
  wire  _T_40083; // @[Switch.scala 30:53:@18785.4]
  wire  valid_58_33; // @[Switch.scala 30:36:@18786.4]
  wire  _T_40086; // @[Switch.scala 30:53:@18788.4]
  wire  valid_58_34; // @[Switch.scala 30:36:@18789.4]
  wire  _T_40089; // @[Switch.scala 30:53:@18791.4]
  wire  valid_58_35; // @[Switch.scala 30:36:@18792.4]
  wire  _T_40092; // @[Switch.scala 30:53:@18794.4]
  wire  valid_58_36; // @[Switch.scala 30:36:@18795.4]
  wire  _T_40095; // @[Switch.scala 30:53:@18797.4]
  wire  valid_58_37; // @[Switch.scala 30:36:@18798.4]
  wire  _T_40098; // @[Switch.scala 30:53:@18800.4]
  wire  valid_58_38; // @[Switch.scala 30:36:@18801.4]
  wire  _T_40101; // @[Switch.scala 30:53:@18803.4]
  wire  valid_58_39; // @[Switch.scala 30:36:@18804.4]
  wire  _T_40104; // @[Switch.scala 30:53:@18806.4]
  wire  valid_58_40; // @[Switch.scala 30:36:@18807.4]
  wire  _T_40107; // @[Switch.scala 30:53:@18809.4]
  wire  valid_58_41; // @[Switch.scala 30:36:@18810.4]
  wire  _T_40110; // @[Switch.scala 30:53:@18812.4]
  wire  valid_58_42; // @[Switch.scala 30:36:@18813.4]
  wire  _T_40113; // @[Switch.scala 30:53:@18815.4]
  wire  valid_58_43; // @[Switch.scala 30:36:@18816.4]
  wire  _T_40116; // @[Switch.scala 30:53:@18818.4]
  wire  valid_58_44; // @[Switch.scala 30:36:@18819.4]
  wire  _T_40119; // @[Switch.scala 30:53:@18821.4]
  wire  valid_58_45; // @[Switch.scala 30:36:@18822.4]
  wire  _T_40122; // @[Switch.scala 30:53:@18824.4]
  wire  valid_58_46; // @[Switch.scala 30:36:@18825.4]
  wire  _T_40125; // @[Switch.scala 30:53:@18827.4]
  wire  valid_58_47; // @[Switch.scala 30:36:@18828.4]
  wire  _T_40128; // @[Switch.scala 30:53:@18830.4]
  wire  valid_58_48; // @[Switch.scala 30:36:@18831.4]
  wire  _T_40131; // @[Switch.scala 30:53:@18833.4]
  wire  valid_58_49; // @[Switch.scala 30:36:@18834.4]
  wire  _T_40134; // @[Switch.scala 30:53:@18836.4]
  wire  valid_58_50; // @[Switch.scala 30:36:@18837.4]
  wire  _T_40137; // @[Switch.scala 30:53:@18839.4]
  wire  valid_58_51; // @[Switch.scala 30:36:@18840.4]
  wire  _T_40140; // @[Switch.scala 30:53:@18842.4]
  wire  valid_58_52; // @[Switch.scala 30:36:@18843.4]
  wire  _T_40143; // @[Switch.scala 30:53:@18845.4]
  wire  valid_58_53; // @[Switch.scala 30:36:@18846.4]
  wire  _T_40146; // @[Switch.scala 30:53:@18848.4]
  wire  valid_58_54; // @[Switch.scala 30:36:@18849.4]
  wire  _T_40149; // @[Switch.scala 30:53:@18851.4]
  wire  valid_58_55; // @[Switch.scala 30:36:@18852.4]
  wire  _T_40152; // @[Switch.scala 30:53:@18854.4]
  wire  valid_58_56; // @[Switch.scala 30:36:@18855.4]
  wire  _T_40155; // @[Switch.scala 30:53:@18857.4]
  wire  valid_58_57; // @[Switch.scala 30:36:@18858.4]
  wire  _T_40158; // @[Switch.scala 30:53:@18860.4]
  wire  valid_58_58; // @[Switch.scala 30:36:@18861.4]
  wire  _T_40161; // @[Switch.scala 30:53:@18863.4]
  wire  valid_58_59; // @[Switch.scala 30:36:@18864.4]
  wire  _T_40164; // @[Switch.scala 30:53:@18866.4]
  wire  valid_58_60; // @[Switch.scala 30:36:@18867.4]
  wire  _T_40167; // @[Switch.scala 30:53:@18869.4]
  wire  valid_58_61; // @[Switch.scala 30:36:@18870.4]
  wire  _T_40170; // @[Switch.scala 30:53:@18872.4]
  wire  valid_58_62; // @[Switch.scala 30:36:@18873.4]
  wire  _T_40173; // @[Switch.scala 30:53:@18875.4]
  wire  valid_58_63; // @[Switch.scala 30:36:@18876.4]
  wire [5:0] _T_40239; // @[Mux.scala 31:69:@18878.4]
  wire [5:0] _T_40240; // @[Mux.scala 31:69:@18879.4]
  wire [5:0] _T_40241; // @[Mux.scala 31:69:@18880.4]
  wire [5:0] _T_40242; // @[Mux.scala 31:69:@18881.4]
  wire [5:0] _T_40243; // @[Mux.scala 31:69:@18882.4]
  wire [5:0] _T_40244; // @[Mux.scala 31:69:@18883.4]
  wire [5:0] _T_40245; // @[Mux.scala 31:69:@18884.4]
  wire [5:0] _T_40246; // @[Mux.scala 31:69:@18885.4]
  wire [5:0] _T_40247; // @[Mux.scala 31:69:@18886.4]
  wire [5:0] _T_40248; // @[Mux.scala 31:69:@18887.4]
  wire [5:0] _T_40249; // @[Mux.scala 31:69:@18888.4]
  wire [5:0] _T_40250; // @[Mux.scala 31:69:@18889.4]
  wire [5:0] _T_40251; // @[Mux.scala 31:69:@18890.4]
  wire [5:0] _T_40252; // @[Mux.scala 31:69:@18891.4]
  wire [5:0] _T_40253; // @[Mux.scala 31:69:@18892.4]
  wire [5:0] _T_40254; // @[Mux.scala 31:69:@18893.4]
  wire [5:0] _T_40255; // @[Mux.scala 31:69:@18894.4]
  wire [5:0] _T_40256; // @[Mux.scala 31:69:@18895.4]
  wire [5:0] _T_40257; // @[Mux.scala 31:69:@18896.4]
  wire [5:0] _T_40258; // @[Mux.scala 31:69:@18897.4]
  wire [5:0] _T_40259; // @[Mux.scala 31:69:@18898.4]
  wire [5:0] _T_40260; // @[Mux.scala 31:69:@18899.4]
  wire [5:0] _T_40261; // @[Mux.scala 31:69:@18900.4]
  wire [5:0] _T_40262; // @[Mux.scala 31:69:@18901.4]
  wire [5:0] _T_40263; // @[Mux.scala 31:69:@18902.4]
  wire [5:0] _T_40264; // @[Mux.scala 31:69:@18903.4]
  wire [5:0] _T_40265; // @[Mux.scala 31:69:@18904.4]
  wire [5:0] _T_40266; // @[Mux.scala 31:69:@18905.4]
  wire [5:0] _T_40267; // @[Mux.scala 31:69:@18906.4]
  wire [5:0] _T_40268; // @[Mux.scala 31:69:@18907.4]
  wire [5:0] _T_40269; // @[Mux.scala 31:69:@18908.4]
  wire [5:0] _T_40270; // @[Mux.scala 31:69:@18909.4]
  wire [5:0] _T_40271; // @[Mux.scala 31:69:@18910.4]
  wire [5:0] _T_40272; // @[Mux.scala 31:69:@18911.4]
  wire [5:0] _T_40273; // @[Mux.scala 31:69:@18912.4]
  wire [5:0] _T_40274; // @[Mux.scala 31:69:@18913.4]
  wire [5:0] _T_40275; // @[Mux.scala 31:69:@18914.4]
  wire [5:0] _T_40276; // @[Mux.scala 31:69:@18915.4]
  wire [5:0] _T_40277; // @[Mux.scala 31:69:@18916.4]
  wire [5:0] _T_40278; // @[Mux.scala 31:69:@18917.4]
  wire [5:0] _T_40279; // @[Mux.scala 31:69:@18918.4]
  wire [5:0] _T_40280; // @[Mux.scala 31:69:@18919.4]
  wire [5:0] _T_40281; // @[Mux.scala 31:69:@18920.4]
  wire [5:0] _T_40282; // @[Mux.scala 31:69:@18921.4]
  wire [5:0] _T_40283; // @[Mux.scala 31:69:@18922.4]
  wire [5:0] _T_40284; // @[Mux.scala 31:69:@18923.4]
  wire [5:0] _T_40285; // @[Mux.scala 31:69:@18924.4]
  wire [5:0] _T_40286; // @[Mux.scala 31:69:@18925.4]
  wire [5:0] _T_40287; // @[Mux.scala 31:69:@18926.4]
  wire [5:0] _T_40288; // @[Mux.scala 31:69:@18927.4]
  wire [5:0] _T_40289; // @[Mux.scala 31:69:@18928.4]
  wire [5:0] _T_40290; // @[Mux.scala 31:69:@18929.4]
  wire [5:0] _T_40291; // @[Mux.scala 31:69:@18930.4]
  wire [5:0] _T_40292; // @[Mux.scala 31:69:@18931.4]
  wire [5:0] _T_40293; // @[Mux.scala 31:69:@18932.4]
  wire [5:0] _T_40294; // @[Mux.scala 31:69:@18933.4]
  wire [5:0] _T_40295; // @[Mux.scala 31:69:@18934.4]
  wire [5:0] _T_40296; // @[Mux.scala 31:69:@18935.4]
  wire [5:0] _T_40297; // @[Mux.scala 31:69:@18936.4]
  wire [5:0] _T_40298; // @[Mux.scala 31:69:@18937.4]
  wire [5:0] _T_40299; // @[Mux.scala 31:69:@18938.4]
  wire [5:0] _T_40300; // @[Mux.scala 31:69:@18939.4]
  wire [5:0] select_58; // @[Mux.scala 31:69:@18940.4]
  wire [47:0] _GEN_3713; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3714; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3715; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3716; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3717; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3718; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3719; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3720; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3721; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3722; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3723; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3724; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3725; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3726; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3727; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3728; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3729; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3730; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3731; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3732; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3733; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3734; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3735; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3736; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3737; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3738; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3739; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3740; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3741; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3742; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3743; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3744; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3745; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3746; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3747; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3748; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3749; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3750; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3751; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3752; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3753; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3754; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3755; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3756; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3757; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3758; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3759; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3760; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3761; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3762; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3763; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3764; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3765; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3766; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3767; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3768; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3769; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3770; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3771; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3772; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3773; // @[Switch.scala 33:19:@18942.4]
  wire [47:0] _GEN_3774; // @[Switch.scala 33:19:@18942.4]
  wire [7:0] _T_40309; // @[Switch.scala 34:32:@18949.4]
  wire [15:0] _T_40317; // @[Switch.scala 34:32:@18957.4]
  wire [7:0] _T_40324; // @[Switch.scala 34:32:@18964.4]
  wire [31:0] _T_40333; // @[Switch.scala 34:32:@18973.4]
  wire [7:0] _T_40340; // @[Switch.scala 34:32:@18980.4]
  wire [15:0] _T_40348; // @[Switch.scala 34:32:@18988.4]
  wire [7:0] _T_40355; // @[Switch.scala 34:32:@18995.4]
  wire [31:0] _T_40364; // @[Switch.scala 34:32:@19004.4]
  wire [63:0] _T_40365; // @[Switch.scala 34:32:@19005.4]
  wire  _T_40369; // @[Switch.scala 30:53:@19008.4]
  wire  valid_59_0; // @[Switch.scala 30:36:@19009.4]
  wire  _T_40372; // @[Switch.scala 30:53:@19011.4]
  wire  valid_59_1; // @[Switch.scala 30:36:@19012.4]
  wire  _T_40375; // @[Switch.scala 30:53:@19014.4]
  wire  valid_59_2; // @[Switch.scala 30:36:@19015.4]
  wire  _T_40378; // @[Switch.scala 30:53:@19017.4]
  wire  valid_59_3; // @[Switch.scala 30:36:@19018.4]
  wire  _T_40381; // @[Switch.scala 30:53:@19020.4]
  wire  valid_59_4; // @[Switch.scala 30:36:@19021.4]
  wire  _T_40384; // @[Switch.scala 30:53:@19023.4]
  wire  valid_59_5; // @[Switch.scala 30:36:@19024.4]
  wire  _T_40387; // @[Switch.scala 30:53:@19026.4]
  wire  valid_59_6; // @[Switch.scala 30:36:@19027.4]
  wire  _T_40390; // @[Switch.scala 30:53:@19029.4]
  wire  valid_59_7; // @[Switch.scala 30:36:@19030.4]
  wire  _T_40393; // @[Switch.scala 30:53:@19032.4]
  wire  valid_59_8; // @[Switch.scala 30:36:@19033.4]
  wire  _T_40396; // @[Switch.scala 30:53:@19035.4]
  wire  valid_59_9; // @[Switch.scala 30:36:@19036.4]
  wire  _T_40399; // @[Switch.scala 30:53:@19038.4]
  wire  valid_59_10; // @[Switch.scala 30:36:@19039.4]
  wire  _T_40402; // @[Switch.scala 30:53:@19041.4]
  wire  valid_59_11; // @[Switch.scala 30:36:@19042.4]
  wire  _T_40405; // @[Switch.scala 30:53:@19044.4]
  wire  valid_59_12; // @[Switch.scala 30:36:@19045.4]
  wire  _T_40408; // @[Switch.scala 30:53:@19047.4]
  wire  valid_59_13; // @[Switch.scala 30:36:@19048.4]
  wire  _T_40411; // @[Switch.scala 30:53:@19050.4]
  wire  valid_59_14; // @[Switch.scala 30:36:@19051.4]
  wire  _T_40414; // @[Switch.scala 30:53:@19053.4]
  wire  valid_59_15; // @[Switch.scala 30:36:@19054.4]
  wire  _T_40417; // @[Switch.scala 30:53:@19056.4]
  wire  valid_59_16; // @[Switch.scala 30:36:@19057.4]
  wire  _T_40420; // @[Switch.scala 30:53:@19059.4]
  wire  valid_59_17; // @[Switch.scala 30:36:@19060.4]
  wire  _T_40423; // @[Switch.scala 30:53:@19062.4]
  wire  valid_59_18; // @[Switch.scala 30:36:@19063.4]
  wire  _T_40426; // @[Switch.scala 30:53:@19065.4]
  wire  valid_59_19; // @[Switch.scala 30:36:@19066.4]
  wire  _T_40429; // @[Switch.scala 30:53:@19068.4]
  wire  valid_59_20; // @[Switch.scala 30:36:@19069.4]
  wire  _T_40432; // @[Switch.scala 30:53:@19071.4]
  wire  valid_59_21; // @[Switch.scala 30:36:@19072.4]
  wire  _T_40435; // @[Switch.scala 30:53:@19074.4]
  wire  valid_59_22; // @[Switch.scala 30:36:@19075.4]
  wire  _T_40438; // @[Switch.scala 30:53:@19077.4]
  wire  valid_59_23; // @[Switch.scala 30:36:@19078.4]
  wire  _T_40441; // @[Switch.scala 30:53:@19080.4]
  wire  valid_59_24; // @[Switch.scala 30:36:@19081.4]
  wire  _T_40444; // @[Switch.scala 30:53:@19083.4]
  wire  valid_59_25; // @[Switch.scala 30:36:@19084.4]
  wire  _T_40447; // @[Switch.scala 30:53:@19086.4]
  wire  valid_59_26; // @[Switch.scala 30:36:@19087.4]
  wire  _T_40450; // @[Switch.scala 30:53:@19089.4]
  wire  valid_59_27; // @[Switch.scala 30:36:@19090.4]
  wire  _T_40453; // @[Switch.scala 30:53:@19092.4]
  wire  valid_59_28; // @[Switch.scala 30:36:@19093.4]
  wire  _T_40456; // @[Switch.scala 30:53:@19095.4]
  wire  valid_59_29; // @[Switch.scala 30:36:@19096.4]
  wire  _T_40459; // @[Switch.scala 30:53:@19098.4]
  wire  valid_59_30; // @[Switch.scala 30:36:@19099.4]
  wire  _T_40462; // @[Switch.scala 30:53:@19101.4]
  wire  valid_59_31; // @[Switch.scala 30:36:@19102.4]
  wire  _T_40465; // @[Switch.scala 30:53:@19104.4]
  wire  valid_59_32; // @[Switch.scala 30:36:@19105.4]
  wire  _T_40468; // @[Switch.scala 30:53:@19107.4]
  wire  valid_59_33; // @[Switch.scala 30:36:@19108.4]
  wire  _T_40471; // @[Switch.scala 30:53:@19110.4]
  wire  valid_59_34; // @[Switch.scala 30:36:@19111.4]
  wire  _T_40474; // @[Switch.scala 30:53:@19113.4]
  wire  valid_59_35; // @[Switch.scala 30:36:@19114.4]
  wire  _T_40477; // @[Switch.scala 30:53:@19116.4]
  wire  valid_59_36; // @[Switch.scala 30:36:@19117.4]
  wire  _T_40480; // @[Switch.scala 30:53:@19119.4]
  wire  valid_59_37; // @[Switch.scala 30:36:@19120.4]
  wire  _T_40483; // @[Switch.scala 30:53:@19122.4]
  wire  valid_59_38; // @[Switch.scala 30:36:@19123.4]
  wire  _T_40486; // @[Switch.scala 30:53:@19125.4]
  wire  valid_59_39; // @[Switch.scala 30:36:@19126.4]
  wire  _T_40489; // @[Switch.scala 30:53:@19128.4]
  wire  valid_59_40; // @[Switch.scala 30:36:@19129.4]
  wire  _T_40492; // @[Switch.scala 30:53:@19131.4]
  wire  valid_59_41; // @[Switch.scala 30:36:@19132.4]
  wire  _T_40495; // @[Switch.scala 30:53:@19134.4]
  wire  valid_59_42; // @[Switch.scala 30:36:@19135.4]
  wire  _T_40498; // @[Switch.scala 30:53:@19137.4]
  wire  valid_59_43; // @[Switch.scala 30:36:@19138.4]
  wire  _T_40501; // @[Switch.scala 30:53:@19140.4]
  wire  valid_59_44; // @[Switch.scala 30:36:@19141.4]
  wire  _T_40504; // @[Switch.scala 30:53:@19143.4]
  wire  valid_59_45; // @[Switch.scala 30:36:@19144.4]
  wire  _T_40507; // @[Switch.scala 30:53:@19146.4]
  wire  valid_59_46; // @[Switch.scala 30:36:@19147.4]
  wire  _T_40510; // @[Switch.scala 30:53:@19149.4]
  wire  valid_59_47; // @[Switch.scala 30:36:@19150.4]
  wire  _T_40513; // @[Switch.scala 30:53:@19152.4]
  wire  valid_59_48; // @[Switch.scala 30:36:@19153.4]
  wire  _T_40516; // @[Switch.scala 30:53:@19155.4]
  wire  valid_59_49; // @[Switch.scala 30:36:@19156.4]
  wire  _T_40519; // @[Switch.scala 30:53:@19158.4]
  wire  valid_59_50; // @[Switch.scala 30:36:@19159.4]
  wire  _T_40522; // @[Switch.scala 30:53:@19161.4]
  wire  valid_59_51; // @[Switch.scala 30:36:@19162.4]
  wire  _T_40525; // @[Switch.scala 30:53:@19164.4]
  wire  valid_59_52; // @[Switch.scala 30:36:@19165.4]
  wire  _T_40528; // @[Switch.scala 30:53:@19167.4]
  wire  valid_59_53; // @[Switch.scala 30:36:@19168.4]
  wire  _T_40531; // @[Switch.scala 30:53:@19170.4]
  wire  valid_59_54; // @[Switch.scala 30:36:@19171.4]
  wire  _T_40534; // @[Switch.scala 30:53:@19173.4]
  wire  valid_59_55; // @[Switch.scala 30:36:@19174.4]
  wire  _T_40537; // @[Switch.scala 30:53:@19176.4]
  wire  valid_59_56; // @[Switch.scala 30:36:@19177.4]
  wire  _T_40540; // @[Switch.scala 30:53:@19179.4]
  wire  valid_59_57; // @[Switch.scala 30:36:@19180.4]
  wire  _T_40543; // @[Switch.scala 30:53:@19182.4]
  wire  valid_59_58; // @[Switch.scala 30:36:@19183.4]
  wire  _T_40546; // @[Switch.scala 30:53:@19185.4]
  wire  valid_59_59; // @[Switch.scala 30:36:@19186.4]
  wire  _T_40549; // @[Switch.scala 30:53:@19188.4]
  wire  valid_59_60; // @[Switch.scala 30:36:@19189.4]
  wire  _T_40552; // @[Switch.scala 30:53:@19191.4]
  wire  valid_59_61; // @[Switch.scala 30:36:@19192.4]
  wire  _T_40555; // @[Switch.scala 30:53:@19194.4]
  wire  valid_59_62; // @[Switch.scala 30:36:@19195.4]
  wire  _T_40558; // @[Switch.scala 30:53:@19197.4]
  wire  valid_59_63; // @[Switch.scala 30:36:@19198.4]
  wire [5:0] _T_40624; // @[Mux.scala 31:69:@19200.4]
  wire [5:0] _T_40625; // @[Mux.scala 31:69:@19201.4]
  wire [5:0] _T_40626; // @[Mux.scala 31:69:@19202.4]
  wire [5:0] _T_40627; // @[Mux.scala 31:69:@19203.4]
  wire [5:0] _T_40628; // @[Mux.scala 31:69:@19204.4]
  wire [5:0] _T_40629; // @[Mux.scala 31:69:@19205.4]
  wire [5:0] _T_40630; // @[Mux.scala 31:69:@19206.4]
  wire [5:0] _T_40631; // @[Mux.scala 31:69:@19207.4]
  wire [5:0] _T_40632; // @[Mux.scala 31:69:@19208.4]
  wire [5:0] _T_40633; // @[Mux.scala 31:69:@19209.4]
  wire [5:0] _T_40634; // @[Mux.scala 31:69:@19210.4]
  wire [5:0] _T_40635; // @[Mux.scala 31:69:@19211.4]
  wire [5:0] _T_40636; // @[Mux.scala 31:69:@19212.4]
  wire [5:0] _T_40637; // @[Mux.scala 31:69:@19213.4]
  wire [5:0] _T_40638; // @[Mux.scala 31:69:@19214.4]
  wire [5:0] _T_40639; // @[Mux.scala 31:69:@19215.4]
  wire [5:0] _T_40640; // @[Mux.scala 31:69:@19216.4]
  wire [5:0] _T_40641; // @[Mux.scala 31:69:@19217.4]
  wire [5:0] _T_40642; // @[Mux.scala 31:69:@19218.4]
  wire [5:0] _T_40643; // @[Mux.scala 31:69:@19219.4]
  wire [5:0] _T_40644; // @[Mux.scala 31:69:@19220.4]
  wire [5:0] _T_40645; // @[Mux.scala 31:69:@19221.4]
  wire [5:0] _T_40646; // @[Mux.scala 31:69:@19222.4]
  wire [5:0] _T_40647; // @[Mux.scala 31:69:@19223.4]
  wire [5:0] _T_40648; // @[Mux.scala 31:69:@19224.4]
  wire [5:0] _T_40649; // @[Mux.scala 31:69:@19225.4]
  wire [5:0] _T_40650; // @[Mux.scala 31:69:@19226.4]
  wire [5:0] _T_40651; // @[Mux.scala 31:69:@19227.4]
  wire [5:0] _T_40652; // @[Mux.scala 31:69:@19228.4]
  wire [5:0] _T_40653; // @[Mux.scala 31:69:@19229.4]
  wire [5:0] _T_40654; // @[Mux.scala 31:69:@19230.4]
  wire [5:0] _T_40655; // @[Mux.scala 31:69:@19231.4]
  wire [5:0] _T_40656; // @[Mux.scala 31:69:@19232.4]
  wire [5:0] _T_40657; // @[Mux.scala 31:69:@19233.4]
  wire [5:0] _T_40658; // @[Mux.scala 31:69:@19234.4]
  wire [5:0] _T_40659; // @[Mux.scala 31:69:@19235.4]
  wire [5:0] _T_40660; // @[Mux.scala 31:69:@19236.4]
  wire [5:0] _T_40661; // @[Mux.scala 31:69:@19237.4]
  wire [5:0] _T_40662; // @[Mux.scala 31:69:@19238.4]
  wire [5:0] _T_40663; // @[Mux.scala 31:69:@19239.4]
  wire [5:0] _T_40664; // @[Mux.scala 31:69:@19240.4]
  wire [5:0] _T_40665; // @[Mux.scala 31:69:@19241.4]
  wire [5:0] _T_40666; // @[Mux.scala 31:69:@19242.4]
  wire [5:0] _T_40667; // @[Mux.scala 31:69:@19243.4]
  wire [5:0] _T_40668; // @[Mux.scala 31:69:@19244.4]
  wire [5:0] _T_40669; // @[Mux.scala 31:69:@19245.4]
  wire [5:0] _T_40670; // @[Mux.scala 31:69:@19246.4]
  wire [5:0] _T_40671; // @[Mux.scala 31:69:@19247.4]
  wire [5:0] _T_40672; // @[Mux.scala 31:69:@19248.4]
  wire [5:0] _T_40673; // @[Mux.scala 31:69:@19249.4]
  wire [5:0] _T_40674; // @[Mux.scala 31:69:@19250.4]
  wire [5:0] _T_40675; // @[Mux.scala 31:69:@19251.4]
  wire [5:0] _T_40676; // @[Mux.scala 31:69:@19252.4]
  wire [5:0] _T_40677; // @[Mux.scala 31:69:@19253.4]
  wire [5:0] _T_40678; // @[Mux.scala 31:69:@19254.4]
  wire [5:0] _T_40679; // @[Mux.scala 31:69:@19255.4]
  wire [5:0] _T_40680; // @[Mux.scala 31:69:@19256.4]
  wire [5:0] _T_40681; // @[Mux.scala 31:69:@19257.4]
  wire [5:0] _T_40682; // @[Mux.scala 31:69:@19258.4]
  wire [5:0] _T_40683; // @[Mux.scala 31:69:@19259.4]
  wire [5:0] _T_40684; // @[Mux.scala 31:69:@19260.4]
  wire [5:0] _T_40685; // @[Mux.scala 31:69:@19261.4]
  wire [5:0] select_59; // @[Mux.scala 31:69:@19262.4]
  wire [47:0] _GEN_3777; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3778; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3779; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3780; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3781; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3782; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3783; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3784; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3785; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3786; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3787; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3788; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3789; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3790; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3791; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3792; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3793; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3794; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3795; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3796; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3797; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3798; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3799; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3800; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3801; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3802; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3803; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3804; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3805; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3806; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3807; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3808; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3809; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3810; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3811; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3812; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3813; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3814; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3815; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3816; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3817; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3818; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3819; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3820; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3821; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3822; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3823; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3824; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3825; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3826; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3827; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3828; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3829; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3830; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3831; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3832; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3833; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3834; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3835; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3836; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3837; // @[Switch.scala 33:19:@19264.4]
  wire [47:0] _GEN_3838; // @[Switch.scala 33:19:@19264.4]
  wire [7:0] _T_40694; // @[Switch.scala 34:32:@19271.4]
  wire [15:0] _T_40702; // @[Switch.scala 34:32:@19279.4]
  wire [7:0] _T_40709; // @[Switch.scala 34:32:@19286.4]
  wire [31:0] _T_40718; // @[Switch.scala 34:32:@19295.4]
  wire [7:0] _T_40725; // @[Switch.scala 34:32:@19302.4]
  wire [15:0] _T_40733; // @[Switch.scala 34:32:@19310.4]
  wire [7:0] _T_40740; // @[Switch.scala 34:32:@19317.4]
  wire [31:0] _T_40749; // @[Switch.scala 34:32:@19326.4]
  wire [63:0] _T_40750; // @[Switch.scala 34:32:@19327.4]
  wire  _T_40754; // @[Switch.scala 30:53:@19330.4]
  wire  valid_60_0; // @[Switch.scala 30:36:@19331.4]
  wire  _T_40757; // @[Switch.scala 30:53:@19333.4]
  wire  valid_60_1; // @[Switch.scala 30:36:@19334.4]
  wire  _T_40760; // @[Switch.scala 30:53:@19336.4]
  wire  valid_60_2; // @[Switch.scala 30:36:@19337.4]
  wire  _T_40763; // @[Switch.scala 30:53:@19339.4]
  wire  valid_60_3; // @[Switch.scala 30:36:@19340.4]
  wire  _T_40766; // @[Switch.scala 30:53:@19342.4]
  wire  valid_60_4; // @[Switch.scala 30:36:@19343.4]
  wire  _T_40769; // @[Switch.scala 30:53:@19345.4]
  wire  valid_60_5; // @[Switch.scala 30:36:@19346.4]
  wire  _T_40772; // @[Switch.scala 30:53:@19348.4]
  wire  valid_60_6; // @[Switch.scala 30:36:@19349.4]
  wire  _T_40775; // @[Switch.scala 30:53:@19351.4]
  wire  valid_60_7; // @[Switch.scala 30:36:@19352.4]
  wire  _T_40778; // @[Switch.scala 30:53:@19354.4]
  wire  valid_60_8; // @[Switch.scala 30:36:@19355.4]
  wire  _T_40781; // @[Switch.scala 30:53:@19357.4]
  wire  valid_60_9; // @[Switch.scala 30:36:@19358.4]
  wire  _T_40784; // @[Switch.scala 30:53:@19360.4]
  wire  valid_60_10; // @[Switch.scala 30:36:@19361.4]
  wire  _T_40787; // @[Switch.scala 30:53:@19363.4]
  wire  valid_60_11; // @[Switch.scala 30:36:@19364.4]
  wire  _T_40790; // @[Switch.scala 30:53:@19366.4]
  wire  valid_60_12; // @[Switch.scala 30:36:@19367.4]
  wire  _T_40793; // @[Switch.scala 30:53:@19369.4]
  wire  valid_60_13; // @[Switch.scala 30:36:@19370.4]
  wire  _T_40796; // @[Switch.scala 30:53:@19372.4]
  wire  valid_60_14; // @[Switch.scala 30:36:@19373.4]
  wire  _T_40799; // @[Switch.scala 30:53:@19375.4]
  wire  valid_60_15; // @[Switch.scala 30:36:@19376.4]
  wire  _T_40802; // @[Switch.scala 30:53:@19378.4]
  wire  valid_60_16; // @[Switch.scala 30:36:@19379.4]
  wire  _T_40805; // @[Switch.scala 30:53:@19381.4]
  wire  valid_60_17; // @[Switch.scala 30:36:@19382.4]
  wire  _T_40808; // @[Switch.scala 30:53:@19384.4]
  wire  valid_60_18; // @[Switch.scala 30:36:@19385.4]
  wire  _T_40811; // @[Switch.scala 30:53:@19387.4]
  wire  valid_60_19; // @[Switch.scala 30:36:@19388.4]
  wire  _T_40814; // @[Switch.scala 30:53:@19390.4]
  wire  valid_60_20; // @[Switch.scala 30:36:@19391.4]
  wire  _T_40817; // @[Switch.scala 30:53:@19393.4]
  wire  valid_60_21; // @[Switch.scala 30:36:@19394.4]
  wire  _T_40820; // @[Switch.scala 30:53:@19396.4]
  wire  valid_60_22; // @[Switch.scala 30:36:@19397.4]
  wire  _T_40823; // @[Switch.scala 30:53:@19399.4]
  wire  valid_60_23; // @[Switch.scala 30:36:@19400.4]
  wire  _T_40826; // @[Switch.scala 30:53:@19402.4]
  wire  valid_60_24; // @[Switch.scala 30:36:@19403.4]
  wire  _T_40829; // @[Switch.scala 30:53:@19405.4]
  wire  valid_60_25; // @[Switch.scala 30:36:@19406.4]
  wire  _T_40832; // @[Switch.scala 30:53:@19408.4]
  wire  valid_60_26; // @[Switch.scala 30:36:@19409.4]
  wire  _T_40835; // @[Switch.scala 30:53:@19411.4]
  wire  valid_60_27; // @[Switch.scala 30:36:@19412.4]
  wire  _T_40838; // @[Switch.scala 30:53:@19414.4]
  wire  valid_60_28; // @[Switch.scala 30:36:@19415.4]
  wire  _T_40841; // @[Switch.scala 30:53:@19417.4]
  wire  valid_60_29; // @[Switch.scala 30:36:@19418.4]
  wire  _T_40844; // @[Switch.scala 30:53:@19420.4]
  wire  valid_60_30; // @[Switch.scala 30:36:@19421.4]
  wire  _T_40847; // @[Switch.scala 30:53:@19423.4]
  wire  valid_60_31; // @[Switch.scala 30:36:@19424.4]
  wire  _T_40850; // @[Switch.scala 30:53:@19426.4]
  wire  valid_60_32; // @[Switch.scala 30:36:@19427.4]
  wire  _T_40853; // @[Switch.scala 30:53:@19429.4]
  wire  valid_60_33; // @[Switch.scala 30:36:@19430.4]
  wire  _T_40856; // @[Switch.scala 30:53:@19432.4]
  wire  valid_60_34; // @[Switch.scala 30:36:@19433.4]
  wire  _T_40859; // @[Switch.scala 30:53:@19435.4]
  wire  valid_60_35; // @[Switch.scala 30:36:@19436.4]
  wire  _T_40862; // @[Switch.scala 30:53:@19438.4]
  wire  valid_60_36; // @[Switch.scala 30:36:@19439.4]
  wire  _T_40865; // @[Switch.scala 30:53:@19441.4]
  wire  valid_60_37; // @[Switch.scala 30:36:@19442.4]
  wire  _T_40868; // @[Switch.scala 30:53:@19444.4]
  wire  valid_60_38; // @[Switch.scala 30:36:@19445.4]
  wire  _T_40871; // @[Switch.scala 30:53:@19447.4]
  wire  valid_60_39; // @[Switch.scala 30:36:@19448.4]
  wire  _T_40874; // @[Switch.scala 30:53:@19450.4]
  wire  valid_60_40; // @[Switch.scala 30:36:@19451.4]
  wire  _T_40877; // @[Switch.scala 30:53:@19453.4]
  wire  valid_60_41; // @[Switch.scala 30:36:@19454.4]
  wire  _T_40880; // @[Switch.scala 30:53:@19456.4]
  wire  valid_60_42; // @[Switch.scala 30:36:@19457.4]
  wire  _T_40883; // @[Switch.scala 30:53:@19459.4]
  wire  valid_60_43; // @[Switch.scala 30:36:@19460.4]
  wire  _T_40886; // @[Switch.scala 30:53:@19462.4]
  wire  valid_60_44; // @[Switch.scala 30:36:@19463.4]
  wire  _T_40889; // @[Switch.scala 30:53:@19465.4]
  wire  valid_60_45; // @[Switch.scala 30:36:@19466.4]
  wire  _T_40892; // @[Switch.scala 30:53:@19468.4]
  wire  valid_60_46; // @[Switch.scala 30:36:@19469.4]
  wire  _T_40895; // @[Switch.scala 30:53:@19471.4]
  wire  valid_60_47; // @[Switch.scala 30:36:@19472.4]
  wire  _T_40898; // @[Switch.scala 30:53:@19474.4]
  wire  valid_60_48; // @[Switch.scala 30:36:@19475.4]
  wire  _T_40901; // @[Switch.scala 30:53:@19477.4]
  wire  valid_60_49; // @[Switch.scala 30:36:@19478.4]
  wire  _T_40904; // @[Switch.scala 30:53:@19480.4]
  wire  valid_60_50; // @[Switch.scala 30:36:@19481.4]
  wire  _T_40907; // @[Switch.scala 30:53:@19483.4]
  wire  valid_60_51; // @[Switch.scala 30:36:@19484.4]
  wire  _T_40910; // @[Switch.scala 30:53:@19486.4]
  wire  valid_60_52; // @[Switch.scala 30:36:@19487.4]
  wire  _T_40913; // @[Switch.scala 30:53:@19489.4]
  wire  valid_60_53; // @[Switch.scala 30:36:@19490.4]
  wire  _T_40916; // @[Switch.scala 30:53:@19492.4]
  wire  valid_60_54; // @[Switch.scala 30:36:@19493.4]
  wire  _T_40919; // @[Switch.scala 30:53:@19495.4]
  wire  valid_60_55; // @[Switch.scala 30:36:@19496.4]
  wire  _T_40922; // @[Switch.scala 30:53:@19498.4]
  wire  valid_60_56; // @[Switch.scala 30:36:@19499.4]
  wire  _T_40925; // @[Switch.scala 30:53:@19501.4]
  wire  valid_60_57; // @[Switch.scala 30:36:@19502.4]
  wire  _T_40928; // @[Switch.scala 30:53:@19504.4]
  wire  valid_60_58; // @[Switch.scala 30:36:@19505.4]
  wire  _T_40931; // @[Switch.scala 30:53:@19507.4]
  wire  valid_60_59; // @[Switch.scala 30:36:@19508.4]
  wire  _T_40934; // @[Switch.scala 30:53:@19510.4]
  wire  valid_60_60; // @[Switch.scala 30:36:@19511.4]
  wire  _T_40937; // @[Switch.scala 30:53:@19513.4]
  wire  valid_60_61; // @[Switch.scala 30:36:@19514.4]
  wire  _T_40940; // @[Switch.scala 30:53:@19516.4]
  wire  valid_60_62; // @[Switch.scala 30:36:@19517.4]
  wire  _T_40943; // @[Switch.scala 30:53:@19519.4]
  wire  valid_60_63; // @[Switch.scala 30:36:@19520.4]
  wire [5:0] _T_41009; // @[Mux.scala 31:69:@19522.4]
  wire [5:0] _T_41010; // @[Mux.scala 31:69:@19523.4]
  wire [5:0] _T_41011; // @[Mux.scala 31:69:@19524.4]
  wire [5:0] _T_41012; // @[Mux.scala 31:69:@19525.4]
  wire [5:0] _T_41013; // @[Mux.scala 31:69:@19526.4]
  wire [5:0] _T_41014; // @[Mux.scala 31:69:@19527.4]
  wire [5:0] _T_41015; // @[Mux.scala 31:69:@19528.4]
  wire [5:0] _T_41016; // @[Mux.scala 31:69:@19529.4]
  wire [5:0] _T_41017; // @[Mux.scala 31:69:@19530.4]
  wire [5:0] _T_41018; // @[Mux.scala 31:69:@19531.4]
  wire [5:0] _T_41019; // @[Mux.scala 31:69:@19532.4]
  wire [5:0] _T_41020; // @[Mux.scala 31:69:@19533.4]
  wire [5:0] _T_41021; // @[Mux.scala 31:69:@19534.4]
  wire [5:0] _T_41022; // @[Mux.scala 31:69:@19535.4]
  wire [5:0] _T_41023; // @[Mux.scala 31:69:@19536.4]
  wire [5:0] _T_41024; // @[Mux.scala 31:69:@19537.4]
  wire [5:0] _T_41025; // @[Mux.scala 31:69:@19538.4]
  wire [5:0] _T_41026; // @[Mux.scala 31:69:@19539.4]
  wire [5:0] _T_41027; // @[Mux.scala 31:69:@19540.4]
  wire [5:0] _T_41028; // @[Mux.scala 31:69:@19541.4]
  wire [5:0] _T_41029; // @[Mux.scala 31:69:@19542.4]
  wire [5:0] _T_41030; // @[Mux.scala 31:69:@19543.4]
  wire [5:0] _T_41031; // @[Mux.scala 31:69:@19544.4]
  wire [5:0] _T_41032; // @[Mux.scala 31:69:@19545.4]
  wire [5:0] _T_41033; // @[Mux.scala 31:69:@19546.4]
  wire [5:0] _T_41034; // @[Mux.scala 31:69:@19547.4]
  wire [5:0] _T_41035; // @[Mux.scala 31:69:@19548.4]
  wire [5:0] _T_41036; // @[Mux.scala 31:69:@19549.4]
  wire [5:0] _T_41037; // @[Mux.scala 31:69:@19550.4]
  wire [5:0] _T_41038; // @[Mux.scala 31:69:@19551.4]
  wire [5:0] _T_41039; // @[Mux.scala 31:69:@19552.4]
  wire [5:0] _T_41040; // @[Mux.scala 31:69:@19553.4]
  wire [5:0] _T_41041; // @[Mux.scala 31:69:@19554.4]
  wire [5:0] _T_41042; // @[Mux.scala 31:69:@19555.4]
  wire [5:0] _T_41043; // @[Mux.scala 31:69:@19556.4]
  wire [5:0] _T_41044; // @[Mux.scala 31:69:@19557.4]
  wire [5:0] _T_41045; // @[Mux.scala 31:69:@19558.4]
  wire [5:0] _T_41046; // @[Mux.scala 31:69:@19559.4]
  wire [5:0] _T_41047; // @[Mux.scala 31:69:@19560.4]
  wire [5:0] _T_41048; // @[Mux.scala 31:69:@19561.4]
  wire [5:0] _T_41049; // @[Mux.scala 31:69:@19562.4]
  wire [5:0] _T_41050; // @[Mux.scala 31:69:@19563.4]
  wire [5:0] _T_41051; // @[Mux.scala 31:69:@19564.4]
  wire [5:0] _T_41052; // @[Mux.scala 31:69:@19565.4]
  wire [5:0] _T_41053; // @[Mux.scala 31:69:@19566.4]
  wire [5:0] _T_41054; // @[Mux.scala 31:69:@19567.4]
  wire [5:0] _T_41055; // @[Mux.scala 31:69:@19568.4]
  wire [5:0] _T_41056; // @[Mux.scala 31:69:@19569.4]
  wire [5:0] _T_41057; // @[Mux.scala 31:69:@19570.4]
  wire [5:0] _T_41058; // @[Mux.scala 31:69:@19571.4]
  wire [5:0] _T_41059; // @[Mux.scala 31:69:@19572.4]
  wire [5:0] _T_41060; // @[Mux.scala 31:69:@19573.4]
  wire [5:0] _T_41061; // @[Mux.scala 31:69:@19574.4]
  wire [5:0] _T_41062; // @[Mux.scala 31:69:@19575.4]
  wire [5:0] _T_41063; // @[Mux.scala 31:69:@19576.4]
  wire [5:0] _T_41064; // @[Mux.scala 31:69:@19577.4]
  wire [5:0] _T_41065; // @[Mux.scala 31:69:@19578.4]
  wire [5:0] _T_41066; // @[Mux.scala 31:69:@19579.4]
  wire [5:0] _T_41067; // @[Mux.scala 31:69:@19580.4]
  wire [5:0] _T_41068; // @[Mux.scala 31:69:@19581.4]
  wire [5:0] _T_41069; // @[Mux.scala 31:69:@19582.4]
  wire [5:0] _T_41070; // @[Mux.scala 31:69:@19583.4]
  wire [5:0] select_60; // @[Mux.scala 31:69:@19584.4]
  wire [47:0] _GEN_3841; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3842; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3843; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3844; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3845; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3846; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3847; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3848; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3849; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3850; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3851; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3852; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3853; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3854; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3855; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3856; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3857; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3858; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3859; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3860; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3861; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3862; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3863; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3864; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3865; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3866; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3867; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3868; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3869; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3870; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3871; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3872; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3873; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3874; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3875; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3876; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3877; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3878; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3879; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3880; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3881; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3882; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3883; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3884; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3885; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3886; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3887; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3888; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3889; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3890; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3891; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3892; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3893; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3894; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3895; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3896; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3897; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3898; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3899; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3900; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3901; // @[Switch.scala 33:19:@19586.4]
  wire [47:0] _GEN_3902; // @[Switch.scala 33:19:@19586.4]
  wire [7:0] _T_41079; // @[Switch.scala 34:32:@19593.4]
  wire [15:0] _T_41087; // @[Switch.scala 34:32:@19601.4]
  wire [7:0] _T_41094; // @[Switch.scala 34:32:@19608.4]
  wire [31:0] _T_41103; // @[Switch.scala 34:32:@19617.4]
  wire [7:0] _T_41110; // @[Switch.scala 34:32:@19624.4]
  wire [15:0] _T_41118; // @[Switch.scala 34:32:@19632.4]
  wire [7:0] _T_41125; // @[Switch.scala 34:32:@19639.4]
  wire [31:0] _T_41134; // @[Switch.scala 34:32:@19648.4]
  wire [63:0] _T_41135; // @[Switch.scala 34:32:@19649.4]
  wire  _T_41139; // @[Switch.scala 30:53:@19652.4]
  wire  valid_61_0; // @[Switch.scala 30:36:@19653.4]
  wire  _T_41142; // @[Switch.scala 30:53:@19655.4]
  wire  valid_61_1; // @[Switch.scala 30:36:@19656.4]
  wire  _T_41145; // @[Switch.scala 30:53:@19658.4]
  wire  valid_61_2; // @[Switch.scala 30:36:@19659.4]
  wire  _T_41148; // @[Switch.scala 30:53:@19661.4]
  wire  valid_61_3; // @[Switch.scala 30:36:@19662.4]
  wire  _T_41151; // @[Switch.scala 30:53:@19664.4]
  wire  valid_61_4; // @[Switch.scala 30:36:@19665.4]
  wire  _T_41154; // @[Switch.scala 30:53:@19667.4]
  wire  valid_61_5; // @[Switch.scala 30:36:@19668.4]
  wire  _T_41157; // @[Switch.scala 30:53:@19670.4]
  wire  valid_61_6; // @[Switch.scala 30:36:@19671.4]
  wire  _T_41160; // @[Switch.scala 30:53:@19673.4]
  wire  valid_61_7; // @[Switch.scala 30:36:@19674.4]
  wire  _T_41163; // @[Switch.scala 30:53:@19676.4]
  wire  valid_61_8; // @[Switch.scala 30:36:@19677.4]
  wire  _T_41166; // @[Switch.scala 30:53:@19679.4]
  wire  valid_61_9; // @[Switch.scala 30:36:@19680.4]
  wire  _T_41169; // @[Switch.scala 30:53:@19682.4]
  wire  valid_61_10; // @[Switch.scala 30:36:@19683.4]
  wire  _T_41172; // @[Switch.scala 30:53:@19685.4]
  wire  valid_61_11; // @[Switch.scala 30:36:@19686.4]
  wire  _T_41175; // @[Switch.scala 30:53:@19688.4]
  wire  valid_61_12; // @[Switch.scala 30:36:@19689.4]
  wire  _T_41178; // @[Switch.scala 30:53:@19691.4]
  wire  valid_61_13; // @[Switch.scala 30:36:@19692.4]
  wire  _T_41181; // @[Switch.scala 30:53:@19694.4]
  wire  valid_61_14; // @[Switch.scala 30:36:@19695.4]
  wire  _T_41184; // @[Switch.scala 30:53:@19697.4]
  wire  valid_61_15; // @[Switch.scala 30:36:@19698.4]
  wire  _T_41187; // @[Switch.scala 30:53:@19700.4]
  wire  valid_61_16; // @[Switch.scala 30:36:@19701.4]
  wire  _T_41190; // @[Switch.scala 30:53:@19703.4]
  wire  valid_61_17; // @[Switch.scala 30:36:@19704.4]
  wire  _T_41193; // @[Switch.scala 30:53:@19706.4]
  wire  valid_61_18; // @[Switch.scala 30:36:@19707.4]
  wire  _T_41196; // @[Switch.scala 30:53:@19709.4]
  wire  valid_61_19; // @[Switch.scala 30:36:@19710.4]
  wire  _T_41199; // @[Switch.scala 30:53:@19712.4]
  wire  valid_61_20; // @[Switch.scala 30:36:@19713.4]
  wire  _T_41202; // @[Switch.scala 30:53:@19715.4]
  wire  valid_61_21; // @[Switch.scala 30:36:@19716.4]
  wire  _T_41205; // @[Switch.scala 30:53:@19718.4]
  wire  valid_61_22; // @[Switch.scala 30:36:@19719.4]
  wire  _T_41208; // @[Switch.scala 30:53:@19721.4]
  wire  valid_61_23; // @[Switch.scala 30:36:@19722.4]
  wire  _T_41211; // @[Switch.scala 30:53:@19724.4]
  wire  valid_61_24; // @[Switch.scala 30:36:@19725.4]
  wire  _T_41214; // @[Switch.scala 30:53:@19727.4]
  wire  valid_61_25; // @[Switch.scala 30:36:@19728.4]
  wire  _T_41217; // @[Switch.scala 30:53:@19730.4]
  wire  valid_61_26; // @[Switch.scala 30:36:@19731.4]
  wire  _T_41220; // @[Switch.scala 30:53:@19733.4]
  wire  valid_61_27; // @[Switch.scala 30:36:@19734.4]
  wire  _T_41223; // @[Switch.scala 30:53:@19736.4]
  wire  valid_61_28; // @[Switch.scala 30:36:@19737.4]
  wire  _T_41226; // @[Switch.scala 30:53:@19739.4]
  wire  valid_61_29; // @[Switch.scala 30:36:@19740.4]
  wire  _T_41229; // @[Switch.scala 30:53:@19742.4]
  wire  valid_61_30; // @[Switch.scala 30:36:@19743.4]
  wire  _T_41232; // @[Switch.scala 30:53:@19745.4]
  wire  valid_61_31; // @[Switch.scala 30:36:@19746.4]
  wire  _T_41235; // @[Switch.scala 30:53:@19748.4]
  wire  valid_61_32; // @[Switch.scala 30:36:@19749.4]
  wire  _T_41238; // @[Switch.scala 30:53:@19751.4]
  wire  valid_61_33; // @[Switch.scala 30:36:@19752.4]
  wire  _T_41241; // @[Switch.scala 30:53:@19754.4]
  wire  valid_61_34; // @[Switch.scala 30:36:@19755.4]
  wire  _T_41244; // @[Switch.scala 30:53:@19757.4]
  wire  valid_61_35; // @[Switch.scala 30:36:@19758.4]
  wire  _T_41247; // @[Switch.scala 30:53:@19760.4]
  wire  valid_61_36; // @[Switch.scala 30:36:@19761.4]
  wire  _T_41250; // @[Switch.scala 30:53:@19763.4]
  wire  valid_61_37; // @[Switch.scala 30:36:@19764.4]
  wire  _T_41253; // @[Switch.scala 30:53:@19766.4]
  wire  valid_61_38; // @[Switch.scala 30:36:@19767.4]
  wire  _T_41256; // @[Switch.scala 30:53:@19769.4]
  wire  valid_61_39; // @[Switch.scala 30:36:@19770.4]
  wire  _T_41259; // @[Switch.scala 30:53:@19772.4]
  wire  valid_61_40; // @[Switch.scala 30:36:@19773.4]
  wire  _T_41262; // @[Switch.scala 30:53:@19775.4]
  wire  valid_61_41; // @[Switch.scala 30:36:@19776.4]
  wire  _T_41265; // @[Switch.scala 30:53:@19778.4]
  wire  valid_61_42; // @[Switch.scala 30:36:@19779.4]
  wire  _T_41268; // @[Switch.scala 30:53:@19781.4]
  wire  valid_61_43; // @[Switch.scala 30:36:@19782.4]
  wire  _T_41271; // @[Switch.scala 30:53:@19784.4]
  wire  valid_61_44; // @[Switch.scala 30:36:@19785.4]
  wire  _T_41274; // @[Switch.scala 30:53:@19787.4]
  wire  valid_61_45; // @[Switch.scala 30:36:@19788.4]
  wire  _T_41277; // @[Switch.scala 30:53:@19790.4]
  wire  valid_61_46; // @[Switch.scala 30:36:@19791.4]
  wire  _T_41280; // @[Switch.scala 30:53:@19793.4]
  wire  valid_61_47; // @[Switch.scala 30:36:@19794.4]
  wire  _T_41283; // @[Switch.scala 30:53:@19796.4]
  wire  valid_61_48; // @[Switch.scala 30:36:@19797.4]
  wire  _T_41286; // @[Switch.scala 30:53:@19799.4]
  wire  valid_61_49; // @[Switch.scala 30:36:@19800.4]
  wire  _T_41289; // @[Switch.scala 30:53:@19802.4]
  wire  valid_61_50; // @[Switch.scala 30:36:@19803.4]
  wire  _T_41292; // @[Switch.scala 30:53:@19805.4]
  wire  valid_61_51; // @[Switch.scala 30:36:@19806.4]
  wire  _T_41295; // @[Switch.scala 30:53:@19808.4]
  wire  valid_61_52; // @[Switch.scala 30:36:@19809.4]
  wire  _T_41298; // @[Switch.scala 30:53:@19811.4]
  wire  valid_61_53; // @[Switch.scala 30:36:@19812.4]
  wire  _T_41301; // @[Switch.scala 30:53:@19814.4]
  wire  valid_61_54; // @[Switch.scala 30:36:@19815.4]
  wire  _T_41304; // @[Switch.scala 30:53:@19817.4]
  wire  valid_61_55; // @[Switch.scala 30:36:@19818.4]
  wire  _T_41307; // @[Switch.scala 30:53:@19820.4]
  wire  valid_61_56; // @[Switch.scala 30:36:@19821.4]
  wire  _T_41310; // @[Switch.scala 30:53:@19823.4]
  wire  valid_61_57; // @[Switch.scala 30:36:@19824.4]
  wire  _T_41313; // @[Switch.scala 30:53:@19826.4]
  wire  valid_61_58; // @[Switch.scala 30:36:@19827.4]
  wire  _T_41316; // @[Switch.scala 30:53:@19829.4]
  wire  valid_61_59; // @[Switch.scala 30:36:@19830.4]
  wire  _T_41319; // @[Switch.scala 30:53:@19832.4]
  wire  valid_61_60; // @[Switch.scala 30:36:@19833.4]
  wire  _T_41322; // @[Switch.scala 30:53:@19835.4]
  wire  valid_61_61; // @[Switch.scala 30:36:@19836.4]
  wire  _T_41325; // @[Switch.scala 30:53:@19838.4]
  wire  valid_61_62; // @[Switch.scala 30:36:@19839.4]
  wire  _T_41328; // @[Switch.scala 30:53:@19841.4]
  wire  valid_61_63; // @[Switch.scala 30:36:@19842.4]
  wire [5:0] _T_41394; // @[Mux.scala 31:69:@19844.4]
  wire [5:0] _T_41395; // @[Mux.scala 31:69:@19845.4]
  wire [5:0] _T_41396; // @[Mux.scala 31:69:@19846.4]
  wire [5:0] _T_41397; // @[Mux.scala 31:69:@19847.4]
  wire [5:0] _T_41398; // @[Mux.scala 31:69:@19848.4]
  wire [5:0] _T_41399; // @[Mux.scala 31:69:@19849.4]
  wire [5:0] _T_41400; // @[Mux.scala 31:69:@19850.4]
  wire [5:0] _T_41401; // @[Mux.scala 31:69:@19851.4]
  wire [5:0] _T_41402; // @[Mux.scala 31:69:@19852.4]
  wire [5:0] _T_41403; // @[Mux.scala 31:69:@19853.4]
  wire [5:0] _T_41404; // @[Mux.scala 31:69:@19854.4]
  wire [5:0] _T_41405; // @[Mux.scala 31:69:@19855.4]
  wire [5:0] _T_41406; // @[Mux.scala 31:69:@19856.4]
  wire [5:0] _T_41407; // @[Mux.scala 31:69:@19857.4]
  wire [5:0] _T_41408; // @[Mux.scala 31:69:@19858.4]
  wire [5:0] _T_41409; // @[Mux.scala 31:69:@19859.4]
  wire [5:0] _T_41410; // @[Mux.scala 31:69:@19860.4]
  wire [5:0] _T_41411; // @[Mux.scala 31:69:@19861.4]
  wire [5:0] _T_41412; // @[Mux.scala 31:69:@19862.4]
  wire [5:0] _T_41413; // @[Mux.scala 31:69:@19863.4]
  wire [5:0] _T_41414; // @[Mux.scala 31:69:@19864.4]
  wire [5:0] _T_41415; // @[Mux.scala 31:69:@19865.4]
  wire [5:0] _T_41416; // @[Mux.scala 31:69:@19866.4]
  wire [5:0] _T_41417; // @[Mux.scala 31:69:@19867.4]
  wire [5:0] _T_41418; // @[Mux.scala 31:69:@19868.4]
  wire [5:0] _T_41419; // @[Mux.scala 31:69:@19869.4]
  wire [5:0] _T_41420; // @[Mux.scala 31:69:@19870.4]
  wire [5:0] _T_41421; // @[Mux.scala 31:69:@19871.4]
  wire [5:0] _T_41422; // @[Mux.scala 31:69:@19872.4]
  wire [5:0] _T_41423; // @[Mux.scala 31:69:@19873.4]
  wire [5:0] _T_41424; // @[Mux.scala 31:69:@19874.4]
  wire [5:0] _T_41425; // @[Mux.scala 31:69:@19875.4]
  wire [5:0] _T_41426; // @[Mux.scala 31:69:@19876.4]
  wire [5:0] _T_41427; // @[Mux.scala 31:69:@19877.4]
  wire [5:0] _T_41428; // @[Mux.scala 31:69:@19878.4]
  wire [5:0] _T_41429; // @[Mux.scala 31:69:@19879.4]
  wire [5:0] _T_41430; // @[Mux.scala 31:69:@19880.4]
  wire [5:0] _T_41431; // @[Mux.scala 31:69:@19881.4]
  wire [5:0] _T_41432; // @[Mux.scala 31:69:@19882.4]
  wire [5:0] _T_41433; // @[Mux.scala 31:69:@19883.4]
  wire [5:0] _T_41434; // @[Mux.scala 31:69:@19884.4]
  wire [5:0] _T_41435; // @[Mux.scala 31:69:@19885.4]
  wire [5:0] _T_41436; // @[Mux.scala 31:69:@19886.4]
  wire [5:0] _T_41437; // @[Mux.scala 31:69:@19887.4]
  wire [5:0] _T_41438; // @[Mux.scala 31:69:@19888.4]
  wire [5:0] _T_41439; // @[Mux.scala 31:69:@19889.4]
  wire [5:0] _T_41440; // @[Mux.scala 31:69:@19890.4]
  wire [5:0] _T_41441; // @[Mux.scala 31:69:@19891.4]
  wire [5:0] _T_41442; // @[Mux.scala 31:69:@19892.4]
  wire [5:0] _T_41443; // @[Mux.scala 31:69:@19893.4]
  wire [5:0] _T_41444; // @[Mux.scala 31:69:@19894.4]
  wire [5:0] _T_41445; // @[Mux.scala 31:69:@19895.4]
  wire [5:0] _T_41446; // @[Mux.scala 31:69:@19896.4]
  wire [5:0] _T_41447; // @[Mux.scala 31:69:@19897.4]
  wire [5:0] _T_41448; // @[Mux.scala 31:69:@19898.4]
  wire [5:0] _T_41449; // @[Mux.scala 31:69:@19899.4]
  wire [5:0] _T_41450; // @[Mux.scala 31:69:@19900.4]
  wire [5:0] _T_41451; // @[Mux.scala 31:69:@19901.4]
  wire [5:0] _T_41452; // @[Mux.scala 31:69:@19902.4]
  wire [5:0] _T_41453; // @[Mux.scala 31:69:@19903.4]
  wire [5:0] _T_41454; // @[Mux.scala 31:69:@19904.4]
  wire [5:0] _T_41455; // @[Mux.scala 31:69:@19905.4]
  wire [5:0] select_61; // @[Mux.scala 31:69:@19906.4]
  wire [47:0] _GEN_3905; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3906; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3907; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3908; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3909; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3910; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3911; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3912; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3913; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3914; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3915; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3916; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3917; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3918; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3919; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3920; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3921; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3922; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3923; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3924; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3925; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3926; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3927; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3928; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3929; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3930; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3931; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3932; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3933; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3934; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3935; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3936; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3937; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3938; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3939; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3940; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3941; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3942; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3943; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3944; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3945; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3946; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3947; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3948; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3949; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3950; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3951; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3952; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3953; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3954; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3955; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3956; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3957; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3958; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3959; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3960; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3961; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3962; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3963; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3964; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3965; // @[Switch.scala 33:19:@19908.4]
  wire [47:0] _GEN_3966; // @[Switch.scala 33:19:@19908.4]
  wire [7:0] _T_41464; // @[Switch.scala 34:32:@19915.4]
  wire [15:0] _T_41472; // @[Switch.scala 34:32:@19923.4]
  wire [7:0] _T_41479; // @[Switch.scala 34:32:@19930.4]
  wire [31:0] _T_41488; // @[Switch.scala 34:32:@19939.4]
  wire [7:0] _T_41495; // @[Switch.scala 34:32:@19946.4]
  wire [15:0] _T_41503; // @[Switch.scala 34:32:@19954.4]
  wire [7:0] _T_41510; // @[Switch.scala 34:32:@19961.4]
  wire [31:0] _T_41519; // @[Switch.scala 34:32:@19970.4]
  wire [63:0] _T_41520; // @[Switch.scala 34:32:@19971.4]
  wire  _T_41524; // @[Switch.scala 30:53:@19974.4]
  wire  valid_62_0; // @[Switch.scala 30:36:@19975.4]
  wire  _T_41527; // @[Switch.scala 30:53:@19977.4]
  wire  valid_62_1; // @[Switch.scala 30:36:@19978.4]
  wire  _T_41530; // @[Switch.scala 30:53:@19980.4]
  wire  valid_62_2; // @[Switch.scala 30:36:@19981.4]
  wire  _T_41533; // @[Switch.scala 30:53:@19983.4]
  wire  valid_62_3; // @[Switch.scala 30:36:@19984.4]
  wire  _T_41536; // @[Switch.scala 30:53:@19986.4]
  wire  valid_62_4; // @[Switch.scala 30:36:@19987.4]
  wire  _T_41539; // @[Switch.scala 30:53:@19989.4]
  wire  valid_62_5; // @[Switch.scala 30:36:@19990.4]
  wire  _T_41542; // @[Switch.scala 30:53:@19992.4]
  wire  valid_62_6; // @[Switch.scala 30:36:@19993.4]
  wire  _T_41545; // @[Switch.scala 30:53:@19995.4]
  wire  valid_62_7; // @[Switch.scala 30:36:@19996.4]
  wire  _T_41548; // @[Switch.scala 30:53:@19998.4]
  wire  valid_62_8; // @[Switch.scala 30:36:@19999.4]
  wire  _T_41551; // @[Switch.scala 30:53:@20001.4]
  wire  valid_62_9; // @[Switch.scala 30:36:@20002.4]
  wire  _T_41554; // @[Switch.scala 30:53:@20004.4]
  wire  valid_62_10; // @[Switch.scala 30:36:@20005.4]
  wire  _T_41557; // @[Switch.scala 30:53:@20007.4]
  wire  valid_62_11; // @[Switch.scala 30:36:@20008.4]
  wire  _T_41560; // @[Switch.scala 30:53:@20010.4]
  wire  valid_62_12; // @[Switch.scala 30:36:@20011.4]
  wire  _T_41563; // @[Switch.scala 30:53:@20013.4]
  wire  valid_62_13; // @[Switch.scala 30:36:@20014.4]
  wire  _T_41566; // @[Switch.scala 30:53:@20016.4]
  wire  valid_62_14; // @[Switch.scala 30:36:@20017.4]
  wire  _T_41569; // @[Switch.scala 30:53:@20019.4]
  wire  valid_62_15; // @[Switch.scala 30:36:@20020.4]
  wire  _T_41572; // @[Switch.scala 30:53:@20022.4]
  wire  valid_62_16; // @[Switch.scala 30:36:@20023.4]
  wire  _T_41575; // @[Switch.scala 30:53:@20025.4]
  wire  valid_62_17; // @[Switch.scala 30:36:@20026.4]
  wire  _T_41578; // @[Switch.scala 30:53:@20028.4]
  wire  valid_62_18; // @[Switch.scala 30:36:@20029.4]
  wire  _T_41581; // @[Switch.scala 30:53:@20031.4]
  wire  valid_62_19; // @[Switch.scala 30:36:@20032.4]
  wire  _T_41584; // @[Switch.scala 30:53:@20034.4]
  wire  valid_62_20; // @[Switch.scala 30:36:@20035.4]
  wire  _T_41587; // @[Switch.scala 30:53:@20037.4]
  wire  valid_62_21; // @[Switch.scala 30:36:@20038.4]
  wire  _T_41590; // @[Switch.scala 30:53:@20040.4]
  wire  valid_62_22; // @[Switch.scala 30:36:@20041.4]
  wire  _T_41593; // @[Switch.scala 30:53:@20043.4]
  wire  valid_62_23; // @[Switch.scala 30:36:@20044.4]
  wire  _T_41596; // @[Switch.scala 30:53:@20046.4]
  wire  valid_62_24; // @[Switch.scala 30:36:@20047.4]
  wire  _T_41599; // @[Switch.scala 30:53:@20049.4]
  wire  valid_62_25; // @[Switch.scala 30:36:@20050.4]
  wire  _T_41602; // @[Switch.scala 30:53:@20052.4]
  wire  valid_62_26; // @[Switch.scala 30:36:@20053.4]
  wire  _T_41605; // @[Switch.scala 30:53:@20055.4]
  wire  valid_62_27; // @[Switch.scala 30:36:@20056.4]
  wire  _T_41608; // @[Switch.scala 30:53:@20058.4]
  wire  valid_62_28; // @[Switch.scala 30:36:@20059.4]
  wire  _T_41611; // @[Switch.scala 30:53:@20061.4]
  wire  valid_62_29; // @[Switch.scala 30:36:@20062.4]
  wire  _T_41614; // @[Switch.scala 30:53:@20064.4]
  wire  valid_62_30; // @[Switch.scala 30:36:@20065.4]
  wire  _T_41617; // @[Switch.scala 30:53:@20067.4]
  wire  valid_62_31; // @[Switch.scala 30:36:@20068.4]
  wire  _T_41620; // @[Switch.scala 30:53:@20070.4]
  wire  valid_62_32; // @[Switch.scala 30:36:@20071.4]
  wire  _T_41623; // @[Switch.scala 30:53:@20073.4]
  wire  valid_62_33; // @[Switch.scala 30:36:@20074.4]
  wire  _T_41626; // @[Switch.scala 30:53:@20076.4]
  wire  valid_62_34; // @[Switch.scala 30:36:@20077.4]
  wire  _T_41629; // @[Switch.scala 30:53:@20079.4]
  wire  valid_62_35; // @[Switch.scala 30:36:@20080.4]
  wire  _T_41632; // @[Switch.scala 30:53:@20082.4]
  wire  valid_62_36; // @[Switch.scala 30:36:@20083.4]
  wire  _T_41635; // @[Switch.scala 30:53:@20085.4]
  wire  valid_62_37; // @[Switch.scala 30:36:@20086.4]
  wire  _T_41638; // @[Switch.scala 30:53:@20088.4]
  wire  valid_62_38; // @[Switch.scala 30:36:@20089.4]
  wire  _T_41641; // @[Switch.scala 30:53:@20091.4]
  wire  valid_62_39; // @[Switch.scala 30:36:@20092.4]
  wire  _T_41644; // @[Switch.scala 30:53:@20094.4]
  wire  valid_62_40; // @[Switch.scala 30:36:@20095.4]
  wire  _T_41647; // @[Switch.scala 30:53:@20097.4]
  wire  valid_62_41; // @[Switch.scala 30:36:@20098.4]
  wire  _T_41650; // @[Switch.scala 30:53:@20100.4]
  wire  valid_62_42; // @[Switch.scala 30:36:@20101.4]
  wire  _T_41653; // @[Switch.scala 30:53:@20103.4]
  wire  valid_62_43; // @[Switch.scala 30:36:@20104.4]
  wire  _T_41656; // @[Switch.scala 30:53:@20106.4]
  wire  valid_62_44; // @[Switch.scala 30:36:@20107.4]
  wire  _T_41659; // @[Switch.scala 30:53:@20109.4]
  wire  valid_62_45; // @[Switch.scala 30:36:@20110.4]
  wire  _T_41662; // @[Switch.scala 30:53:@20112.4]
  wire  valid_62_46; // @[Switch.scala 30:36:@20113.4]
  wire  _T_41665; // @[Switch.scala 30:53:@20115.4]
  wire  valid_62_47; // @[Switch.scala 30:36:@20116.4]
  wire  _T_41668; // @[Switch.scala 30:53:@20118.4]
  wire  valid_62_48; // @[Switch.scala 30:36:@20119.4]
  wire  _T_41671; // @[Switch.scala 30:53:@20121.4]
  wire  valid_62_49; // @[Switch.scala 30:36:@20122.4]
  wire  _T_41674; // @[Switch.scala 30:53:@20124.4]
  wire  valid_62_50; // @[Switch.scala 30:36:@20125.4]
  wire  _T_41677; // @[Switch.scala 30:53:@20127.4]
  wire  valid_62_51; // @[Switch.scala 30:36:@20128.4]
  wire  _T_41680; // @[Switch.scala 30:53:@20130.4]
  wire  valid_62_52; // @[Switch.scala 30:36:@20131.4]
  wire  _T_41683; // @[Switch.scala 30:53:@20133.4]
  wire  valid_62_53; // @[Switch.scala 30:36:@20134.4]
  wire  _T_41686; // @[Switch.scala 30:53:@20136.4]
  wire  valid_62_54; // @[Switch.scala 30:36:@20137.4]
  wire  _T_41689; // @[Switch.scala 30:53:@20139.4]
  wire  valid_62_55; // @[Switch.scala 30:36:@20140.4]
  wire  _T_41692; // @[Switch.scala 30:53:@20142.4]
  wire  valid_62_56; // @[Switch.scala 30:36:@20143.4]
  wire  _T_41695; // @[Switch.scala 30:53:@20145.4]
  wire  valid_62_57; // @[Switch.scala 30:36:@20146.4]
  wire  _T_41698; // @[Switch.scala 30:53:@20148.4]
  wire  valid_62_58; // @[Switch.scala 30:36:@20149.4]
  wire  _T_41701; // @[Switch.scala 30:53:@20151.4]
  wire  valid_62_59; // @[Switch.scala 30:36:@20152.4]
  wire  _T_41704; // @[Switch.scala 30:53:@20154.4]
  wire  valid_62_60; // @[Switch.scala 30:36:@20155.4]
  wire  _T_41707; // @[Switch.scala 30:53:@20157.4]
  wire  valid_62_61; // @[Switch.scala 30:36:@20158.4]
  wire  _T_41710; // @[Switch.scala 30:53:@20160.4]
  wire  valid_62_62; // @[Switch.scala 30:36:@20161.4]
  wire  _T_41713; // @[Switch.scala 30:53:@20163.4]
  wire  valid_62_63; // @[Switch.scala 30:36:@20164.4]
  wire [5:0] _T_41779; // @[Mux.scala 31:69:@20166.4]
  wire [5:0] _T_41780; // @[Mux.scala 31:69:@20167.4]
  wire [5:0] _T_41781; // @[Mux.scala 31:69:@20168.4]
  wire [5:0] _T_41782; // @[Mux.scala 31:69:@20169.4]
  wire [5:0] _T_41783; // @[Mux.scala 31:69:@20170.4]
  wire [5:0] _T_41784; // @[Mux.scala 31:69:@20171.4]
  wire [5:0] _T_41785; // @[Mux.scala 31:69:@20172.4]
  wire [5:0] _T_41786; // @[Mux.scala 31:69:@20173.4]
  wire [5:0] _T_41787; // @[Mux.scala 31:69:@20174.4]
  wire [5:0] _T_41788; // @[Mux.scala 31:69:@20175.4]
  wire [5:0] _T_41789; // @[Mux.scala 31:69:@20176.4]
  wire [5:0] _T_41790; // @[Mux.scala 31:69:@20177.4]
  wire [5:0] _T_41791; // @[Mux.scala 31:69:@20178.4]
  wire [5:0] _T_41792; // @[Mux.scala 31:69:@20179.4]
  wire [5:0] _T_41793; // @[Mux.scala 31:69:@20180.4]
  wire [5:0] _T_41794; // @[Mux.scala 31:69:@20181.4]
  wire [5:0] _T_41795; // @[Mux.scala 31:69:@20182.4]
  wire [5:0] _T_41796; // @[Mux.scala 31:69:@20183.4]
  wire [5:0] _T_41797; // @[Mux.scala 31:69:@20184.4]
  wire [5:0] _T_41798; // @[Mux.scala 31:69:@20185.4]
  wire [5:0] _T_41799; // @[Mux.scala 31:69:@20186.4]
  wire [5:0] _T_41800; // @[Mux.scala 31:69:@20187.4]
  wire [5:0] _T_41801; // @[Mux.scala 31:69:@20188.4]
  wire [5:0] _T_41802; // @[Mux.scala 31:69:@20189.4]
  wire [5:0] _T_41803; // @[Mux.scala 31:69:@20190.4]
  wire [5:0] _T_41804; // @[Mux.scala 31:69:@20191.4]
  wire [5:0] _T_41805; // @[Mux.scala 31:69:@20192.4]
  wire [5:0] _T_41806; // @[Mux.scala 31:69:@20193.4]
  wire [5:0] _T_41807; // @[Mux.scala 31:69:@20194.4]
  wire [5:0] _T_41808; // @[Mux.scala 31:69:@20195.4]
  wire [5:0] _T_41809; // @[Mux.scala 31:69:@20196.4]
  wire [5:0] _T_41810; // @[Mux.scala 31:69:@20197.4]
  wire [5:0] _T_41811; // @[Mux.scala 31:69:@20198.4]
  wire [5:0] _T_41812; // @[Mux.scala 31:69:@20199.4]
  wire [5:0] _T_41813; // @[Mux.scala 31:69:@20200.4]
  wire [5:0] _T_41814; // @[Mux.scala 31:69:@20201.4]
  wire [5:0] _T_41815; // @[Mux.scala 31:69:@20202.4]
  wire [5:0] _T_41816; // @[Mux.scala 31:69:@20203.4]
  wire [5:0] _T_41817; // @[Mux.scala 31:69:@20204.4]
  wire [5:0] _T_41818; // @[Mux.scala 31:69:@20205.4]
  wire [5:0] _T_41819; // @[Mux.scala 31:69:@20206.4]
  wire [5:0] _T_41820; // @[Mux.scala 31:69:@20207.4]
  wire [5:0] _T_41821; // @[Mux.scala 31:69:@20208.4]
  wire [5:0] _T_41822; // @[Mux.scala 31:69:@20209.4]
  wire [5:0] _T_41823; // @[Mux.scala 31:69:@20210.4]
  wire [5:0] _T_41824; // @[Mux.scala 31:69:@20211.4]
  wire [5:0] _T_41825; // @[Mux.scala 31:69:@20212.4]
  wire [5:0] _T_41826; // @[Mux.scala 31:69:@20213.4]
  wire [5:0] _T_41827; // @[Mux.scala 31:69:@20214.4]
  wire [5:0] _T_41828; // @[Mux.scala 31:69:@20215.4]
  wire [5:0] _T_41829; // @[Mux.scala 31:69:@20216.4]
  wire [5:0] _T_41830; // @[Mux.scala 31:69:@20217.4]
  wire [5:0] _T_41831; // @[Mux.scala 31:69:@20218.4]
  wire [5:0] _T_41832; // @[Mux.scala 31:69:@20219.4]
  wire [5:0] _T_41833; // @[Mux.scala 31:69:@20220.4]
  wire [5:0] _T_41834; // @[Mux.scala 31:69:@20221.4]
  wire [5:0] _T_41835; // @[Mux.scala 31:69:@20222.4]
  wire [5:0] _T_41836; // @[Mux.scala 31:69:@20223.4]
  wire [5:0] _T_41837; // @[Mux.scala 31:69:@20224.4]
  wire [5:0] _T_41838; // @[Mux.scala 31:69:@20225.4]
  wire [5:0] _T_41839; // @[Mux.scala 31:69:@20226.4]
  wire [5:0] _T_41840; // @[Mux.scala 31:69:@20227.4]
  wire [5:0] select_62; // @[Mux.scala 31:69:@20228.4]
  wire [47:0] _GEN_3969; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_3970; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_3971; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_3972; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_3973; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_3974; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_3975; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_3976; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_3977; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_3978; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_3979; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_3980; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_3981; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_3982; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_3983; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_3984; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_3985; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_3986; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_3987; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_3988; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_3989; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_3990; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_3991; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_3992; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_3993; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_3994; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_3995; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_3996; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_3997; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_3998; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_3999; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_4000; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_4001; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_4002; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_4003; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_4004; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_4005; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_4006; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_4007; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_4008; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_4009; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_4010; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_4011; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_4012; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_4013; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_4014; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_4015; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_4016; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_4017; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_4018; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_4019; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_4020; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_4021; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_4022; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_4023; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_4024; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_4025; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_4026; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_4027; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_4028; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_4029; // @[Switch.scala 33:19:@20230.4]
  wire [47:0] _GEN_4030; // @[Switch.scala 33:19:@20230.4]
  wire [7:0] _T_41849; // @[Switch.scala 34:32:@20237.4]
  wire [15:0] _T_41857; // @[Switch.scala 34:32:@20245.4]
  wire [7:0] _T_41864; // @[Switch.scala 34:32:@20252.4]
  wire [31:0] _T_41873; // @[Switch.scala 34:32:@20261.4]
  wire [7:0] _T_41880; // @[Switch.scala 34:32:@20268.4]
  wire [15:0] _T_41888; // @[Switch.scala 34:32:@20276.4]
  wire [7:0] _T_41895; // @[Switch.scala 34:32:@20283.4]
  wire [31:0] _T_41904; // @[Switch.scala 34:32:@20292.4]
  wire [63:0] _T_41905; // @[Switch.scala 34:32:@20293.4]
  wire  _T_41909; // @[Switch.scala 30:53:@20296.4]
  wire  valid_63_0; // @[Switch.scala 30:36:@20297.4]
  wire  _T_41912; // @[Switch.scala 30:53:@20299.4]
  wire  valid_63_1; // @[Switch.scala 30:36:@20300.4]
  wire  _T_41915; // @[Switch.scala 30:53:@20302.4]
  wire  valid_63_2; // @[Switch.scala 30:36:@20303.4]
  wire  _T_41918; // @[Switch.scala 30:53:@20305.4]
  wire  valid_63_3; // @[Switch.scala 30:36:@20306.4]
  wire  _T_41921; // @[Switch.scala 30:53:@20308.4]
  wire  valid_63_4; // @[Switch.scala 30:36:@20309.4]
  wire  _T_41924; // @[Switch.scala 30:53:@20311.4]
  wire  valid_63_5; // @[Switch.scala 30:36:@20312.4]
  wire  _T_41927; // @[Switch.scala 30:53:@20314.4]
  wire  valid_63_6; // @[Switch.scala 30:36:@20315.4]
  wire  _T_41930; // @[Switch.scala 30:53:@20317.4]
  wire  valid_63_7; // @[Switch.scala 30:36:@20318.4]
  wire  _T_41933; // @[Switch.scala 30:53:@20320.4]
  wire  valid_63_8; // @[Switch.scala 30:36:@20321.4]
  wire  _T_41936; // @[Switch.scala 30:53:@20323.4]
  wire  valid_63_9; // @[Switch.scala 30:36:@20324.4]
  wire  _T_41939; // @[Switch.scala 30:53:@20326.4]
  wire  valid_63_10; // @[Switch.scala 30:36:@20327.4]
  wire  _T_41942; // @[Switch.scala 30:53:@20329.4]
  wire  valid_63_11; // @[Switch.scala 30:36:@20330.4]
  wire  _T_41945; // @[Switch.scala 30:53:@20332.4]
  wire  valid_63_12; // @[Switch.scala 30:36:@20333.4]
  wire  _T_41948; // @[Switch.scala 30:53:@20335.4]
  wire  valid_63_13; // @[Switch.scala 30:36:@20336.4]
  wire  _T_41951; // @[Switch.scala 30:53:@20338.4]
  wire  valid_63_14; // @[Switch.scala 30:36:@20339.4]
  wire  _T_41954; // @[Switch.scala 30:53:@20341.4]
  wire  valid_63_15; // @[Switch.scala 30:36:@20342.4]
  wire  _T_41957; // @[Switch.scala 30:53:@20344.4]
  wire  valid_63_16; // @[Switch.scala 30:36:@20345.4]
  wire  _T_41960; // @[Switch.scala 30:53:@20347.4]
  wire  valid_63_17; // @[Switch.scala 30:36:@20348.4]
  wire  _T_41963; // @[Switch.scala 30:53:@20350.4]
  wire  valid_63_18; // @[Switch.scala 30:36:@20351.4]
  wire  _T_41966; // @[Switch.scala 30:53:@20353.4]
  wire  valid_63_19; // @[Switch.scala 30:36:@20354.4]
  wire  _T_41969; // @[Switch.scala 30:53:@20356.4]
  wire  valid_63_20; // @[Switch.scala 30:36:@20357.4]
  wire  _T_41972; // @[Switch.scala 30:53:@20359.4]
  wire  valid_63_21; // @[Switch.scala 30:36:@20360.4]
  wire  _T_41975; // @[Switch.scala 30:53:@20362.4]
  wire  valid_63_22; // @[Switch.scala 30:36:@20363.4]
  wire  _T_41978; // @[Switch.scala 30:53:@20365.4]
  wire  valid_63_23; // @[Switch.scala 30:36:@20366.4]
  wire  _T_41981; // @[Switch.scala 30:53:@20368.4]
  wire  valid_63_24; // @[Switch.scala 30:36:@20369.4]
  wire  _T_41984; // @[Switch.scala 30:53:@20371.4]
  wire  valid_63_25; // @[Switch.scala 30:36:@20372.4]
  wire  _T_41987; // @[Switch.scala 30:53:@20374.4]
  wire  valid_63_26; // @[Switch.scala 30:36:@20375.4]
  wire  _T_41990; // @[Switch.scala 30:53:@20377.4]
  wire  valid_63_27; // @[Switch.scala 30:36:@20378.4]
  wire  _T_41993; // @[Switch.scala 30:53:@20380.4]
  wire  valid_63_28; // @[Switch.scala 30:36:@20381.4]
  wire  _T_41996; // @[Switch.scala 30:53:@20383.4]
  wire  valid_63_29; // @[Switch.scala 30:36:@20384.4]
  wire  _T_41999; // @[Switch.scala 30:53:@20386.4]
  wire  valid_63_30; // @[Switch.scala 30:36:@20387.4]
  wire  _T_42002; // @[Switch.scala 30:53:@20389.4]
  wire  valid_63_31; // @[Switch.scala 30:36:@20390.4]
  wire  _T_42005; // @[Switch.scala 30:53:@20392.4]
  wire  valid_63_32; // @[Switch.scala 30:36:@20393.4]
  wire  _T_42008; // @[Switch.scala 30:53:@20395.4]
  wire  valid_63_33; // @[Switch.scala 30:36:@20396.4]
  wire  _T_42011; // @[Switch.scala 30:53:@20398.4]
  wire  valid_63_34; // @[Switch.scala 30:36:@20399.4]
  wire  _T_42014; // @[Switch.scala 30:53:@20401.4]
  wire  valid_63_35; // @[Switch.scala 30:36:@20402.4]
  wire  _T_42017; // @[Switch.scala 30:53:@20404.4]
  wire  valid_63_36; // @[Switch.scala 30:36:@20405.4]
  wire  _T_42020; // @[Switch.scala 30:53:@20407.4]
  wire  valid_63_37; // @[Switch.scala 30:36:@20408.4]
  wire  _T_42023; // @[Switch.scala 30:53:@20410.4]
  wire  valid_63_38; // @[Switch.scala 30:36:@20411.4]
  wire  _T_42026; // @[Switch.scala 30:53:@20413.4]
  wire  valid_63_39; // @[Switch.scala 30:36:@20414.4]
  wire  _T_42029; // @[Switch.scala 30:53:@20416.4]
  wire  valid_63_40; // @[Switch.scala 30:36:@20417.4]
  wire  _T_42032; // @[Switch.scala 30:53:@20419.4]
  wire  valid_63_41; // @[Switch.scala 30:36:@20420.4]
  wire  _T_42035; // @[Switch.scala 30:53:@20422.4]
  wire  valid_63_42; // @[Switch.scala 30:36:@20423.4]
  wire  _T_42038; // @[Switch.scala 30:53:@20425.4]
  wire  valid_63_43; // @[Switch.scala 30:36:@20426.4]
  wire  _T_42041; // @[Switch.scala 30:53:@20428.4]
  wire  valid_63_44; // @[Switch.scala 30:36:@20429.4]
  wire  _T_42044; // @[Switch.scala 30:53:@20431.4]
  wire  valid_63_45; // @[Switch.scala 30:36:@20432.4]
  wire  _T_42047; // @[Switch.scala 30:53:@20434.4]
  wire  valid_63_46; // @[Switch.scala 30:36:@20435.4]
  wire  _T_42050; // @[Switch.scala 30:53:@20437.4]
  wire  valid_63_47; // @[Switch.scala 30:36:@20438.4]
  wire  _T_42053; // @[Switch.scala 30:53:@20440.4]
  wire  valid_63_48; // @[Switch.scala 30:36:@20441.4]
  wire  _T_42056; // @[Switch.scala 30:53:@20443.4]
  wire  valid_63_49; // @[Switch.scala 30:36:@20444.4]
  wire  _T_42059; // @[Switch.scala 30:53:@20446.4]
  wire  valid_63_50; // @[Switch.scala 30:36:@20447.4]
  wire  _T_42062; // @[Switch.scala 30:53:@20449.4]
  wire  valid_63_51; // @[Switch.scala 30:36:@20450.4]
  wire  _T_42065; // @[Switch.scala 30:53:@20452.4]
  wire  valid_63_52; // @[Switch.scala 30:36:@20453.4]
  wire  _T_42068; // @[Switch.scala 30:53:@20455.4]
  wire  valid_63_53; // @[Switch.scala 30:36:@20456.4]
  wire  _T_42071; // @[Switch.scala 30:53:@20458.4]
  wire  valid_63_54; // @[Switch.scala 30:36:@20459.4]
  wire  _T_42074; // @[Switch.scala 30:53:@20461.4]
  wire  valid_63_55; // @[Switch.scala 30:36:@20462.4]
  wire  _T_42077; // @[Switch.scala 30:53:@20464.4]
  wire  valid_63_56; // @[Switch.scala 30:36:@20465.4]
  wire  _T_42080; // @[Switch.scala 30:53:@20467.4]
  wire  valid_63_57; // @[Switch.scala 30:36:@20468.4]
  wire  _T_42083; // @[Switch.scala 30:53:@20470.4]
  wire  valid_63_58; // @[Switch.scala 30:36:@20471.4]
  wire  _T_42086; // @[Switch.scala 30:53:@20473.4]
  wire  valid_63_59; // @[Switch.scala 30:36:@20474.4]
  wire  _T_42089; // @[Switch.scala 30:53:@20476.4]
  wire  valid_63_60; // @[Switch.scala 30:36:@20477.4]
  wire  _T_42092; // @[Switch.scala 30:53:@20479.4]
  wire  valid_63_61; // @[Switch.scala 30:36:@20480.4]
  wire  _T_42095; // @[Switch.scala 30:53:@20482.4]
  wire  valid_63_62; // @[Switch.scala 30:36:@20483.4]
  wire  _T_42098; // @[Switch.scala 30:53:@20485.4]
  wire  valid_63_63; // @[Switch.scala 30:36:@20486.4]
  wire [5:0] _T_42164; // @[Mux.scala 31:69:@20488.4]
  wire [5:0] _T_42165; // @[Mux.scala 31:69:@20489.4]
  wire [5:0] _T_42166; // @[Mux.scala 31:69:@20490.4]
  wire [5:0] _T_42167; // @[Mux.scala 31:69:@20491.4]
  wire [5:0] _T_42168; // @[Mux.scala 31:69:@20492.4]
  wire [5:0] _T_42169; // @[Mux.scala 31:69:@20493.4]
  wire [5:0] _T_42170; // @[Mux.scala 31:69:@20494.4]
  wire [5:0] _T_42171; // @[Mux.scala 31:69:@20495.4]
  wire [5:0] _T_42172; // @[Mux.scala 31:69:@20496.4]
  wire [5:0] _T_42173; // @[Mux.scala 31:69:@20497.4]
  wire [5:0] _T_42174; // @[Mux.scala 31:69:@20498.4]
  wire [5:0] _T_42175; // @[Mux.scala 31:69:@20499.4]
  wire [5:0] _T_42176; // @[Mux.scala 31:69:@20500.4]
  wire [5:0] _T_42177; // @[Mux.scala 31:69:@20501.4]
  wire [5:0] _T_42178; // @[Mux.scala 31:69:@20502.4]
  wire [5:0] _T_42179; // @[Mux.scala 31:69:@20503.4]
  wire [5:0] _T_42180; // @[Mux.scala 31:69:@20504.4]
  wire [5:0] _T_42181; // @[Mux.scala 31:69:@20505.4]
  wire [5:0] _T_42182; // @[Mux.scala 31:69:@20506.4]
  wire [5:0] _T_42183; // @[Mux.scala 31:69:@20507.4]
  wire [5:0] _T_42184; // @[Mux.scala 31:69:@20508.4]
  wire [5:0] _T_42185; // @[Mux.scala 31:69:@20509.4]
  wire [5:0] _T_42186; // @[Mux.scala 31:69:@20510.4]
  wire [5:0] _T_42187; // @[Mux.scala 31:69:@20511.4]
  wire [5:0] _T_42188; // @[Mux.scala 31:69:@20512.4]
  wire [5:0] _T_42189; // @[Mux.scala 31:69:@20513.4]
  wire [5:0] _T_42190; // @[Mux.scala 31:69:@20514.4]
  wire [5:0] _T_42191; // @[Mux.scala 31:69:@20515.4]
  wire [5:0] _T_42192; // @[Mux.scala 31:69:@20516.4]
  wire [5:0] _T_42193; // @[Mux.scala 31:69:@20517.4]
  wire [5:0] _T_42194; // @[Mux.scala 31:69:@20518.4]
  wire [5:0] _T_42195; // @[Mux.scala 31:69:@20519.4]
  wire [5:0] _T_42196; // @[Mux.scala 31:69:@20520.4]
  wire [5:0] _T_42197; // @[Mux.scala 31:69:@20521.4]
  wire [5:0] _T_42198; // @[Mux.scala 31:69:@20522.4]
  wire [5:0] _T_42199; // @[Mux.scala 31:69:@20523.4]
  wire [5:0] _T_42200; // @[Mux.scala 31:69:@20524.4]
  wire [5:0] _T_42201; // @[Mux.scala 31:69:@20525.4]
  wire [5:0] _T_42202; // @[Mux.scala 31:69:@20526.4]
  wire [5:0] _T_42203; // @[Mux.scala 31:69:@20527.4]
  wire [5:0] _T_42204; // @[Mux.scala 31:69:@20528.4]
  wire [5:0] _T_42205; // @[Mux.scala 31:69:@20529.4]
  wire [5:0] _T_42206; // @[Mux.scala 31:69:@20530.4]
  wire [5:0] _T_42207; // @[Mux.scala 31:69:@20531.4]
  wire [5:0] _T_42208; // @[Mux.scala 31:69:@20532.4]
  wire [5:0] _T_42209; // @[Mux.scala 31:69:@20533.4]
  wire [5:0] _T_42210; // @[Mux.scala 31:69:@20534.4]
  wire [5:0] _T_42211; // @[Mux.scala 31:69:@20535.4]
  wire [5:0] _T_42212; // @[Mux.scala 31:69:@20536.4]
  wire [5:0] _T_42213; // @[Mux.scala 31:69:@20537.4]
  wire [5:0] _T_42214; // @[Mux.scala 31:69:@20538.4]
  wire [5:0] _T_42215; // @[Mux.scala 31:69:@20539.4]
  wire [5:0] _T_42216; // @[Mux.scala 31:69:@20540.4]
  wire [5:0] _T_42217; // @[Mux.scala 31:69:@20541.4]
  wire [5:0] _T_42218; // @[Mux.scala 31:69:@20542.4]
  wire [5:0] _T_42219; // @[Mux.scala 31:69:@20543.4]
  wire [5:0] _T_42220; // @[Mux.scala 31:69:@20544.4]
  wire [5:0] _T_42221; // @[Mux.scala 31:69:@20545.4]
  wire [5:0] _T_42222; // @[Mux.scala 31:69:@20546.4]
  wire [5:0] _T_42223; // @[Mux.scala 31:69:@20547.4]
  wire [5:0] _T_42224; // @[Mux.scala 31:69:@20548.4]
  wire [5:0] _T_42225; // @[Mux.scala 31:69:@20549.4]
  wire [5:0] select_63; // @[Mux.scala 31:69:@20550.4]
  wire [47:0] _GEN_4033; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4034; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4035; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4036; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4037; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4038; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4039; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4040; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4041; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4042; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4043; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4044; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4045; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4046; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4047; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4048; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4049; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4050; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4051; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4052; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4053; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4054; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4055; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4056; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4057; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4058; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4059; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4060; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4061; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4062; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4063; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4064; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4065; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4066; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4067; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4068; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4069; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4070; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4071; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4072; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4073; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4074; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4075; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4076; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4077; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4078; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4079; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4080; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4081; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4082; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4083; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4084; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4085; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4086; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4087; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4088; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4089; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4090; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4091; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4092; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4093; // @[Switch.scala 33:19:@20552.4]
  wire [47:0] _GEN_4094; // @[Switch.scala 33:19:@20552.4]
  wire [7:0] _T_42234; // @[Switch.scala 34:32:@20559.4]
  wire [15:0] _T_42242; // @[Switch.scala 34:32:@20567.4]
  wire [7:0] _T_42249; // @[Switch.scala 34:32:@20574.4]
  wire [31:0] _T_42258; // @[Switch.scala 34:32:@20583.4]
  wire [7:0] _T_42265; // @[Switch.scala 34:32:@20590.4]
  wire [15:0] _T_42273; // @[Switch.scala 34:32:@20598.4]
  wire [7:0] _T_42280; // @[Switch.scala 34:32:@20605.4]
  wire [31:0] _T_42289; // @[Switch.scala 34:32:@20614.4]
  wire [63:0] _T_42290; // @[Switch.scala 34:32:@20615.4]
  wire  _T_59460; // @[Switch.scala 41:52:@20619.4]
  wire  output_0_0; // @[Switch.scala 41:38:@20620.4]
  wire  _T_59463; // @[Switch.scala 41:52:@20622.4]
  wire  output_0_1; // @[Switch.scala 41:38:@20623.4]
  wire  _T_59466; // @[Switch.scala 41:52:@20625.4]
  wire  output_0_2; // @[Switch.scala 41:38:@20626.4]
  wire  _T_59469; // @[Switch.scala 41:52:@20628.4]
  wire  output_0_3; // @[Switch.scala 41:38:@20629.4]
  wire  _T_59472; // @[Switch.scala 41:52:@20631.4]
  wire  output_0_4; // @[Switch.scala 41:38:@20632.4]
  wire  _T_59475; // @[Switch.scala 41:52:@20634.4]
  wire  output_0_5; // @[Switch.scala 41:38:@20635.4]
  wire  _T_59478; // @[Switch.scala 41:52:@20637.4]
  wire  output_0_6; // @[Switch.scala 41:38:@20638.4]
  wire  _T_59481; // @[Switch.scala 41:52:@20640.4]
  wire  output_0_7; // @[Switch.scala 41:38:@20641.4]
  wire  _T_59484; // @[Switch.scala 41:52:@20643.4]
  wire  output_0_8; // @[Switch.scala 41:38:@20644.4]
  wire  _T_59487; // @[Switch.scala 41:52:@20646.4]
  wire  output_0_9; // @[Switch.scala 41:38:@20647.4]
  wire  _T_59490; // @[Switch.scala 41:52:@20649.4]
  wire  output_0_10; // @[Switch.scala 41:38:@20650.4]
  wire  _T_59493; // @[Switch.scala 41:52:@20652.4]
  wire  output_0_11; // @[Switch.scala 41:38:@20653.4]
  wire  _T_59496; // @[Switch.scala 41:52:@20655.4]
  wire  output_0_12; // @[Switch.scala 41:38:@20656.4]
  wire  _T_59499; // @[Switch.scala 41:52:@20658.4]
  wire  output_0_13; // @[Switch.scala 41:38:@20659.4]
  wire  _T_59502; // @[Switch.scala 41:52:@20661.4]
  wire  output_0_14; // @[Switch.scala 41:38:@20662.4]
  wire  _T_59505; // @[Switch.scala 41:52:@20664.4]
  wire  output_0_15; // @[Switch.scala 41:38:@20665.4]
  wire  _T_59508; // @[Switch.scala 41:52:@20667.4]
  wire  output_0_16; // @[Switch.scala 41:38:@20668.4]
  wire  _T_59511; // @[Switch.scala 41:52:@20670.4]
  wire  output_0_17; // @[Switch.scala 41:38:@20671.4]
  wire  _T_59514; // @[Switch.scala 41:52:@20673.4]
  wire  output_0_18; // @[Switch.scala 41:38:@20674.4]
  wire  _T_59517; // @[Switch.scala 41:52:@20676.4]
  wire  output_0_19; // @[Switch.scala 41:38:@20677.4]
  wire  _T_59520; // @[Switch.scala 41:52:@20679.4]
  wire  output_0_20; // @[Switch.scala 41:38:@20680.4]
  wire  _T_59523; // @[Switch.scala 41:52:@20682.4]
  wire  output_0_21; // @[Switch.scala 41:38:@20683.4]
  wire  _T_59526; // @[Switch.scala 41:52:@20685.4]
  wire  output_0_22; // @[Switch.scala 41:38:@20686.4]
  wire  _T_59529; // @[Switch.scala 41:52:@20688.4]
  wire  output_0_23; // @[Switch.scala 41:38:@20689.4]
  wire  _T_59532; // @[Switch.scala 41:52:@20691.4]
  wire  output_0_24; // @[Switch.scala 41:38:@20692.4]
  wire  _T_59535; // @[Switch.scala 41:52:@20694.4]
  wire  output_0_25; // @[Switch.scala 41:38:@20695.4]
  wire  _T_59538; // @[Switch.scala 41:52:@20697.4]
  wire  output_0_26; // @[Switch.scala 41:38:@20698.4]
  wire  _T_59541; // @[Switch.scala 41:52:@20700.4]
  wire  output_0_27; // @[Switch.scala 41:38:@20701.4]
  wire  _T_59544; // @[Switch.scala 41:52:@20703.4]
  wire  output_0_28; // @[Switch.scala 41:38:@20704.4]
  wire  _T_59547; // @[Switch.scala 41:52:@20706.4]
  wire  output_0_29; // @[Switch.scala 41:38:@20707.4]
  wire  _T_59550; // @[Switch.scala 41:52:@20709.4]
  wire  output_0_30; // @[Switch.scala 41:38:@20710.4]
  wire  _T_59553; // @[Switch.scala 41:52:@20712.4]
  wire  output_0_31; // @[Switch.scala 41:38:@20713.4]
  wire  _T_59556; // @[Switch.scala 41:52:@20715.4]
  wire  output_0_32; // @[Switch.scala 41:38:@20716.4]
  wire  _T_59559; // @[Switch.scala 41:52:@20718.4]
  wire  output_0_33; // @[Switch.scala 41:38:@20719.4]
  wire  _T_59562; // @[Switch.scala 41:52:@20721.4]
  wire  output_0_34; // @[Switch.scala 41:38:@20722.4]
  wire  _T_59565; // @[Switch.scala 41:52:@20724.4]
  wire  output_0_35; // @[Switch.scala 41:38:@20725.4]
  wire  _T_59568; // @[Switch.scala 41:52:@20727.4]
  wire  output_0_36; // @[Switch.scala 41:38:@20728.4]
  wire  _T_59571; // @[Switch.scala 41:52:@20730.4]
  wire  output_0_37; // @[Switch.scala 41:38:@20731.4]
  wire  _T_59574; // @[Switch.scala 41:52:@20733.4]
  wire  output_0_38; // @[Switch.scala 41:38:@20734.4]
  wire  _T_59577; // @[Switch.scala 41:52:@20736.4]
  wire  output_0_39; // @[Switch.scala 41:38:@20737.4]
  wire  _T_59580; // @[Switch.scala 41:52:@20739.4]
  wire  output_0_40; // @[Switch.scala 41:38:@20740.4]
  wire  _T_59583; // @[Switch.scala 41:52:@20742.4]
  wire  output_0_41; // @[Switch.scala 41:38:@20743.4]
  wire  _T_59586; // @[Switch.scala 41:52:@20745.4]
  wire  output_0_42; // @[Switch.scala 41:38:@20746.4]
  wire  _T_59589; // @[Switch.scala 41:52:@20748.4]
  wire  output_0_43; // @[Switch.scala 41:38:@20749.4]
  wire  _T_59592; // @[Switch.scala 41:52:@20751.4]
  wire  output_0_44; // @[Switch.scala 41:38:@20752.4]
  wire  _T_59595; // @[Switch.scala 41:52:@20754.4]
  wire  output_0_45; // @[Switch.scala 41:38:@20755.4]
  wire  _T_59598; // @[Switch.scala 41:52:@20757.4]
  wire  output_0_46; // @[Switch.scala 41:38:@20758.4]
  wire  _T_59601; // @[Switch.scala 41:52:@20760.4]
  wire  output_0_47; // @[Switch.scala 41:38:@20761.4]
  wire  _T_59604; // @[Switch.scala 41:52:@20763.4]
  wire  output_0_48; // @[Switch.scala 41:38:@20764.4]
  wire  _T_59607; // @[Switch.scala 41:52:@20766.4]
  wire  output_0_49; // @[Switch.scala 41:38:@20767.4]
  wire  _T_59610; // @[Switch.scala 41:52:@20769.4]
  wire  output_0_50; // @[Switch.scala 41:38:@20770.4]
  wire  _T_59613; // @[Switch.scala 41:52:@20772.4]
  wire  output_0_51; // @[Switch.scala 41:38:@20773.4]
  wire  _T_59616; // @[Switch.scala 41:52:@20775.4]
  wire  output_0_52; // @[Switch.scala 41:38:@20776.4]
  wire  _T_59619; // @[Switch.scala 41:52:@20778.4]
  wire  output_0_53; // @[Switch.scala 41:38:@20779.4]
  wire  _T_59622; // @[Switch.scala 41:52:@20781.4]
  wire  output_0_54; // @[Switch.scala 41:38:@20782.4]
  wire  _T_59625; // @[Switch.scala 41:52:@20784.4]
  wire  output_0_55; // @[Switch.scala 41:38:@20785.4]
  wire  _T_59628; // @[Switch.scala 41:52:@20787.4]
  wire  output_0_56; // @[Switch.scala 41:38:@20788.4]
  wire  _T_59631; // @[Switch.scala 41:52:@20790.4]
  wire  output_0_57; // @[Switch.scala 41:38:@20791.4]
  wire  _T_59634; // @[Switch.scala 41:52:@20793.4]
  wire  output_0_58; // @[Switch.scala 41:38:@20794.4]
  wire  _T_59637; // @[Switch.scala 41:52:@20796.4]
  wire  output_0_59; // @[Switch.scala 41:38:@20797.4]
  wire  _T_59640; // @[Switch.scala 41:52:@20799.4]
  wire  output_0_60; // @[Switch.scala 41:38:@20800.4]
  wire  _T_59643; // @[Switch.scala 41:52:@20802.4]
  wire  output_0_61; // @[Switch.scala 41:38:@20803.4]
  wire  _T_59646; // @[Switch.scala 41:52:@20805.4]
  wire  output_0_62; // @[Switch.scala 41:38:@20806.4]
  wire  _T_59649; // @[Switch.scala 41:52:@20808.4]
  wire  output_0_63; // @[Switch.scala 41:38:@20809.4]
  wire [7:0] _T_59657; // @[Switch.scala 43:31:@20817.4]
  wire [15:0] _T_59665; // @[Switch.scala 43:31:@20825.4]
  wire [7:0] _T_59672; // @[Switch.scala 43:31:@20832.4]
  wire [31:0] _T_59681; // @[Switch.scala 43:31:@20841.4]
  wire [7:0] _T_59688; // @[Switch.scala 43:31:@20848.4]
  wire [15:0] _T_59696; // @[Switch.scala 43:31:@20856.4]
  wire [7:0] _T_59703; // @[Switch.scala 43:31:@20863.4]
  wire [31:0] _T_59712; // @[Switch.scala 43:31:@20872.4]
  wire [63:0] _T_59713; // @[Switch.scala 43:31:@20873.4]
  wire  _T_59717; // @[Switch.scala 41:52:@20876.4]
  wire  output_1_0; // @[Switch.scala 41:38:@20877.4]
  wire  _T_59720; // @[Switch.scala 41:52:@20879.4]
  wire  output_1_1; // @[Switch.scala 41:38:@20880.4]
  wire  _T_59723; // @[Switch.scala 41:52:@20882.4]
  wire  output_1_2; // @[Switch.scala 41:38:@20883.4]
  wire  _T_59726; // @[Switch.scala 41:52:@20885.4]
  wire  output_1_3; // @[Switch.scala 41:38:@20886.4]
  wire  _T_59729; // @[Switch.scala 41:52:@20888.4]
  wire  output_1_4; // @[Switch.scala 41:38:@20889.4]
  wire  _T_59732; // @[Switch.scala 41:52:@20891.4]
  wire  output_1_5; // @[Switch.scala 41:38:@20892.4]
  wire  _T_59735; // @[Switch.scala 41:52:@20894.4]
  wire  output_1_6; // @[Switch.scala 41:38:@20895.4]
  wire  _T_59738; // @[Switch.scala 41:52:@20897.4]
  wire  output_1_7; // @[Switch.scala 41:38:@20898.4]
  wire  _T_59741; // @[Switch.scala 41:52:@20900.4]
  wire  output_1_8; // @[Switch.scala 41:38:@20901.4]
  wire  _T_59744; // @[Switch.scala 41:52:@20903.4]
  wire  output_1_9; // @[Switch.scala 41:38:@20904.4]
  wire  _T_59747; // @[Switch.scala 41:52:@20906.4]
  wire  output_1_10; // @[Switch.scala 41:38:@20907.4]
  wire  _T_59750; // @[Switch.scala 41:52:@20909.4]
  wire  output_1_11; // @[Switch.scala 41:38:@20910.4]
  wire  _T_59753; // @[Switch.scala 41:52:@20912.4]
  wire  output_1_12; // @[Switch.scala 41:38:@20913.4]
  wire  _T_59756; // @[Switch.scala 41:52:@20915.4]
  wire  output_1_13; // @[Switch.scala 41:38:@20916.4]
  wire  _T_59759; // @[Switch.scala 41:52:@20918.4]
  wire  output_1_14; // @[Switch.scala 41:38:@20919.4]
  wire  _T_59762; // @[Switch.scala 41:52:@20921.4]
  wire  output_1_15; // @[Switch.scala 41:38:@20922.4]
  wire  _T_59765; // @[Switch.scala 41:52:@20924.4]
  wire  output_1_16; // @[Switch.scala 41:38:@20925.4]
  wire  _T_59768; // @[Switch.scala 41:52:@20927.4]
  wire  output_1_17; // @[Switch.scala 41:38:@20928.4]
  wire  _T_59771; // @[Switch.scala 41:52:@20930.4]
  wire  output_1_18; // @[Switch.scala 41:38:@20931.4]
  wire  _T_59774; // @[Switch.scala 41:52:@20933.4]
  wire  output_1_19; // @[Switch.scala 41:38:@20934.4]
  wire  _T_59777; // @[Switch.scala 41:52:@20936.4]
  wire  output_1_20; // @[Switch.scala 41:38:@20937.4]
  wire  _T_59780; // @[Switch.scala 41:52:@20939.4]
  wire  output_1_21; // @[Switch.scala 41:38:@20940.4]
  wire  _T_59783; // @[Switch.scala 41:52:@20942.4]
  wire  output_1_22; // @[Switch.scala 41:38:@20943.4]
  wire  _T_59786; // @[Switch.scala 41:52:@20945.4]
  wire  output_1_23; // @[Switch.scala 41:38:@20946.4]
  wire  _T_59789; // @[Switch.scala 41:52:@20948.4]
  wire  output_1_24; // @[Switch.scala 41:38:@20949.4]
  wire  _T_59792; // @[Switch.scala 41:52:@20951.4]
  wire  output_1_25; // @[Switch.scala 41:38:@20952.4]
  wire  _T_59795; // @[Switch.scala 41:52:@20954.4]
  wire  output_1_26; // @[Switch.scala 41:38:@20955.4]
  wire  _T_59798; // @[Switch.scala 41:52:@20957.4]
  wire  output_1_27; // @[Switch.scala 41:38:@20958.4]
  wire  _T_59801; // @[Switch.scala 41:52:@20960.4]
  wire  output_1_28; // @[Switch.scala 41:38:@20961.4]
  wire  _T_59804; // @[Switch.scala 41:52:@20963.4]
  wire  output_1_29; // @[Switch.scala 41:38:@20964.4]
  wire  _T_59807; // @[Switch.scala 41:52:@20966.4]
  wire  output_1_30; // @[Switch.scala 41:38:@20967.4]
  wire  _T_59810; // @[Switch.scala 41:52:@20969.4]
  wire  output_1_31; // @[Switch.scala 41:38:@20970.4]
  wire  _T_59813; // @[Switch.scala 41:52:@20972.4]
  wire  output_1_32; // @[Switch.scala 41:38:@20973.4]
  wire  _T_59816; // @[Switch.scala 41:52:@20975.4]
  wire  output_1_33; // @[Switch.scala 41:38:@20976.4]
  wire  _T_59819; // @[Switch.scala 41:52:@20978.4]
  wire  output_1_34; // @[Switch.scala 41:38:@20979.4]
  wire  _T_59822; // @[Switch.scala 41:52:@20981.4]
  wire  output_1_35; // @[Switch.scala 41:38:@20982.4]
  wire  _T_59825; // @[Switch.scala 41:52:@20984.4]
  wire  output_1_36; // @[Switch.scala 41:38:@20985.4]
  wire  _T_59828; // @[Switch.scala 41:52:@20987.4]
  wire  output_1_37; // @[Switch.scala 41:38:@20988.4]
  wire  _T_59831; // @[Switch.scala 41:52:@20990.4]
  wire  output_1_38; // @[Switch.scala 41:38:@20991.4]
  wire  _T_59834; // @[Switch.scala 41:52:@20993.4]
  wire  output_1_39; // @[Switch.scala 41:38:@20994.4]
  wire  _T_59837; // @[Switch.scala 41:52:@20996.4]
  wire  output_1_40; // @[Switch.scala 41:38:@20997.4]
  wire  _T_59840; // @[Switch.scala 41:52:@20999.4]
  wire  output_1_41; // @[Switch.scala 41:38:@21000.4]
  wire  _T_59843; // @[Switch.scala 41:52:@21002.4]
  wire  output_1_42; // @[Switch.scala 41:38:@21003.4]
  wire  _T_59846; // @[Switch.scala 41:52:@21005.4]
  wire  output_1_43; // @[Switch.scala 41:38:@21006.4]
  wire  _T_59849; // @[Switch.scala 41:52:@21008.4]
  wire  output_1_44; // @[Switch.scala 41:38:@21009.4]
  wire  _T_59852; // @[Switch.scala 41:52:@21011.4]
  wire  output_1_45; // @[Switch.scala 41:38:@21012.4]
  wire  _T_59855; // @[Switch.scala 41:52:@21014.4]
  wire  output_1_46; // @[Switch.scala 41:38:@21015.4]
  wire  _T_59858; // @[Switch.scala 41:52:@21017.4]
  wire  output_1_47; // @[Switch.scala 41:38:@21018.4]
  wire  _T_59861; // @[Switch.scala 41:52:@21020.4]
  wire  output_1_48; // @[Switch.scala 41:38:@21021.4]
  wire  _T_59864; // @[Switch.scala 41:52:@21023.4]
  wire  output_1_49; // @[Switch.scala 41:38:@21024.4]
  wire  _T_59867; // @[Switch.scala 41:52:@21026.4]
  wire  output_1_50; // @[Switch.scala 41:38:@21027.4]
  wire  _T_59870; // @[Switch.scala 41:52:@21029.4]
  wire  output_1_51; // @[Switch.scala 41:38:@21030.4]
  wire  _T_59873; // @[Switch.scala 41:52:@21032.4]
  wire  output_1_52; // @[Switch.scala 41:38:@21033.4]
  wire  _T_59876; // @[Switch.scala 41:52:@21035.4]
  wire  output_1_53; // @[Switch.scala 41:38:@21036.4]
  wire  _T_59879; // @[Switch.scala 41:52:@21038.4]
  wire  output_1_54; // @[Switch.scala 41:38:@21039.4]
  wire  _T_59882; // @[Switch.scala 41:52:@21041.4]
  wire  output_1_55; // @[Switch.scala 41:38:@21042.4]
  wire  _T_59885; // @[Switch.scala 41:52:@21044.4]
  wire  output_1_56; // @[Switch.scala 41:38:@21045.4]
  wire  _T_59888; // @[Switch.scala 41:52:@21047.4]
  wire  output_1_57; // @[Switch.scala 41:38:@21048.4]
  wire  _T_59891; // @[Switch.scala 41:52:@21050.4]
  wire  output_1_58; // @[Switch.scala 41:38:@21051.4]
  wire  _T_59894; // @[Switch.scala 41:52:@21053.4]
  wire  output_1_59; // @[Switch.scala 41:38:@21054.4]
  wire  _T_59897; // @[Switch.scala 41:52:@21056.4]
  wire  output_1_60; // @[Switch.scala 41:38:@21057.4]
  wire  _T_59900; // @[Switch.scala 41:52:@21059.4]
  wire  output_1_61; // @[Switch.scala 41:38:@21060.4]
  wire  _T_59903; // @[Switch.scala 41:52:@21062.4]
  wire  output_1_62; // @[Switch.scala 41:38:@21063.4]
  wire  _T_59906; // @[Switch.scala 41:52:@21065.4]
  wire  output_1_63; // @[Switch.scala 41:38:@21066.4]
  wire [7:0] _T_59914; // @[Switch.scala 43:31:@21074.4]
  wire [15:0] _T_59922; // @[Switch.scala 43:31:@21082.4]
  wire [7:0] _T_59929; // @[Switch.scala 43:31:@21089.4]
  wire [31:0] _T_59938; // @[Switch.scala 43:31:@21098.4]
  wire [7:0] _T_59945; // @[Switch.scala 43:31:@21105.4]
  wire [15:0] _T_59953; // @[Switch.scala 43:31:@21113.4]
  wire [7:0] _T_59960; // @[Switch.scala 43:31:@21120.4]
  wire [31:0] _T_59969; // @[Switch.scala 43:31:@21129.4]
  wire [63:0] _T_59970; // @[Switch.scala 43:31:@21130.4]
  wire  _T_59974; // @[Switch.scala 41:52:@21133.4]
  wire  output_2_0; // @[Switch.scala 41:38:@21134.4]
  wire  _T_59977; // @[Switch.scala 41:52:@21136.4]
  wire  output_2_1; // @[Switch.scala 41:38:@21137.4]
  wire  _T_59980; // @[Switch.scala 41:52:@21139.4]
  wire  output_2_2; // @[Switch.scala 41:38:@21140.4]
  wire  _T_59983; // @[Switch.scala 41:52:@21142.4]
  wire  output_2_3; // @[Switch.scala 41:38:@21143.4]
  wire  _T_59986; // @[Switch.scala 41:52:@21145.4]
  wire  output_2_4; // @[Switch.scala 41:38:@21146.4]
  wire  _T_59989; // @[Switch.scala 41:52:@21148.4]
  wire  output_2_5; // @[Switch.scala 41:38:@21149.4]
  wire  _T_59992; // @[Switch.scala 41:52:@21151.4]
  wire  output_2_6; // @[Switch.scala 41:38:@21152.4]
  wire  _T_59995; // @[Switch.scala 41:52:@21154.4]
  wire  output_2_7; // @[Switch.scala 41:38:@21155.4]
  wire  _T_59998; // @[Switch.scala 41:52:@21157.4]
  wire  output_2_8; // @[Switch.scala 41:38:@21158.4]
  wire  _T_60001; // @[Switch.scala 41:52:@21160.4]
  wire  output_2_9; // @[Switch.scala 41:38:@21161.4]
  wire  _T_60004; // @[Switch.scala 41:52:@21163.4]
  wire  output_2_10; // @[Switch.scala 41:38:@21164.4]
  wire  _T_60007; // @[Switch.scala 41:52:@21166.4]
  wire  output_2_11; // @[Switch.scala 41:38:@21167.4]
  wire  _T_60010; // @[Switch.scala 41:52:@21169.4]
  wire  output_2_12; // @[Switch.scala 41:38:@21170.4]
  wire  _T_60013; // @[Switch.scala 41:52:@21172.4]
  wire  output_2_13; // @[Switch.scala 41:38:@21173.4]
  wire  _T_60016; // @[Switch.scala 41:52:@21175.4]
  wire  output_2_14; // @[Switch.scala 41:38:@21176.4]
  wire  _T_60019; // @[Switch.scala 41:52:@21178.4]
  wire  output_2_15; // @[Switch.scala 41:38:@21179.4]
  wire  _T_60022; // @[Switch.scala 41:52:@21181.4]
  wire  output_2_16; // @[Switch.scala 41:38:@21182.4]
  wire  _T_60025; // @[Switch.scala 41:52:@21184.4]
  wire  output_2_17; // @[Switch.scala 41:38:@21185.4]
  wire  _T_60028; // @[Switch.scala 41:52:@21187.4]
  wire  output_2_18; // @[Switch.scala 41:38:@21188.4]
  wire  _T_60031; // @[Switch.scala 41:52:@21190.4]
  wire  output_2_19; // @[Switch.scala 41:38:@21191.4]
  wire  _T_60034; // @[Switch.scala 41:52:@21193.4]
  wire  output_2_20; // @[Switch.scala 41:38:@21194.4]
  wire  _T_60037; // @[Switch.scala 41:52:@21196.4]
  wire  output_2_21; // @[Switch.scala 41:38:@21197.4]
  wire  _T_60040; // @[Switch.scala 41:52:@21199.4]
  wire  output_2_22; // @[Switch.scala 41:38:@21200.4]
  wire  _T_60043; // @[Switch.scala 41:52:@21202.4]
  wire  output_2_23; // @[Switch.scala 41:38:@21203.4]
  wire  _T_60046; // @[Switch.scala 41:52:@21205.4]
  wire  output_2_24; // @[Switch.scala 41:38:@21206.4]
  wire  _T_60049; // @[Switch.scala 41:52:@21208.4]
  wire  output_2_25; // @[Switch.scala 41:38:@21209.4]
  wire  _T_60052; // @[Switch.scala 41:52:@21211.4]
  wire  output_2_26; // @[Switch.scala 41:38:@21212.4]
  wire  _T_60055; // @[Switch.scala 41:52:@21214.4]
  wire  output_2_27; // @[Switch.scala 41:38:@21215.4]
  wire  _T_60058; // @[Switch.scala 41:52:@21217.4]
  wire  output_2_28; // @[Switch.scala 41:38:@21218.4]
  wire  _T_60061; // @[Switch.scala 41:52:@21220.4]
  wire  output_2_29; // @[Switch.scala 41:38:@21221.4]
  wire  _T_60064; // @[Switch.scala 41:52:@21223.4]
  wire  output_2_30; // @[Switch.scala 41:38:@21224.4]
  wire  _T_60067; // @[Switch.scala 41:52:@21226.4]
  wire  output_2_31; // @[Switch.scala 41:38:@21227.4]
  wire  _T_60070; // @[Switch.scala 41:52:@21229.4]
  wire  output_2_32; // @[Switch.scala 41:38:@21230.4]
  wire  _T_60073; // @[Switch.scala 41:52:@21232.4]
  wire  output_2_33; // @[Switch.scala 41:38:@21233.4]
  wire  _T_60076; // @[Switch.scala 41:52:@21235.4]
  wire  output_2_34; // @[Switch.scala 41:38:@21236.4]
  wire  _T_60079; // @[Switch.scala 41:52:@21238.4]
  wire  output_2_35; // @[Switch.scala 41:38:@21239.4]
  wire  _T_60082; // @[Switch.scala 41:52:@21241.4]
  wire  output_2_36; // @[Switch.scala 41:38:@21242.4]
  wire  _T_60085; // @[Switch.scala 41:52:@21244.4]
  wire  output_2_37; // @[Switch.scala 41:38:@21245.4]
  wire  _T_60088; // @[Switch.scala 41:52:@21247.4]
  wire  output_2_38; // @[Switch.scala 41:38:@21248.4]
  wire  _T_60091; // @[Switch.scala 41:52:@21250.4]
  wire  output_2_39; // @[Switch.scala 41:38:@21251.4]
  wire  _T_60094; // @[Switch.scala 41:52:@21253.4]
  wire  output_2_40; // @[Switch.scala 41:38:@21254.4]
  wire  _T_60097; // @[Switch.scala 41:52:@21256.4]
  wire  output_2_41; // @[Switch.scala 41:38:@21257.4]
  wire  _T_60100; // @[Switch.scala 41:52:@21259.4]
  wire  output_2_42; // @[Switch.scala 41:38:@21260.4]
  wire  _T_60103; // @[Switch.scala 41:52:@21262.4]
  wire  output_2_43; // @[Switch.scala 41:38:@21263.4]
  wire  _T_60106; // @[Switch.scala 41:52:@21265.4]
  wire  output_2_44; // @[Switch.scala 41:38:@21266.4]
  wire  _T_60109; // @[Switch.scala 41:52:@21268.4]
  wire  output_2_45; // @[Switch.scala 41:38:@21269.4]
  wire  _T_60112; // @[Switch.scala 41:52:@21271.4]
  wire  output_2_46; // @[Switch.scala 41:38:@21272.4]
  wire  _T_60115; // @[Switch.scala 41:52:@21274.4]
  wire  output_2_47; // @[Switch.scala 41:38:@21275.4]
  wire  _T_60118; // @[Switch.scala 41:52:@21277.4]
  wire  output_2_48; // @[Switch.scala 41:38:@21278.4]
  wire  _T_60121; // @[Switch.scala 41:52:@21280.4]
  wire  output_2_49; // @[Switch.scala 41:38:@21281.4]
  wire  _T_60124; // @[Switch.scala 41:52:@21283.4]
  wire  output_2_50; // @[Switch.scala 41:38:@21284.4]
  wire  _T_60127; // @[Switch.scala 41:52:@21286.4]
  wire  output_2_51; // @[Switch.scala 41:38:@21287.4]
  wire  _T_60130; // @[Switch.scala 41:52:@21289.4]
  wire  output_2_52; // @[Switch.scala 41:38:@21290.4]
  wire  _T_60133; // @[Switch.scala 41:52:@21292.4]
  wire  output_2_53; // @[Switch.scala 41:38:@21293.4]
  wire  _T_60136; // @[Switch.scala 41:52:@21295.4]
  wire  output_2_54; // @[Switch.scala 41:38:@21296.4]
  wire  _T_60139; // @[Switch.scala 41:52:@21298.4]
  wire  output_2_55; // @[Switch.scala 41:38:@21299.4]
  wire  _T_60142; // @[Switch.scala 41:52:@21301.4]
  wire  output_2_56; // @[Switch.scala 41:38:@21302.4]
  wire  _T_60145; // @[Switch.scala 41:52:@21304.4]
  wire  output_2_57; // @[Switch.scala 41:38:@21305.4]
  wire  _T_60148; // @[Switch.scala 41:52:@21307.4]
  wire  output_2_58; // @[Switch.scala 41:38:@21308.4]
  wire  _T_60151; // @[Switch.scala 41:52:@21310.4]
  wire  output_2_59; // @[Switch.scala 41:38:@21311.4]
  wire  _T_60154; // @[Switch.scala 41:52:@21313.4]
  wire  output_2_60; // @[Switch.scala 41:38:@21314.4]
  wire  _T_60157; // @[Switch.scala 41:52:@21316.4]
  wire  output_2_61; // @[Switch.scala 41:38:@21317.4]
  wire  _T_60160; // @[Switch.scala 41:52:@21319.4]
  wire  output_2_62; // @[Switch.scala 41:38:@21320.4]
  wire  _T_60163; // @[Switch.scala 41:52:@21322.4]
  wire  output_2_63; // @[Switch.scala 41:38:@21323.4]
  wire [7:0] _T_60171; // @[Switch.scala 43:31:@21331.4]
  wire [15:0] _T_60179; // @[Switch.scala 43:31:@21339.4]
  wire [7:0] _T_60186; // @[Switch.scala 43:31:@21346.4]
  wire [31:0] _T_60195; // @[Switch.scala 43:31:@21355.4]
  wire [7:0] _T_60202; // @[Switch.scala 43:31:@21362.4]
  wire [15:0] _T_60210; // @[Switch.scala 43:31:@21370.4]
  wire [7:0] _T_60217; // @[Switch.scala 43:31:@21377.4]
  wire [31:0] _T_60226; // @[Switch.scala 43:31:@21386.4]
  wire [63:0] _T_60227; // @[Switch.scala 43:31:@21387.4]
  wire  _T_60231; // @[Switch.scala 41:52:@21390.4]
  wire  output_3_0; // @[Switch.scala 41:38:@21391.4]
  wire  _T_60234; // @[Switch.scala 41:52:@21393.4]
  wire  output_3_1; // @[Switch.scala 41:38:@21394.4]
  wire  _T_60237; // @[Switch.scala 41:52:@21396.4]
  wire  output_3_2; // @[Switch.scala 41:38:@21397.4]
  wire  _T_60240; // @[Switch.scala 41:52:@21399.4]
  wire  output_3_3; // @[Switch.scala 41:38:@21400.4]
  wire  _T_60243; // @[Switch.scala 41:52:@21402.4]
  wire  output_3_4; // @[Switch.scala 41:38:@21403.4]
  wire  _T_60246; // @[Switch.scala 41:52:@21405.4]
  wire  output_3_5; // @[Switch.scala 41:38:@21406.4]
  wire  _T_60249; // @[Switch.scala 41:52:@21408.4]
  wire  output_3_6; // @[Switch.scala 41:38:@21409.4]
  wire  _T_60252; // @[Switch.scala 41:52:@21411.4]
  wire  output_3_7; // @[Switch.scala 41:38:@21412.4]
  wire  _T_60255; // @[Switch.scala 41:52:@21414.4]
  wire  output_3_8; // @[Switch.scala 41:38:@21415.4]
  wire  _T_60258; // @[Switch.scala 41:52:@21417.4]
  wire  output_3_9; // @[Switch.scala 41:38:@21418.4]
  wire  _T_60261; // @[Switch.scala 41:52:@21420.4]
  wire  output_3_10; // @[Switch.scala 41:38:@21421.4]
  wire  _T_60264; // @[Switch.scala 41:52:@21423.4]
  wire  output_3_11; // @[Switch.scala 41:38:@21424.4]
  wire  _T_60267; // @[Switch.scala 41:52:@21426.4]
  wire  output_3_12; // @[Switch.scala 41:38:@21427.4]
  wire  _T_60270; // @[Switch.scala 41:52:@21429.4]
  wire  output_3_13; // @[Switch.scala 41:38:@21430.4]
  wire  _T_60273; // @[Switch.scala 41:52:@21432.4]
  wire  output_3_14; // @[Switch.scala 41:38:@21433.4]
  wire  _T_60276; // @[Switch.scala 41:52:@21435.4]
  wire  output_3_15; // @[Switch.scala 41:38:@21436.4]
  wire  _T_60279; // @[Switch.scala 41:52:@21438.4]
  wire  output_3_16; // @[Switch.scala 41:38:@21439.4]
  wire  _T_60282; // @[Switch.scala 41:52:@21441.4]
  wire  output_3_17; // @[Switch.scala 41:38:@21442.4]
  wire  _T_60285; // @[Switch.scala 41:52:@21444.4]
  wire  output_3_18; // @[Switch.scala 41:38:@21445.4]
  wire  _T_60288; // @[Switch.scala 41:52:@21447.4]
  wire  output_3_19; // @[Switch.scala 41:38:@21448.4]
  wire  _T_60291; // @[Switch.scala 41:52:@21450.4]
  wire  output_3_20; // @[Switch.scala 41:38:@21451.4]
  wire  _T_60294; // @[Switch.scala 41:52:@21453.4]
  wire  output_3_21; // @[Switch.scala 41:38:@21454.4]
  wire  _T_60297; // @[Switch.scala 41:52:@21456.4]
  wire  output_3_22; // @[Switch.scala 41:38:@21457.4]
  wire  _T_60300; // @[Switch.scala 41:52:@21459.4]
  wire  output_3_23; // @[Switch.scala 41:38:@21460.4]
  wire  _T_60303; // @[Switch.scala 41:52:@21462.4]
  wire  output_3_24; // @[Switch.scala 41:38:@21463.4]
  wire  _T_60306; // @[Switch.scala 41:52:@21465.4]
  wire  output_3_25; // @[Switch.scala 41:38:@21466.4]
  wire  _T_60309; // @[Switch.scala 41:52:@21468.4]
  wire  output_3_26; // @[Switch.scala 41:38:@21469.4]
  wire  _T_60312; // @[Switch.scala 41:52:@21471.4]
  wire  output_3_27; // @[Switch.scala 41:38:@21472.4]
  wire  _T_60315; // @[Switch.scala 41:52:@21474.4]
  wire  output_3_28; // @[Switch.scala 41:38:@21475.4]
  wire  _T_60318; // @[Switch.scala 41:52:@21477.4]
  wire  output_3_29; // @[Switch.scala 41:38:@21478.4]
  wire  _T_60321; // @[Switch.scala 41:52:@21480.4]
  wire  output_3_30; // @[Switch.scala 41:38:@21481.4]
  wire  _T_60324; // @[Switch.scala 41:52:@21483.4]
  wire  output_3_31; // @[Switch.scala 41:38:@21484.4]
  wire  _T_60327; // @[Switch.scala 41:52:@21486.4]
  wire  output_3_32; // @[Switch.scala 41:38:@21487.4]
  wire  _T_60330; // @[Switch.scala 41:52:@21489.4]
  wire  output_3_33; // @[Switch.scala 41:38:@21490.4]
  wire  _T_60333; // @[Switch.scala 41:52:@21492.4]
  wire  output_3_34; // @[Switch.scala 41:38:@21493.4]
  wire  _T_60336; // @[Switch.scala 41:52:@21495.4]
  wire  output_3_35; // @[Switch.scala 41:38:@21496.4]
  wire  _T_60339; // @[Switch.scala 41:52:@21498.4]
  wire  output_3_36; // @[Switch.scala 41:38:@21499.4]
  wire  _T_60342; // @[Switch.scala 41:52:@21501.4]
  wire  output_3_37; // @[Switch.scala 41:38:@21502.4]
  wire  _T_60345; // @[Switch.scala 41:52:@21504.4]
  wire  output_3_38; // @[Switch.scala 41:38:@21505.4]
  wire  _T_60348; // @[Switch.scala 41:52:@21507.4]
  wire  output_3_39; // @[Switch.scala 41:38:@21508.4]
  wire  _T_60351; // @[Switch.scala 41:52:@21510.4]
  wire  output_3_40; // @[Switch.scala 41:38:@21511.4]
  wire  _T_60354; // @[Switch.scala 41:52:@21513.4]
  wire  output_3_41; // @[Switch.scala 41:38:@21514.4]
  wire  _T_60357; // @[Switch.scala 41:52:@21516.4]
  wire  output_3_42; // @[Switch.scala 41:38:@21517.4]
  wire  _T_60360; // @[Switch.scala 41:52:@21519.4]
  wire  output_3_43; // @[Switch.scala 41:38:@21520.4]
  wire  _T_60363; // @[Switch.scala 41:52:@21522.4]
  wire  output_3_44; // @[Switch.scala 41:38:@21523.4]
  wire  _T_60366; // @[Switch.scala 41:52:@21525.4]
  wire  output_3_45; // @[Switch.scala 41:38:@21526.4]
  wire  _T_60369; // @[Switch.scala 41:52:@21528.4]
  wire  output_3_46; // @[Switch.scala 41:38:@21529.4]
  wire  _T_60372; // @[Switch.scala 41:52:@21531.4]
  wire  output_3_47; // @[Switch.scala 41:38:@21532.4]
  wire  _T_60375; // @[Switch.scala 41:52:@21534.4]
  wire  output_3_48; // @[Switch.scala 41:38:@21535.4]
  wire  _T_60378; // @[Switch.scala 41:52:@21537.4]
  wire  output_3_49; // @[Switch.scala 41:38:@21538.4]
  wire  _T_60381; // @[Switch.scala 41:52:@21540.4]
  wire  output_3_50; // @[Switch.scala 41:38:@21541.4]
  wire  _T_60384; // @[Switch.scala 41:52:@21543.4]
  wire  output_3_51; // @[Switch.scala 41:38:@21544.4]
  wire  _T_60387; // @[Switch.scala 41:52:@21546.4]
  wire  output_3_52; // @[Switch.scala 41:38:@21547.4]
  wire  _T_60390; // @[Switch.scala 41:52:@21549.4]
  wire  output_3_53; // @[Switch.scala 41:38:@21550.4]
  wire  _T_60393; // @[Switch.scala 41:52:@21552.4]
  wire  output_3_54; // @[Switch.scala 41:38:@21553.4]
  wire  _T_60396; // @[Switch.scala 41:52:@21555.4]
  wire  output_3_55; // @[Switch.scala 41:38:@21556.4]
  wire  _T_60399; // @[Switch.scala 41:52:@21558.4]
  wire  output_3_56; // @[Switch.scala 41:38:@21559.4]
  wire  _T_60402; // @[Switch.scala 41:52:@21561.4]
  wire  output_3_57; // @[Switch.scala 41:38:@21562.4]
  wire  _T_60405; // @[Switch.scala 41:52:@21564.4]
  wire  output_3_58; // @[Switch.scala 41:38:@21565.4]
  wire  _T_60408; // @[Switch.scala 41:52:@21567.4]
  wire  output_3_59; // @[Switch.scala 41:38:@21568.4]
  wire  _T_60411; // @[Switch.scala 41:52:@21570.4]
  wire  output_3_60; // @[Switch.scala 41:38:@21571.4]
  wire  _T_60414; // @[Switch.scala 41:52:@21573.4]
  wire  output_3_61; // @[Switch.scala 41:38:@21574.4]
  wire  _T_60417; // @[Switch.scala 41:52:@21576.4]
  wire  output_3_62; // @[Switch.scala 41:38:@21577.4]
  wire  _T_60420; // @[Switch.scala 41:52:@21579.4]
  wire  output_3_63; // @[Switch.scala 41:38:@21580.4]
  wire [7:0] _T_60428; // @[Switch.scala 43:31:@21588.4]
  wire [15:0] _T_60436; // @[Switch.scala 43:31:@21596.4]
  wire [7:0] _T_60443; // @[Switch.scala 43:31:@21603.4]
  wire [31:0] _T_60452; // @[Switch.scala 43:31:@21612.4]
  wire [7:0] _T_60459; // @[Switch.scala 43:31:@21619.4]
  wire [15:0] _T_60467; // @[Switch.scala 43:31:@21627.4]
  wire [7:0] _T_60474; // @[Switch.scala 43:31:@21634.4]
  wire [31:0] _T_60483; // @[Switch.scala 43:31:@21643.4]
  wire [63:0] _T_60484; // @[Switch.scala 43:31:@21644.4]
  wire  _T_60488; // @[Switch.scala 41:52:@21647.4]
  wire  output_4_0; // @[Switch.scala 41:38:@21648.4]
  wire  _T_60491; // @[Switch.scala 41:52:@21650.4]
  wire  output_4_1; // @[Switch.scala 41:38:@21651.4]
  wire  _T_60494; // @[Switch.scala 41:52:@21653.4]
  wire  output_4_2; // @[Switch.scala 41:38:@21654.4]
  wire  _T_60497; // @[Switch.scala 41:52:@21656.4]
  wire  output_4_3; // @[Switch.scala 41:38:@21657.4]
  wire  _T_60500; // @[Switch.scala 41:52:@21659.4]
  wire  output_4_4; // @[Switch.scala 41:38:@21660.4]
  wire  _T_60503; // @[Switch.scala 41:52:@21662.4]
  wire  output_4_5; // @[Switch.scala 41:38:@21663.4]
  wire  _T_60506; // @[Switch.scala 41:52:@21665.4]
  wire  output_4_6; // @[Switch.scala 41:38:@21666.4]
  wire  _T_60509; // @[Switch.scala 41:52:@21668.4]
  wire  output_4_7; // @[Switch.scala 41:38:@21669.4]
  wire  _T_60512; // @[Switch.scala 41:52:@21671.4]
  wire  output_4_8; // @[Switch.scala 41:38:@21672.4]
  wire  _T_60515; // @[Switch.scala 41:52:@21674.4]
  wire  output_4_9; // @[Switch.scala 41:38:@21675.4]
  wire  _T_60518; // @[Switch.scala 41:52:@21677.4]
  wire  output_4_10; // @[Switch.scala 41:38:@21678.4]
  wire  _T_60521; // @[Switch.scala 41:52:@21680.4]
  wire  output_4_11; // @[Switch.scala 41:38:@21681.4]
  wire  _T_60524; // @[Switch.scala 41:52:@21683.4]
  wire  output_4_12; // @[Switch.scala 41:38:@21684.4]
  wire  _T_60527; // @[Switch.scala 41:52:@21686.4]
  wire  output_4_13; // @[Switch.scala 41:38:@21687.4]
  wire  _T_60530; // @[Switch.scala 41:52:@21689.4]
  wire  output_4_14; // @[Switch.scala 41:38:@21690.4]
  wire  _T_60533; // @[Switch.scala 41:52:@21692.4]
  wire  output_4_15; // @[Switch.scala 41:38:@21693.4]
  wire  _T_60536; // @[Switch.scala 41:52:@21695.4]
  wire  output_4_16; // @[Switch.scala 41:38:@21696.4]
  wire  _T_60539; // @[Switch.scala 41:52:@21698.4]
  wire  output_4_17; // @[Switch.scala 41:38:@21699.4]
  wire  _T_60542; // @[Switch.scala 41:52:@21701.4]
  wire  output_4_18; // @[Switch.scala 41:38:@21702.4]
  wire  _T_60545; // @[Switch.scala 41:52:@21704.4]
  wire  output_4_19; // @[Switch.scala 41:38:@21705.4]
  wire  _T_60548; // @[Switch.scala 41:52:@21707.4]
  wire  output_4_20; // @[Switch.scala 41:38:@21708.4]
  wire  _T_60551; // @[Switch.scala 41:52:@21710.4]
  wire  output_4_21; // @[Switch.scala 41:38:@21711.4]
  wire  _T_60554; // @[Switch.scala 41:52:@21713.4]
  wire  output_4_22; // @[Switch.scala 41:38:@21714.4]
  wire  _T_60557; // @[Switch.scala 41:52:@21716.4]
  wire  output_4_23; // @[Switch.scala 41:38:@21717.4]
  wire  _T_60560; // @[Switch.scala 41:52:@21719.4]
  wire  output_4_24; // @[Switch.scala 41:38:@21720.4]
  wire  _T_60563; // @[Switch.scala 41:52:@21722.4]
  wire  output_4_25; // @[Switch.scala 41:38:@21723.4]
  wire  _T_60566; // @[Switch.scala 41:52:@21725.4]
  wire  output_4_26; // @[Switch.scala 41:38:@21726.4]
  wire  _T_60569; // @[Switch.scala 41:52:@21728.4]
  wire  output_4_27; // @[Switch.scala 41:38:@21729.4]
  wire  _T_60572; // @[Switch.scala 41:52:@21731.4]
  wire  output_4_28; // @[Switch.scala 41:38:@21732.4]
  wire  _T_60575; // @[Switch.scala 41:52:@21734.4]
  wire  output_4_29; // @[Switch.scala 41:38:@21735.4]
  wire  _T_60578; // @[Switch.scala 41:52:@21737.4]
  wire  output_4_30; // @[Switch.scala 41:38:@21738.4]
  wire  _T_60581; // @[Switch.scala 41:52:@21740.4]
  wire  output_4_31; // @[Switch.scala 41:38:@21741.4]
  wire  _T_60584; // @[Switch.scala 41:52:@21743.4]
  wire  output_4_32; // @[Switch.scala 41:38:@21744.4]
  wire  _T_60587; // @[Switch.scala 41:52:@21746.4]
  wire  output_4_33; // @[Switch.scala 41:38:@21747.4]
  wire  _T_60590; // @[Switch.scala 41:52:@21749.4]
  wire  output_4_34; // @[Switch.scala 41:38:@21750.4]
  wire  _T_60593; // @[Switch.scala 41:52:@21752.4]
  wire  output_4_35; // @[Switch.scala 41:38:@21753.4]
  wire  _T_60596; // @[Switch.scala 41:52:@21755.4]
  wire  output_4_36; // @[Switch.scala 41:38:@21756.4]
  wire  _T_60599; // @[Switch.scala 41:52:@21758.4]
  wire  output_4_37; // @[Switch.scala 41:38:@21759.4]
  wire  _T_60602; // @[Switch.scala 41:52:@21761.4]
  wire  output_4_38; // @[Switch.scala 41:38:@21762.4]
  wire  _T_60605; // @[Switch.scala 41:52:@21764.4]
  wire  output_4_39; // @[Switch.scala 41:38:@21765.4]
  wire  _T_60608; // @[Switch.scala 41:52:@21767.4]
  wire  output_4_40; // @[Switch.scala 41:38:@21768.4]
  wire  _T_60611; // @[Switch.scala 41:52:@21770.4]
  wire  output_4_41; // @[Switch.scala 41:38:@21771.4]
  wire  _T_60614; // @[Switch.scala 41:52:@21773.4]
  wire  output_4_42; // @[Switch.scala 41:38:@21774.4]
  wire  _T_60617; // @[Switch.scala 41:52:@21776.4]
  wire  output_4_43; // @[Switch.scala 41:38:@21777.4]
  wire  _T_60620; // @[Switch.scala 41:52:@21779.4]
  wire  output_4_44; // @[Switch.scala 41:38:@21780.4]
  wire  _T_60623; // @[Switch.scala 41:52:@21782.4]
  wire  output_4_45; // @[Switch.scala 41:38:@21783.4]
  wire  _T_60626; // @[Switch.scala 41:52:@21785.4]
  wire  output_4_46; // @[Switch.scala 41:38:@21786.4]
  wire  _T_60629; // @[Switch.scala 41:52:@21788.4]
  wire  output_4_47; // @[Switch.scala 41:38:@21789.4]
  wire  _T_60632; // @[Switch.scala 41:52:@21791.4]
  wire  output_4_48; // @[Switch.scala 41:38:@21792.4]
  wire  _T_60635; // @[Switch.scala 41:52:@21794.4]
  wire  output_4_49; // @[Switch.scala 41:38:@21795.4]
  wire  _T_60638; // @[Switch.scala 41:52:@21797.4]
  wire  output_4_50; // @[Switch.scala 41:38:@21798.4]
  wire  _T_60641; // @[Switch.scala 41:52:@21800.4]
  wire  output_4_51; // @[Switch.scala 41:38:@21801.4]
  wire  _T_60644; // @[Switch.scala 41:52:@21803.4]
  wire  output_4_52; // @[Switch.scala 41:38:@21804.4]
  wire  _T_60647; // @[Switch.scala 41:52:@21806.4]
  wire  output_4_53; // @[Switch.scala 41:38:@21807.4]
  wire  _T_60650; // @[Switch.scala 41:52:@21809.4]
  wire  output_4_54; // @[Switch.scala 41:38:@21810.4]
  wire  _T_60653; // @[Switch.scala 41:52:@21812.4]
  wire  output_4_55; // @[Switch.scala 41:38:@21813.4]
  wire  _T_60656; // @[Switch.scala 41:52:@21815.4]
  wire  output_4_56; // @[Switch.scala 41:38:@21816.4]
  wire  _T_60659; // @[Switch.scala 41:52:@21818.4]
  wire  output_4_57; // @[Switch.scala 41:38:@21819.4]
  wire  _T_60662; // @[Switch.scala 41:52:@21821.4]
  wire  output_4_58; // @[Switch.scala 41:38:@21822.4]
  wire  _T_60665; // @[Switch.scala 41:52:@21824.4]
  wire  output_4_59; // @[Switch.scala 41:38:@21825.4]
  wire  _T_60668; // @[Switch.scala 41:52:@21827.4]
  wire  output_4_60; // @[Switch.scala 41:38:@21828.4]
  wire  _T_60671; // @[Switch.scala 41:52:@21830.4]
  wire  output_4_61; // @[Switch.scala 41:38:@21831.4]
  wire  _T_60674; // @[Switch.scala 41:52:@21833.4]
  wire  output_4_62; // @[Switch.scala 41:38:@21834.4]
  wire  _T_60677; // @[Switch.scala 41:52:@21836.4]
  wire  output_4_63; // @[Switch.scala 41:38:@21837.4]
  wire [7:0] _T_60685; // @[Switch.scala 43:31:@21845.4]
  wire [15:0] _T_60693; // @[Switch.scala 43:31:@21853.4]
  wire [7:0] _T_60700; // @[Switch.scala 43:31:@21860.4]
  wire [31:0] _T_60709; // @[Switch.scala 43:31:@21869.4]
  wire [7:0] _T_60716; // @[Switch.scala 43:31:@21876.4]
  wire [15:0] _T_60724; // @[Switch.scala 43:31:@21884.4]
  wire [7:0] _T_60731; // @[Switch.scala 43:31:@21891.4]
  wire [31:0] _T_60740; // @[Switch.scala 43:31:@21900.4]
  wire [63:0] _T_60741; // @[Switch.scala 43:31:@21901.4]
  wire  _T_60745; // @[Switch.scala 41:52:@21904.4]
  wire  output_5_0; // @[Switch.scala 41:38:@21905.4]
  wire  _T_60748; // @[Switch.scala 41:52:@21907.4]
  wire  output_5_1; // @[Switch.scala 41:38:@21908.4]
  wire  _T_60751; // @[Switch.scala 41:52:@21910.4]
  wire  output_5_2; // @[Switch.scala 41:38:@21911.4]
  wire  _T_60754; // @[Switch.scala 41:52:@21913.4]
  wire  output_5_3; // @[Switch.scala 41:38:@21914.4]
  wire  _T_60757; // @[Switch.scala 41:52:@21916.4]
  wire  output_5_4; // @[Switch.scala 41:38:@21917.4]
  wire  _T_60760; // @[Switch.scala 41:52:@21919.4]
  wire  output_5_5; // @[Switch.scala 41:38:@21920.4]
  wire  _T_60763; // @[Switch.scala 41:52:@21922.4]
  wire  output_5_6; // @[Switch.scala 41:38:@21923.4]
  wire  _T_60766; // @[Switch.scala 41:52:@21925.4]
  wire  output_5_7; // @[Switch.scala 41:38:@21926.4]
  wire  _T_60769; // @[Switch.scala 41:52:@21928.4]
  wire  output_5_8; // @[Switch.scala 41:38:@21929.4]
  wire  _T_60772; // @[Switch.scala 41:52:@21931.4]
  wire  output_5_9; // @[Switch.scala 41:38:@21932.4]
  wire  _T_60775; // @[Switch.scala 41:52:@21934.4]
  wire  output_5_10; // @[Switch.scala 41:38:@21935.4]
  wire  _T_60778; // @[Switch.scala 41:52:@21937.4]
  wire  output_5_11; // @[Switch.scala 41:38:@21938.4]
  wire  _T_60781; // @[Switch.scala 41:52:@21940.4]
  wire  output_5_12; // @[Switch.scala 41:38:@21941.4]
  wire  _T_60784; // @[Switch.scala 41:52:@21943.4]
  wire  output_5_13; // @[Switch.scala 41:38:@21944.4]
  wire  _T_60787; // @[Switch.scala 41:52:@21946.4]
  wire  output_5_14; // @[Switch.scala 41:38:@21947.4]
  wire  _T_60790; // @[Switch.scala 41:52:@21949.4]
  wire  output_5_15; // @[Switch.scala 41:38:@21950.4]
  wire  _T_60793; // @[Switch.scala 41:52:@21952.4]
  wire  output_5_16; // @[Switch.scala 41:38:@21953.4]
  wire  _T_60796; // @[Switch.scala 41:52:@21955.4]
  wire  output_5_17; // @[Switch.scala 41:38:@21956.4]
  wire  _T_60799; // @[Switch.scala 41:52:@21958.4]
  wire  output_5_18; // @[Switch.scala 41:38:@21959.4]
  wire  _T_60802; // @[Switch.scala 41:52:@21961.4]
  wire  output_5_19; // @[Switch.scala 41:38:@21962.4]
  wire  _T_60805; // @[Switch.scala 41:52:@21964.4]
  wire  output_5_20; // @[Switch.scala 41:38:@21965.4]
  wire  _T_60808; // @[Switch.scala 41:52:@21967.4]
  wire  output_5_21; // @[Switch.scala 41:38:@21968.4]
  wire  _T_60811; // @[Switch.scala 41:52:@21970.4]
  wire  output_5_22; // @[Switch.scala 41:38:@21971.4]
  wire  _T_60814; // @[Switch.scala 41:52:@21973.4]
  wire  output_5_23; // @[Switch.scala 41:38:@21974.4]
  wire  _T_60817; // @[Switch.scala 41:52:@21976.4]
  wire  output_5_24; // @[Switch.scala 41:38:@21977.4]
  wire  _T_60820; // @[Switch.scala 41:52:@21979.4]
  wire  output_5_25; // @[Switch.scala 41:38:@21980.4]
  wire  _T_60823; // @[Switch.scala 41:52:@21982.4]
  wire  output_5_26; // @[Switch.scala 41:38:@21983.4]
  wire  _T_60826; // @[Switch.scala 41:52:@21985.4]
  wire  output_5_27; // @[Switch.scala 41:38:@21986.4]
  wire  _T_60829; // @[Switch.scala 41:52:@21988.4]
  wire  output_5_28; // @[Switch.scala 41:38:@21989.4]
  wire  _T_60832; // @[Switch.scala 41:52:@21991.4]
  wire  output_5_29; // @[Switch.scala 41:38:@21992.4]
  wire  _T_60835; // @[Switch.scala 41:52:@21994.4]
  wire  output_5_30; // @[Switch.scala 41:38:@21995.4]
  wire  _T_60838; // @[Switch.scala 41:52:@21997.4]
  wire  output_5_31; // @[Switch.scala 41:38:@21998.4]
  wire  _T_60841; // @[Switch.scala 41:52:@22000.4]
  wire  output_5_32; // @[Switch.scala 41:38:@22001.4]
  wire  _T_60844; // @[Switch.scala 41:52:@22003.4]
  wire  output_5_33; // @[Switch.scala 41:38:@22004.4]
  wire  _T_60847; // @[Switch.scala 41:52:@22006.4]
  wire  output_5_34; // @[Switch.scala 41:38:@22007.4]
  wire  _T_60850; // @[Switch.scala 41:52:@22009.4]
  wire  output_5_35; // @[Switch.scala 41:38:@22010.4]
  wire  _T_60853; // @[Switch.scala 41:52:@22012.4]
  wire  output_5_36; // @[Switch.scala 41:38:@22013.4]
  wire  _T_60856; // @[Switch.scala 41:52:@22015.4]
  wire  output_5_37; // @[Switch.scala 41:38:@22016.4]
  wire  _T_60859; // @[Switch.scala 41:52:@22018.4]
  wire  output_5_38; // @[Switch.scala 41:38:@22019.4]
  wire  _T_60862; // @[Switch.scala 41:52:@22021.4]
  wire  output_5_39; // @[Switch.scala 41:38:@22022.4]
  wire  _T_60865; // @[Switch.scala 41:52:@22024.4]
  wire  output_5_40; // @[Switch.scala 41:38:@22025.4]
  wire  _T_60868; // @[Switch.scala 41:52:@22027.4]
  wire  output_5_41; // @[Switch.scala 41:38:@22028.4]
  wire  _T_60871; // @[Switch.scala 41:52:@22030.4]
  wire  output_5_42; // @[Switch.scala 41:38:@22031.4]
  wire  _T_60874; // @[Switch.scala 41:52:@22033.4]
  wire  output_5_43; // @[Switch.scala 41:38:@22034.4]
  wire  _T_60877; // @[Switch.scala 41:52:@22036.4]
  wire  output_5_44; // @[Switch.scala 41:38:@22037.4]
  wire  _T_60880; // @[Switch.scala 41:52:@22039.4]
  wire  output_5_45; // @[Switch.scala 41:38:@22040.4]
  wire  _T_60883; // @[Switch.scala 41:52:@22042.4]
  wire  output_5_46; // @[Switch.scala 41:38:@22043.4]
  wire  _T_60886; // @[Switch.scala 41:52:@22045.4]
  wire  output_5_47; // @[Switch.scala 41:38:@22046.4]
  wire  _T_60889; // @[Switch.scala 41:52:@22048.4]
  wire  output_5_48; // @[Switch.scala 41:38:@22049.4]
  wire  _T_60892; // @[Switch.scala 41:52:@22051.4]
  wire  output_5_49; // @[Switch.scala 41:38:@22052.4]
  wire  _T_60895; // @[Switch.scala 41:52:@22054.4]
  wire  output_5_50; // @[Switch.scala 41:38:@22055.4]
  wire  _T_60898; // @[Switch.scala 41:52:@22057.4]
  wire  output_5_51; // @[Switch.scala 41:38:@22058.4]
  wire  _T_60901; // @[Switch.scala 41:52:@22060.4]
  wire  output_5_52; // @[Switch.scala 41:38:@22061.4]
  wire  _T_60904; // @[Switch.scala 41:52:@22063.4]
  wire  output_5_53; // @[Switch.scala 41:38:@22064.4]
  wire  _T_60907; // @[Switch.scala 41:52:@22066.4]
  wire  output_5_54; // @[Switch.scala 41:38:@22067.4]
  wire  _T_60910; // @[Switch.scala 41:52:@22069.4]
  wire  output_5_55; // @[Switch.scala 41:38:@22070.4]
  wire  _T_60913; // @[Switch.scala 41:52:@22072.4]
  wire  output_5_56; // @[Switch.scala 41:38:@22073.4]
  wire  _T_60916; // @[Switch.scala 41:52:@22075.4]
  wire  output_5_57; // @[Switch.scala 41:38:@22076.4]
  wire  _T_60919; // @[Switch.scala 41:52:@22078.4]
  wire  output_5_58; // @[Switch.scala 41:38:@22079.4]
  wire  _T_60922; // @[Switch.scala 41:52:@22081.4]
  wire  output_5_59; // @[Switch.scala 41:38:@22082.4]
  wire  _T_60925; // @[Switch.scala 41:52:@22084.4]
  wire  output_5_60; // @[Switch.scala 41:38:@22085.4]
  wire  _T_60928; // @[Switch.scala 41:52:@22087.4]
  wire  output_5_61; // @[Switch.scala 41:38:@22088.4]
  wire  _T_60931; // @[Switch.scala 41:52:@22090.4]
  wire  output_5_62; // @[Switch.scala 41:38:@22091.4]
  wire  _T_60934; // @[Switch.scala 41:52:@22093.4]
  wire  output_5_63; // @[Switch.scala 41:38:@22094.4]
  wire [7:0] _T_60942; // @[Switch.scala 43:31:@22102.4]
  wire [15:0] _T_60950; // @[Switch.scala 43:31:@22110.4]
  wire [7:0] _T_60957; // @[Switch.scala 43:31:@22117.4]
  wire [31:0] _T_60966; // @[Switch.scala 43:31:@22126.4]
  wire [7:0] _T_60973; // @[Switch.scala 43:31:@22133.4]
  wire [15:0] _T_60981; // @[Switch.scala 43:31:@22141.4]
  wire [7:0] _T_60988; // @[Switch.scala 43:31:@22148.4]
  wire [31:0] _T_60997; // @[Switch.scala 43:31:@22157.4]
  wire [63:0] _T_60998; // @[Switch.scala 43:31:@22158.4]
  wire  _T_61002; // @[Switch.scala 41:52:@22161.4]
  wire  output_6_0; // @[Switch.scala 41:38:@22162.4]
  wire  _T_61005; // @[Switch.scala 41:52:@22164.4]
  wire  output_6_1; // @[Switch.scala 41:38:@22165.4]
  wire  _T_61008; // @[Switch.scala 41:52:@22167.4]
  wire  output_6_2; // @[Switch.scala 41:38:@22168.4]
  wire  _T_61011; // @[Switch.scala 41:52:@22170.4]
  wire  output_6_3; // @[Switch.scala 41:38:@22171.4]
  wire  _T_61014; // @[Switch.scala 41:52:@22173.4]
  wire  output_6_4; // @[Switch.scala 41:38:@22174.4]
  wire  _T_61017; // @[Switch.scala 41:52:@22176.4]
  wire  output_6_5; // @[Switch.scala 41:38:@22177.4]
  wire  _T_61020; // @[Switch.scala 41:52:@22179.4]
  wire  output_6_6; // @[Switch.scala 41:38:@22180.4]
  wire  _T_61023; // @[Switch.scala 41:52:@22182.4]
  wire  output_6_7; // @[Switch.scala 41:38:@22183.4]
  wire  _T_61026; // @[Switch.scala 41:52:@22185.4]
  wire  output_6_8; // @[Switch.scala 41:38:@22186.4]
  wire  _T_61029; // @[Switch.scala 41:52:@22188.4]
  wire  output_6_9; // @[Switch.scala 41:38:@22189.4]
  wire  _T_61032; // @[Switch.scala 41:52:@22191.4]
  wire  output_6_10; // @[Switch.scala 41:38:@22192.4]
  wire  _T_61035; // @[Switch.scala 41:52:@22194.4]
  wire  output_6_11; // @[Switch.scala 41:38:@22195.4]
  wire  _T_61038; // @[Switch.scala 41:52:@22197.4]
  wire  output_6_12; // @[Switch.scala 41:38:@22198.4]
  wire  _T_61041; // @[Switch.scala 41:52:@22200.4]
  wire  output_6_13; // @[Switch.scala 41:38:@22201.4]
  wire  _T_61044; // @[Switch.scala 41:52:@22203.4]
  wire  output_6_14; // @[Switch.scala 41:38:@22204.4]
  wire  _T_61047; // @[Switch.scala 41:52:@22206.4]
  wire  output_6_15; // @[Switch.scala 41:38:@22207.4]
  wire  _T_61050; // @[Switch.scala 41:52:@22209.4]
  wire  output_6_16; // @[Switch.scala 41:38:@22210.4]
  wire  _T_61053; // @[Switch.scala 41:52:@22212.4]
  wire  output_6_17; // @[Switch.scala 41:38:@22213.4]
  wire  _T_61056; // @[Switch.scala 41:52:@22215.4]
  wire  output_6_18; // @[Switch.scala 41:38:@22216.4]
  wire  _T_61059; // @[Switch.scala 41:52:@22218.4]
  wire  output_6_19; // @[Switch.scala 41:38:@22219.4]
  wire  _T_61062; // @[Switch.scala 41:52:@22221.4]
  wire  output_6_20; // @[Switch.scala 41:38:@22222.4]
  wire  _T_61065; // @[Switch.scala 41:52:@22224.4]
  wire  output_6_21; // @[Switch.scala 41:38:@22225.4]
  wire  _T_61068; // @[Switch.scala 41:52:@22227.4]
  wire  output_6_22; // @[Switch.scala 41:38:@22228.4]
  wire  _T_61071; // @[Switch.scala 41:52:@22230.4]
  wire  output_6_23; // @[Switch.scala 41:38:@22231.4]
  wire  _T_61074; // @[Switch.scala 41:52:@22233.4]
  wire  output_6_24; // @[Switch.scala 41:38:@22234.4]
  wire  _T_61077; // @[Switch.scala 41:52:@22236.4]
  wire  output_6_25; // @[Switch.scala 41:38:@22237.4]
  wire  _T_61080; // @[Switch.scala 41:52:@22239.4]
  wire  output_6_26; // @[Switch.scala 41:38:@22240.4]
  wire  _T_61083; // @[Switch.scala 41:52:@22242.4]
  wire  output_6_27; // @[Switch.scala 41:38:@22243.4]
  wire  _T_61086; // @[Switch.scala 41:52:@22245.4]
  wire  output_6_28; // @[Switch.scala 41:38:@22246.4]
  wire  _T_61089; // @[Switch.scala 41:52:@22248.4]
  wire  output_6_29; // @[Switch.scala 41:38:@22249.4]
  wire  _T_61092; // @[Switch.scala 41:52:@22251.4]
  wire  output_6_30; // @[Switch.scala 41:38:@22252.4]
  wire  _T_61095; // @[Switch.scala 41:52:@22254.4]
  wire  output_6_31; // @[Switch.scala 41:38:@22255.4]
  wire  _T_61098; // @[Switch.scala 41:52:@22257.4]
  wire  output_6_32; // @[Switch.scala 41:38:@22258.4]
  wire  _T_61101; // @[Switch.scala 41:52:@22260.4]
  wire  output_6_33; // @[Switch.scala 41:38:@22261.4]
  wire  _T_61104; // @[Switch.scala 41:52:@22263.4]
  wire  output_6_34; // @[Switch.scala 41:38:@22264.4]
  wire  _T_61107; // @[Switch.scala 41:52:@22266.4]
  wire  output_6_35; // @[Switch.scala 41:38:@22267.4]
  wire  _T_61110; // @[Switch.scala 41:52:@22269.4]
  wire  output_6_36; // @[Switch.scala 41:38:@22270.4]
  wire  _T_61113; // @[Switch.scala 41:52:@22272.4]
  wire  output_6_37; // @[Switch.scala 41:38:@22273.4]
  wire  _T_61116; // @[Switch.scala 41:52:@22275.4]
  wire  output_6_38; // @[Switch.scala 41:38:@22276.4]
  wire  _T_61119; // @[Switch.scala 41:52:@22278.4]
  wire  output_6_39; // @[Switch.scala 41:38:@22279.4]
  wire  _T_61122; // @[Switch.scala 41:52:@22281.4]
  wire  output_6_40; // @[Switch.scala 41:38:@22282.4]
  wire  _T_61125; // @[Switch.scala 41:52:@22284.4]
  wire  output_6_41; // @[Switch.scala 41:38:@22285.4]
  wire  _T_61128; // @[Switch.scala 41:52:@22287.4]
  wire  output_6_42; // @[Switch.scala 41:38:@22288.4]
  wire  _T_61131; // @[Switch.scala 41:52:@22290.4]
  wire  output_6_43; // @[Switch.scala 41:38:@22291.4]
  wire  _T_61134; // @[Switch.scala 41:52:@22293.4]
  wire  output_6_44; // @[Switch.scala 41:38:@22294.4]
  wire  _T_61137; // @[Switch.scala 41:52:@22296.4]
  wire  output_6_45; // @[Switch.scala 41:38:@22297.4]
  wire  _T_61140; // @[Switch.scala 41:52:@22299.4]
  wire  output_6_46; // @[Switch.scala 41:38:@22300.4]
  wire  _T_61143; // @[Switch.scala 41:52:@22302.4]
  wire  output_6_47; // @[Switch.scala 41:38:@22303.4]
  wire  _T_61146; // @[Switch.scala 41:52:@22305.4]
  wire  output_6_48; // @[Switch.scala 41:38:@22306.4]
  wire  _T_61149; // @[Switch.scala 41:52:@22308.4]
  wire  output_6_49; // @[Switch.scala 41:38:@22309.4]
  wire  _T_61152; // @[Switch.scala 41:52:@22311.4]
  wire  output_6_50; // @[Switch.scala 41:38:@22312.4]
  wire  _T_61155; // @[Switch.scala 41:52:@22314.4]
  wire  output_6_51; // @[Switch.scala 41:38:@22315.4]
  wire  _T_61158; // @[Switch.scala 41:52:@22317.4]
  wire  output_6_52; // @[Switch.scala 41:38:@22318.4]
  wire  _T_61161; // @[Switch.scala 41:52:@22320.4]
  wire  output_6_53; // @[Switch.scala 41:38:@22321.4]
  wire  _T_61164; // @[Switch.scala 41:52:@22323.4]
  wire  output_6_54; // @[Switch.scala 41:38:@22324.4]
  wire  _T_61167; // @[Switch.scala 41:52:@22326.4]
  wire  output_6_55; // @[Switch.scala 41:38:@22327.4]
  wire  _T_61170; // @[Switch.scala 41:52:@22329.4]
  wire  output_6_56; // @[Switch.scala 41:38:@22330.4]
  wire  _T_61173; // @[Switch.scala 41:52:@22332.4]
  wire  output_6_57; // @[Switch.scala 41:38:@22333.4]
  wire  _T_61176; // @[Switch.scala 41:52:@22335.4]
  wire  output_6_58; // @[Switch.scala 41:38:@22336.4]
  wire  _T_61179; // @[Switch.scala 41:52:@22338.4]
  wire  output_6_59; // @[Switch.scala 41:38:@22339.4]
  wire  _T_61182; // @[Switch.scala 41:52:@22341.4]
  wire  output_6_60; // @[Switch.scala 41:38:@22342.4]
  wire  _T_61185; // @[Switch.scala 41:52:@22344.4]
  wire  output_6_61; // @[Switch.scala 41:38:@22345.4]
  wire  _T_61188; // @[Switch.scala 41:52:@22347.4]
  wire  output_6_62; // @[Switch.scala 41:38:@22348.4]
  wire  _T_61191; // @[Switch.scala 41:52:@22350.4]
  wire  output_6_63; // @[Switch.scala 41:38:@22351.4]
  wire [7:0] _T_61199; // @[Switch.scala 43:31:@22359.4]
  wire [15:0] _T_61207; // @[Switch.scala 43:31:@22367.4]
  wire [7:0] _T_61214; // @[Switch.scala 43:31:@22374.4]
  wire [31:0] _T_61223; // @[Switch.scala 43:31:@22383.4]
  wire [7:0] _T_61230; // @[Switch.scala 43:31:@22390.4]
  wire [15:0] _T_61238; // @[Switch.scala 43:31:@22398.4]
  wire [7:0] _T_61245; // @[Switch.scala 43:31:@22405.4]
  wire [31:0] _T_61254; // @[Switch.scala 43:31:@22414.4]
  wire [63:0] _T_61255; // @[Switch.scala 43:31:@22415.4]
  wire  _T_61259; // @[Switch.scala 41:52:@22418.4]
  wire  output_7_0; // @[Switch.scala 41:38:@22419.4]
  wire  _T_61262; // @[Switch.scala 41:52:@22421.4]
  wire  output_7_1; // @[Switch.scala 41:38:@22422.4]
  wire  _T_61265; // @[Switch.scala 41:52:@22424.4]
  wire  output_7_2; // @[Switch.scala 41:38:@22425.4]
  wire  _T_61268; // @[Switch.scala 41:52:@22427.4]
  wire  output_7_3; // @[Switch.scala 41:38:@22428.4]
  wire  _T_61271; // @[Switch.scala 41:52:@22430.4]
  wire  output_7_4; // @[Switch.scala 41:38:@22431.4]
  wire  _T_61274; // @[Switch.scala 41:52:@22433.4]
  wire  output_7_5; // @[Switch.scala 41:38:@22434.4]
  wire  _T_61277; // @[Switch.scala 41:52:@22436.4]
  wire  output_7_6; // @[Switch.scala 41:38:@22437.4]
  wire  _T_61280; // @[Switch.scala 41:52:@22439.4]
  wire  output_7_7; // @[Switch.scala 41:38:@22440.4]
  wire  _T_61283; // @[Switch.scala 41:52:@22442.4]
  wire  output_7_8; // @[Switch.scala 41:38:@22443.4]
  wire  _T_61286; // @[Switch.scala 41:52:@22445.4]
  wire  output_7_9; // @[Switch.scala 41:38:@22446.4]
  wire  _T_61289; // @[Switch.scala 41:52:@22448.4]
  wire  output_7_10; // @[Switch.scala 41:38:@22449.4]
  wire  _T_61292; // @[Switch.scala 41:52:@22451.4]
  wire  output_7_11; // @[Switch.scala 41:38:@22452.4]
  wire  _T_61295; // @[Switch.scala 41:52:@22454.4]
  wire  output_7_12; // @[Switch.scala 41:38:@22455.4]
  wire  _T_61298; // @[Switch.scala 41:52:@22457.4]
  wire  output_7_13; // @[Switch.scala 41:38:@22458.4]
  wire  _T_61301; // @[Switch.scala 41:52:@22460.4]
  wire  output_7_14; // @[Switch.scala 41:38:@22461.4]
  wire  _T_61304; // @[Switch.scala 41:52:@22463.4]
  wire  output_7_15; // @[Switch.scala 41:38:@22464.4]
  wire  _T_61307; // @[Switch.scala 41:52:@22466.4]
  wire  output_7_16; // @[Switch.scala 41:38:@22467.4]
  wire  _T_61310; // @[Switch.scala 41:52:@22469.4]
  wire  output_7_17; // @[Switch.scala 41:38:@22470.4]
  wire  _T_61313; // @[Switch.scala 41:52:@22472.4]
  wire  output_7_18; // @[Switch.scala 41:38:@22473.4]
  wire  _T_61316; // @[Switch.scala 41:52:@22475.4]
  wire  output_7_19; // @[Switch.scala 41:38:@22476.4]
  wire  _T_61319; // @[Switch.scala 41:52:@22478.4]
  wire  output_7_20; // @[Switch.scala 41:38:@22479.4]
  wire  _T_61322; // @[Switch.scala 41:52:@22481.4]
  wire  output_7_21; // @[Switch.scala 41:38:@22482.4]
  wire  _T_61325; // @[Switch.scala 41:52:@22484.4]
  wire  output_7_22; // @[Switch.scala 41:38:@22485.4]
  wire  _T_61328; // @[Switch.scala 41:52:@22487.4]
  wire  output_7_23; // @[Switch.scala 41:38:@22488.4]
  wire  _T_61331; // @[Switch.scala 41:52:@22490.4]
  wire  output_7_24; // @[Switch.scala 41:38:@22491.4]
  wire  _T_61334; // @[Switch.scala 41:52:@22493.4]
  wire  output_7_25; // @[Switch.scala 41:38:@22494.4]
  wire  _T_61337; // @[Switch.scala 41:52:@22496.4]
  wire  output_7_26; // @[Switch.scala 41:38:@22497.4]
  wire  _T_61340; // @[Switch.scala 41:52:@22499.4]
  wire  output_7_27; // @[Switch.scala 41:38:@22500.4]
  wire  _T_61343; // @[Switch.scala 41:52:@22502.4]
  wire  output_7_28; // @[Switch.scala 41:38:@22503.4]
  wire  _T_61346; // @[Switch.scala 41:52:@22505.4]
  wire  output_7_29; // @[Switch.scala 41:38:@22506.4]
  wire  _T_61349; // @[Switch.scala 41:52:@22508.4]
  wire  output_7_30; // @[Switch.scala 41:38:@22509.4]
  wire  _T_61352; // @[Switch.scala 41:52:@22511.4]
  wire  output_7_31; // @[Switch.scala 41:38:@22512.4]
  wire  _T_61355; // @[Switch.scala 41:52:@22514.4]
  wire  output_7_32; // @[Switch.scala 41:38:@22515.4]
  wire  _T_61358; // @[Switch.scala 41:52:@22517.4]
  wire  output_7_33; // @[Switch.scala 41:38:@22518.4]
  wire  _T_61361; // @[Switch.scala 41:52:@22520.4]
  wire  output_7_34; // @[Switch.scala 41:38:@22521.4]
  wire  _T_61364; // @[Switch.scala 41:52:@22523.4]
  wire  output_7_35; // @[Switch.scala 41:38:@22524.4]
  wire  _T_61367; // @[Switch.scala 41:52:@22526.4]
  wire  output_7_36; // @[Switch.scala 41:38:@22527.4]
  wire  _T_61370; // @[Switch.scala 41:52:@22529.4]
  wire  output_7_37; // @[Switch.scala 41:38:@22530.4]
  wire  _T_61373; // @[Switch.scala 41:52:@22532.4]
  wire  output_7_38; // @[Switch.scala 41:38:@22533.4]
  wire  _T_61376; // @[Switch.scala 41:52:@22535.4]
  wire  output_7_39; // @[Switch.scala 41:38:@22536.4]
  wire  _T_61379; // @[Switch.scala 41:52:@22538.4]
  wire  output_7_40; // @[Switch.scala 41:38:@22539.4]
  wire  _T_61382; // @[Switch.scala 41:52:@22541.4]
  wire  output_7_41; // @[Switch.scala 41:38:@22542.4]
  wire  _T_61385; // @[Switch.scala 41:52:@22544.4]
  wire  output_7_42; // @[Switch.scala 41:38:@22545.4]
  wire  _T_61388; // @[Switch.scala 41:52:@22547.4]
  wire  output_7_43; // @[Switch.scala 41:38:@22548.4]
  wire  _T_61391; // @[Switch.scala 41:52:@22550.4]
  wire  output_7_44; // @[Switch.scala 41:38:@22551.4]
  wire  _T_61394; // @[Switch.scala 41:52:@22553.4]
  wire  output_7_45; // @[Switch.scala 41:38:@22554.4]
  wire  _T_61397; // @[Switch.scala 41:52:@22556.4]
  wire  output_7_46; // @[Switch.scala 41:38:@22557.4]
  wire  _T_61400; // @[Switch.scala 41:52:@22559.4]
  wire  output_7_47; // @[Switch.scala 41:38:@22560.4]
  wire  _T_61403; // @[Switch.scala 41:52:@22562.4]
  wire  output_7_48; // @[Switch.scala 41:38:@22563.4]
  wire  _T_61406; // @[Switch.scala 41:52:@22565.4]
  wire  output_7_49; // @[Switch.scala 41:38:@22566.4]
  wire  _T_61409; // @[Switch.scala 41:52:@22568.4]
  wire  output_7_50; // @[Switch.scala 41:38:@22569.4]
  wire  _T_61412; // @[Switch.scala 41:52:@22571.4]
  wire  output_7_51; // @[Switch.scala 41:38:@22572.4]
  wire  _T_61415; // @[Switch.scala 41:52:@22574.4]
  wire  output_7_52; // @[Switch.scala 41:38:@22575.4]
  wire  _T_61418; // @[Switch.scala 41:52:@22577.4]
  wire  output_7_53; // @[Switch.scala 41:38:@22578.4]
  wire  _T_61421; // @[Switch.scala 41:52:@22580.4]
  wire  output_7_54; // @[Switch.scala 41:38:@22581.4]
  wire  _T_61424; // @[Switch.scala 41:52:@22583.4]
  wire  output_7_55; // @[Switch.scala 41:38:@22584.4]
  wire  _T_61427; // @[Switch.scala 41:52:@22586.4]
  wire  output_7_56; // @[Switch.scala 41:38:@22587.4]
  wire  _T_61430; // @[Switch.scala 41:52:@22589.4]
  wire  output_7_57; // @[Switch.scala 41:38:@22590.4]
  wire  _T_61433; // @[Switch.scala 41:52:@22592.4]
  wire  output_7_58; // @[Switch.scala 41:38:@22593.4]
  wire  _T_61436; // @[Switch.scala 41:52:@22595.4]
  wire  output_7_59; // @[Switch.scala 41:38:@22596.4]
  wire  _T_61439; // @[Switch.scala 41:52:@22598.4]
  wire  output_7_60; // @[Switch.scala 41:38:@22599.4]
  wire  _T_61442; // @[Switch.scala 41:52:@22601.4]
  wire  output_7_61; // @[Switch.scala 41:38:@22602.4]
  wire  _T_61445; // @[Switch.scala 41:52:@22604.4]
  wire  output_7_62; // @[Switch.scala 41:38:@22605.4]
  wire  _T_61448; // @[Switch.scala 41:52:@22607.4]
  wire  output_7_63; // @[Switch.scala 41:38:@22608.4]
  wire [7:0] _T_61456; // @[Switch.scala 43:31:@22616.4]
  wire [15:0] _T_61464; // @[Switch.scala 43:31:@22624.4]
  wire [7:0] _T_61471; // @[Switch.scala 43:31:@22631.4]
  wire [31:0] _T_61480; // @[Switch.scala 43:31:@22640.4]
  wire [7:0] _T_61487; // @[Switch.scala 43:31:@22647.4]
  wire [15:0] _T_61495; // @[Switch.scala 43:31:@22655.4]
  wire [7:0] _T_61502; // @[Switch.scala 43:31:@22662.4]
  wire [31:0] _T_61511; // @[Switch.scala 43:31:@22671.4]
  wire [63:0] _T_61512; // @[Switch.scala 43:31:@22672.4]
  wire  _T_61516; // @[Switch.scala 41:52:@22675.4]
  wire  output_8_0; // @[Switch.scala 41:38:@22676.4]
  wire  _T_61519; // @[Switch.scala 41:52:@22678.4]
  wire  output_8_1; // @[Switch.scala 41:38:@22679.4]
  wire  _T_61522; // @[Switch.scala 41:52:@22681.4]
  wire  output_8_2; // @[Switch.scala 41:38:@22682.4]
  wire  _T_61525; // @[Switch.scala 41:52:@22684.4]
  wire  output_8_3; // @[Switch.scala 41:38:@22685.4]
  wire  _T_61528; // @[Switch.scala 41:52:@22687.4]
  wire  output_8_4; // @[Switch.scala 41:38:@22688.4]
  wire  _T_61531; // @[Switch.scala 41:52:@22690.4]
  wire  output_8_5; // @[Switch.scala 41:38:@22691.4]
  wire  _T_61534; // @[Switch.scala 41:52:@22693.4]
  wire  output_8_6; // @[Switch.scala 41:38:@22694.4]
  wire  _T_61537; // @[Switch.scala 41:52:@22696.4]
  wire  output_8_7; // @[Switch.scala 41:38:@22697.4]
  wire  _T_61540; // @[Switch.scala 41:52:@22699.4]
  wire  output_8_8; // @[Switch.scala 41:38:@22700.4]
  wire  _T_61543; // @[Switch.scala 41:52:@22702.4]
  wire  output_8_9; // @[Switch.scala 41:38:@22703.4]
  wire  _T_61546; // @[Switch.scala 41:52:@22705.4]
  wire  output_8_10; // @[Switch.scala 41:38:@22706.4]
  wire  _T_61549; // @[Switch.scala 41:52:@22708.4]
  wire  output_8_11; // @[Switch.scala 41:38:@22709.4]
  wire  _T_61552; // @[Switch.scala 41:52:@22711.4]
  wire  output_8_12; // @[Switch.scala 41:38:@22712.4]
  wire  _T_61555; // @[Switch.scala 41:52:@22714.4]
  wire  output_8_13; // @[Switch.scala 41:38:@22715.4]
  wire  _T_61558; // @[Switch.scala 41:52:@22717.4]
  wire  output_8_14; // @[Switch.scala 41:38:@22718.4]
  wire  _T_61561; // @[Switch.scala 41:52:@22720.4]
  wire  output_8_15; // @[Switch.scala 41:38:@22721.4]
  wire  _T_61564; // @[Switch.scala 41:52:@22723.4]
  wire  output_8_16; // @[Switch.scala 41:38:@22724.4]
  wire  _T_61567; // @[Switch.scala 41:52:@22726.4]
  wire  output_8_17; // @[Switch.scala 41:38:@22727.4]
  wire  _T_61570; // @[Switch.scala 41:52:@22729.4]
  wire  output_8_18; // @[Switch.scala 41:38:@22730.4]
  wire  _T_61573; // @[Switch.scala 41:52:@22732.4]
  wire  output_8_19; // @[Switch.scala 41:38:@22733.4]
  wire  _T_61576; // @[Switch.scala 41:52:@22735.4]
  wire  output_8_20; // @[Switch.scala 41:38:@22736.4]
  wire  _T_61579; // @[Switch.scala 41:52:@22738.4]
  wire  output_8_21; // @[Switch.scala 41:38:@22739.4]
  wire  _T_61582; // @[Switch.scala 41:52:@22741.4]
  wire  output_8_22; // @[Switch.scala 41:38:@22742.4]
  wire  _T_61585; // @[Switch.scala 41:52:@22744.4]
  wire  output_8_23; // @[Switch.scala 41:38:@22745.4]
  wire  _T_61588; // @[Switch.scala 41:52:@22747.4]
  wire  output_8_24; // @[Switch.scala 41:38:@22748.4]
  wire  _T_61591; // @[Switch.scala 41:52:@22750.4]
  wire  output_8_25; // @[Switch.scala 41:38:@22751.4]
  wire  _T_61594; // @[Switch.scala 41:52:@22753.4]
  wire  output_8_26; // @[Switch.scala 41:38:@22754.4]
  wire  _T_61597; // @[Switch.scala 41:52:@22756.4]
  wire  output_8_27; // @[Switch.scala 41:38:@22757.4]
  wire  _T_61600; // @[Switch.scala 41:52:@22759.4]
  wire  output_8_28; // @[Switch.scala 41:38:@22760.4]
  wire  _T_61603; // @[Switch.scala 41:52:@22762.4]
  wire  output_8_29; // @[Switch.scala 41:38:@22763.4]
  wire  _T_61606; // @[Switch.scala 41:52:@22765.4]
  wire  output_8_30; // @[Switch.scala 41:38:@22766.4]
  wire  _T_61609; // @[Switch.scala 41:52:@22768.4]
  wire  output_8_31; // @[Switch.scala 41:38:@22769.4]
  wire  _T_61612; // @[Switch.scala 41:52:@22771.4]
  wire  output_8_32; // @[Switch.scala 41:38:@22772.4]
  wire  _T_61615; // @[Switch.scala 41:52:@22774.4]
  wire  output_8_33; // @[Switch.scala 41:38:@22775.4]
  wire  _T_61618; // @[Switch.scala 41:52:@22777.4]
  wire  output_8_34; // @[Switch.scala 41:38:@22778.4]
  wire  _T_61621; // @[Switch.scala 41:52:@22780.4]
  wire  output_8_35; // @[Switch.scala 41:38:@22781.4]
  wire  _T_61624; // @[Switch.scala 41:52:@22783.4]
  wire  output_8_36; // @[Switch.scala 41:38:@22784.4]
  wire  _T_61627; // @[Switch.scala 41:52:@22786.4]
  wire  output_8_37; // @[Switch.scala 41:38:@22787.4]
  wire  _T_61630; // @[Switch.scala 41:52:@22789.4]
  wire  output_8_38; // @[Switch.scala 41:38:@22790.4]
  wire  _T_61633; // @[Switch.scala 41:52:@22792.4]
  wire  output_8_39; // @[Switch.scala 41:38:@22793.4]
  wire  _T_61636; // @[Switch.scala 41:52:@22795.4]
  wire  output_8_40; // @[Switch.scala 41:38:@22796.4]
  wire  _T_61639; // @[Switch.scala 41:52:@22798.4]
  wire  output_8_41; // @[Switch.scala 41:38:@22799.4]
  wire  _T_61642; // @[Switch.scala 41:52:@22801.4]
  wire  output_8_42; // @[Switch.scala 41:38:@22802.4]
  wire  _T_61645; // @[Switch.scala 41:52:@22804.4]
  wire  output_8_43; // @[Switch.scala 41:38:@22805.4]
  wire  _T_61648; // @[Switch.scala 41:52:@22807.4]
  wire  output_8_44; // @[Switch.scala 41:38:@22808.4]
  wire  _T_61651; // @[Switch.scala 41:52:@22810.4]
  wire  output_8_45; // @[Switch.scala 41:38:@22811.4]
  wire  _T_61654; // @[Switch.scala 41:52:@22813.4]
  wire  output_8_46; // @[Switch.scala 41:38:@22814.4]
  wire  _T_61657; // @[Switch.scala 41:52:@22816.4]
  wire  output_8_47; // @[Switch.scala 41:38:@22817.4]
  wire  _T_61660; // @[Switch.scala 41:52:@22819.4]
  wire  output_8_48; // @[Switch.scala 41:38:@22820.4]
  wire  _T_61663; // @[Switch.scala 41:52:@22822.4]
  wire  output_8_49; // @[Switch.scala 41:38:@22823.4]
  wire  _T_61666; // @[Switch.scala 41:52:@22825.4]
  wire  output_8_50; // @[Switch.scala 41:38:@22826.4]
  wire  _T_61669; // @[Switch.scala 41:52:@22828.4]
  wire  output_8_51; // @[Switch.scala 41:38:@22829.4]
  wire  _T_61672; // @[Switch.scala 41:52:@22831.4]
  wire  output_8_52; // @[Switch.scala 41:38:@22832.4]
  wire  _T_61675; // @[Switch.scala 41:52:@22834.4]
  wire  output_8_53; // @[Switch.scala 41:38:@22835.4]
  wire  _T_61678; // @[Switch.scala 41:52:@22837.4]
  wire  output_8_54; // @[Switch.scala 41:38:@22838.4]
  wire  _T_61681; // @[Switch.scala 41:52:@22840.4]
  wire  output_8_55; // @[Switch.scala 41:38:@22841.4]
  wire  _T_61684; // @[Switch.scala 41:52:@22843.4]
  wire  output_8_56; // @[Switch.scala 41:38:@22844.4]
  wire  _T_61687; // @[Switch.scala 41:52:@22846.4]
  wire  output_8_57; // @[Switch.scala 41:38:@22847.4]
  wire  _T_61690; // @[Switch.scala 41:52:@22849.4]
  wire  output_8_58; // @[Switch.scala 41:38:@22850.4]
  wire  _T_61693; // @[Switch.scala 41:52:@22852.4]
  wire  output_8_59; // @[Switch.scala 41:38:@22853.4]
  wire  _T_61696; // @[Switch.scala 41:52:@22855.4]
  wire  output_8_60; // @[Switch.scala 41:38:@22856.4]
  wire  _T_61699; // @[Switch.scala 41:52:@22858.4]
  wire  output_8_61; // @[Switch.scala 41:38:@22859.4]
  wire  _T_61702; // @[Switch.scala 41:52:@22861.4]
  wire  output_8_62; // @[Switch.scala 41:38:@22862.4]
  wire  _T_61705; // @[Switch.scala 41:52:@22864.4]
  wire  output_8_63; // @[Switch.scala 41:38:@22865.4]
  wire [7:0] _T_61713; // @[Switch.scala 43:31:@22873.4]
  wire [15:0] _T_61721; // @[Switch.scala 43:31:@22881.4]
  wire [7:0] _T_61728; // @[Switch.scala 43:31:@22888.4]
  wire [31:0] _T_61737; // @[Switch.scala 43:31:@22897.4]
  wire [7:0] _T_61744; // @[Switch.scala 43:31:@22904.4]
  wire [15:0] _T_61752; // @[Switch.scala 43:31:@22912.4]
  wire [7:0] _T_61759; // @[Switch.scala 43:31:@22919.4]
  wire [31:0] _T_61768; // @[Switch.scala 43:31:@22928.4]
  wire [63:0] _T_61769; // @[Switch.scala 43:31:@22929.4]
  wire  _T_61773; // @[Switch.scala 41:52:@22932.4]
  wire  output_9_0; // @[Switch.scala 41:38:@22933.4]
  wire  _T_61776; // @[Switch.scala 41:52:@22935.4]
  wire  output_9_1; // @[Switch.scala 41:38:@22936.4]
  wire  _T_61779; // @[Switch.scala 41:52:@22938.4]
  wire  output_9_2; // @[Switch.scala 41:38:@22939.4]
  wire  _T_61782; // @[Switch.scala 41:52:@22941.4]
  wire  output_9_3; // @[Switch.scala 41:38:@22942.4]
  wire  _T_61785; // @[Switch.scala 41:52:@22944.4]
  wire  output_9_4; // @[Switch.scala 41:38:@22945.4]
  wire  _T_61788; // @[Switch.scala 41:52:@22947.4]
  wire  output_9_5; // @[Switch.scala 41:38:@22948.4]
  wire  _T_61791; // @[Switch.scala 41:52:@22950.4]
  wire  output_9_6; // @[Switch.scala 41:38:@22951.4]
  wire  _T_61794; // @[Switch.scala 41:52:@22953.4]
  wire  output_9_7; // @[Switch.scala 41:38:@22954.4]
  wire  _T_61797; // @[Switch.scala 41:52:@22956.4]
  wire  output_9_8; // @[Switch.scala 41:38:@22957.4]
  wire  _T_61800; // @[Switch.scala 41:52:@22959.4]
  wire  output_9_9; // @[Switch.scala 41:38:@22960.4]
  wire  _T_61803; // @[Switch.scala 41:52:@22962.4]
  wire  output_9_10; // @[Switch.scala 41:38:@22963.4]
  wire  _T_61806; // @[Switch.scala 41:52:@22965.4]
  wire  output_9_11; // @[Switch.scala 41:38:@22966.4]
  wire  _T_61809; // @[Switch.scala 41:52:@22968.4]
  wire  output_9_12; // @[Switch.scala 41:38:@22969.4]
  wire  _T_61812; // @[Switch.scala 41:52:@22971.4]
  wire  output_9_13; // @[Switch.scala 41:38:@22972.4]
  wire  _T_61815; // @[Switch.scala 41:52:@22974.4]
  wire  output_9_14; // @[Switch.scala 41:38:@22975.4]
  wire  _T_61818; // @[Switch.scala 41:52:@22977.4]
  wire  output_9_15; // @[Switch.scala 41:38:@22978.4]
  wire  _T_61821; // @[Switch.scala 41:52:@22980.4]
  wire  output_9_16; // @[Switch.scala 41:38:@22981.4]
  wire  _T_61824; // @[Switch.scala 41:52:@22983.4]
  wire  output_9_17; // @[Switch.scala 41:38:@22984.4]
  wire  _T_61827; // @[Switch.scala 41:52:@22986.4]
  wire  output_9_18; // @[Switch.scala 41:38:@22987.4]
  wire  _T_61830; // @[Switch.scala 41:52:@22989.4]
  wire  output_9_19; // @[Switch.scala 41:38:@22990.4]
  wire  _T_61833; // @[Switch.scala 41:52:@22992.4]
  wire  output_9_20; // @[Switch.scala 41:38:@22993.4]
  wire  _T_61836; // @[Switch.scala 41:52:@22995.4]
  wire  output_9_21; // @[Switch.scala 41:38:@22996.4]
  wire  _T_61839; // @[Switch.scala 41:52:@22998.4]
  wire  output_9_22; // @[Switch.scala 41:38:@22999.4]
  wire  _T_61842; // @[Switch.scala 41:52:@23001.4]
  wire  output_9_23; // @[Switch.scala 41:38:@23002.4]
  wire  _T_61845; // @[Switch.scala 41:52:@23004.4]
  wire  output_9_24; // @[Switch.scala 41:38:@23005.4]
  wire  _T_61848; // @[Switch.scala 41:52:@23007.4]
  wire  output_9_25; // @[Switch.scala 41:38:@23008.4]
  wire  _T_61851; // @[Switch.scala 41:52:@23010.4]
  wire  output_9_26; // @[Switch.scala 41:38:@23011.4]
  wire  _T_61854; // @[Switch.scala 41:52:@23013.4]
  wire  output_9_27; // @[Switch.scala 41:38:@23014.4]
  wire  _T_61857; // @[Switch.scala 41:52:@23016.4]
  wire  output_9_28; // @[Switch.scala 41:38:@23017.4]
  wire  _T_61860; // @[Switch.scala 41:52:@23019.4]
  wire  output_9_29; // @[Switch.scala 41:38:@23020.4]
  wire  _T_61863; // @[Switch.scala 41:52:@23022.4]
  wire  output_9_30; // @[Switch.scala 41:38:@23023.4]
  wire  _T_61866; // @[Switch.scala 41:52:@23025.4]
  wire  output_9_31; // @[Switch.scala 41:38:@23026.4]
  wire  _T_61869; // @[Switch.scala 41:52:@23028.4]
  wire  output_9_32; // @[Switch.scala 41:38:@23029.4]
  wire  _T_61872; // @[Switch.scala 41:52:@23031.4]
  wire  output_9_33; // @[Switch.scala 41:38:@23032.4]
  wire  _T_61875; // @[Switch.scala 41:52:@23034.4]
  wire  output_9_34; // @[Switch.scala 41:38:@23035.4]
  wire  _T_61878; // @[Switch.scala 41:52:@23037.4]
  wire  output_9_35; // @[Switch.scala 41:38:@23038.4]
  wire  _T_61881; // @[Switch.scala 41:52:@23040.4]
  wire  output_9_36; // @[Switch.scala 41:38:@23041.4]
  wire  _T_61884; // @[Switch.scala 41:52:@23043.4]
  wire  output_9_37; // @[Switch.scala 41:38:@23044.4]
  wire  _T_61887; // @[Switch.scala 41:52:@23046.4]
  wire  output_9_38; // @[Switch.scala 41:38:@23047.4]
  wire  _T_61890; // @[Switch.scala 41:52:@23049.4]
  wire  output_9_39; // @[Switch.scala 41:38:@23050.4]
  wire  _T_61893; // @[Switch.scala 41:52:@23052.4]
  wire  output_9_40; // @[Switch.scala 41:38:@23053.4]
  wire  _T_61896; // @[Switch.scala 41:52:@23055.4]
  wire  output_9_41; // @[Switch.scala 41:38:@23056.4]
  wire  _T_61899; // @[Switch.scala 41:52:@23058.4]
  wire  output_9_42; // @[Switch.scala 41:38:@23059.4]
  wire  _T_61902; // @[Switch.scala 41:52:@23061.4]
  wire  output_9_43; // @[Switch.scala 41:38:@23062.4]
  wire  _T_61905; // @[Switch.scala 41:52:@23064.4]
  wire  output_9_44; // @[Switch.scala 41:38:@23065.4]
  wire  _T_61908; // @[Switch.scala 41:52:@23067.4]
  wire  output_9_45; // @[Switch.scala 41:38:@23068.4]
  wire  _T_61911; // @[Switch.scala 41:52:@23070.4]
  wire  output_9_46; // @[Switch.scala 41:38:@23071.4]
  wire  _T_61914; // @[Switch.scala 41:52:@23073.4]
  wire  output_9_47; // @[Switch.scala 41:38:@23074.4]
  wire  _T_61917; // @[Switch.scala 41:52:@23076.4]
  wire  output_9_48; // @[Switch.scala 41:38:@23077.4]
  wire  _T_61920; // @[Switch.scala 41:52:@23079.4]
  wire  output_9_49; // @[Switch.scala 41:38:@23080.4]
  wire  _T_61923; // @[Switch.scala 41:52:@23082.4]
  wire  output_9_50; // @[Switch.scala 41:38:@23083.4]
  wire  _T_61926; // @[Switch.scala 41:52:@23085.4]
  wire  output_9_51; // @[Switch.scala 41:38:@23086.4]
  wire  _T_61929; // @[Switch.scala 41:52:@23088.4]
  wire  output_9_52; // @[Switch.scala 41:38:@23089.4]
  wire  _T_61932; // @[Switch.scala 41:52:@23091.4]
  wire  output_9_53; // @[Switch.scala 41:38:@23092.4]
  wire  _T_61935; // @[Switch.scala 41:52:@23094.4]
  wire  output_9_54; // @[Switch.scala 41:38:@23095.4]
  wire  _T_61938; // @[Switch.scala 41:52:@23097.4]
  wire  output_9_55; // @[Switch.scala 41:38:@23098.4]
  wire  _T_61941; // @[Switch.scala 41:52:@23100.4]
  wire  output_9_56; // @[Switch.scala 41:38:@23101.4]
  wire  _T_61944; // @[Switch.scala 41:52:@23103.4]
  wire  output_9_57; // @[Switch.scala 41:38:@23104.4]
  wire  _T_61947; // @[Switch.scala 41:52:@23106.4]
  wire  output_9_58; // @[Switch.scala 41:38:@23107.4]
  wire  _T_61950; // @[Switch.scala 41:52:@23109.4]
  wire  output_9_59; // @[Switch.scala 41:38:@23110.4]
  wire  _T_61953; // @[Switch.scala 41:52:@23112.4]
  wire  output_9_60; // @[Switch.scala 41:38:@23113.4]
  wire  _T_61956; // @[Switch.scala 41:52:@23115.4]
  wire  output_9_61; // @[Switch.scala 41:38:@23116.4]
  wire  _T_61959; // @[Switch.scala 41:52:@23118.4]
  wire  output_9_62; // @[Switch.scala 41:38:@23119.4]
  wire  _T_61962; // @[Switch.scala 41:52:@23121.4]
  wire  output_9_63; // @[Switch.scala 41:38:@23122.4]
  wire [7:0] _T_61970; // @[Switch.scala 43:31:@23130.4]
  wire [15:0] _T_61978; // @[Switch.scala 43:31:@23138.4]
  wire [7:0] _T_61985; // @[Switch.scala 43:31:@23145.4]
  wire [31:0] _T_61994; // @[Switch.scala 43:31:@23154.4]
  wire [7:0] _T_62001; // @[Switch.scala 43:31:@23161.4]
  wire [15:0] _T_62009; // @[Switch.scala 43:31:@23169.4]
  wire [7:0] _T_62016; // @[Switch.scala 43:31:@23176.4]
  wire [31:0] _T_62025; // @[Switch.scala 43:31:@23185.4]
  wire [63:0] _T_62026; // @[Switch.scala 43:31:@23186.4]
  wire  _T_62030; // @[Switch.scala 41:52:@23189.4]
  wire  output_10_0; // @[Switch.scala 41:38:@23190.4]
  wire  _T_62033; // @[Switch.scala 41:52:@23192.4]
  wire  output_10_1; // @[Switch.scala 41:38:@23193.4]
  wire  _T_62036; // @[Switch.scala 41:52:@23195.4]
  wire  output_10_2; // @[Switch.scala 41:38:@23196.4]
  wire  _T_62039; // @[Switch.scala 41:52:@23198.4]
  wire  output_10_3; // @[Switch.scala 41:38:@23199.4]
  wire  _T_62042; // @[Switch.scala 41:52:@23201.4]
  wire  output_10_4; // @[Switch.scala 41:38:@23202.4]
  wire  _T_62045; // @[Switch.scala 41:52:@23204.4]
  wire  output_10_5; // @[Switch.scala 41:38:@23205.4]
  wire  _T_62048; // @[Switch.scala 41:52:@23207.4]
  wire  output_10_6; // @[Switch.scala 41:38:@23208.4]
  wire  _T_62051; // @[Switch.scala 41:52:@23210.4]
  wire  output_10_7; // @[Switch.scala 41:38:@23211.4]
  wire  _T_62054; // @[Switch.scala 41:52:@23213.4]
  wire  output_10_8; // @[Switch.scala 41:38:@23214.4]
  wire  _T_62057; // @[Switch.scala 41:52:@23216.4]
  wire  output_10_9; // @[Switch.scala 41:38:@23217.4]
  wire  _T_62060; // @[Switch.scala 41:52:@23219.4]
  wire  output_10_10; // @[Switch.scala 41:38:@23220.4]
  wire  _T_62063; // @[Switch.scala 41:52:@23222.4]
  wire  output_10_11; // @[Switch.scala 41:38:@23223.4]
  wire  _T_62066; // @[Switch.scala 41:52:@23225.4]
  wire  output_10_12; // @[Switch.scala 41:38:@23226.4]
  wire  _T_62069; // @[Switch.scala 41:52:@23228.4]
  wire  output_10_13; // @[Switch.scala 41:38:@23229.4]
  wire  _T_62072; // @[Switch.scala 41:52:@23231.4]
  wire  output_10_14; // @[Switch.scala 41:38:@23232.4]
  wire  _T_62075; // @[Switch.scala 41:52:@23234.4]
  wire  output_10_15; // @[Switch.scala 41:38:@23235.4]
  wire  _T_62078; // @[Switch.scala 41:52:@23237.4]
  wire  output_10_16; // @[Switch.scala 41:38:@23238.4]
  wire  _T_62081; // @[Switch.scala 41:52:@23240.4]
  wire  output_10_17; // @[Switch.scala 41:38:@23241.4]
  wire  _T_62084; // @[Switch.scala 41:52:@23243.4]
  wire  output_10_18; // @[Switch.scala 41:38:@23244.4]
  wire  _T_62087; // @[Switch.scala 41:52:@23246.4]
  wire  output_10_19; // @[Switch.scala 41:38:@23247.4]
  wire  _T_62090; // @[Switch.scala 41:52:@23249.4]
  wire  output_10_20; // @[Switch.scala 41:38:@23250.4]
  wire  _T_62093; // @[Switch.scala 41:52:@23252.4]
  wire  output_10_21; // @[Switch.scala 41:38:@23253.4]
  wire  _T_62096; // @[Switch.scala 41:52:@23255.4]
  wire  output_10_22; // @[Switch.scala 41:38:@23256.4]
  wire  _T_62099; // @[Switch.scala 41:52:@23258.4]
  wire  output_10_23; // @[Switch.scala 41:38:@23259.4]
  wire  _T_62102; // @[Switch.scala 41:52:@23261.4]
  wire  output_10_24; // @[Switch.scala 41:38:@23262.4]
  wire  _T_62105; // @[Switch.scala 41:52:@23264.4]
  wire  output_10_25; // @[Switch.scala 41:38:@23265.4]
  wire  _T_62108; // @[Switch.scala 41:52:@23267.4]
  wire  output_10_26; // @[Switch.scala 41:38:@23268.4]
  wire  _T_62111; // @[Switch.scala 41:52:@23270.4]
  wire  output_10_27; // @[Switch.scala 41:38:@23271.4]
  wire  _T_62114; // @[Switch.scala 41:52:@23273.4]
  wire  output_10_28; // @[Switch.scala 41:38:@23274.4]
  wire  _T_62117; // @[Switch.scala 41:52:@23276.4]
  wire  output_10_29; // @[Switch.scala 41:38:@23277.4]
  wire  _T_62120; // @[Switch.scala 41:52:@23279.4]
  wire  output_10_30; // @[Switch.scala 41:38:@23280.4]
  wire  _T_62123; // @[Switch.scala 41:52:@23282.4]
  wire  output_10_31; // @[Switch.scala 41:38:@23283.4]
  wire  _T_62126; // @[Switch.scala 41:52:@23285.4]
  wire  output_10_32; // @[Switch.scala 41:38:@23286.4]
  wire  _T_62129; // @[Switch.scala 41:52:@23288.4]
  wire  output_10_33; // @[Switch.scala 41:38:@23289.4]
  wire  _T_62132; // @[Switch.scala 41:52:@23291.4]
  wire  output_10_34; // @[Switch.scala 41:38:@23292.4]
  wire  _T_62135; // @[Switch.scala 41:52:@23294.4]
  wire  output_10_35; // @[Switch.scala 41:38:@23295.4]
  wire  _T_62138; // @[Switch.scala 41:52:@23297.4]
  wire  output_10_36; // @[Switch.scala 41:38:@23298.4]
  wire  _T_62141; // @[Switch.scala 41:52:@23300.4]
  wire  output_10_37; // @[Switch.scala 41:38:@23301.4]
  wire  _T_62144; // @[Switch.scala 41:52:@23303.4]
  wire  output_10_38; // @[Switch.scala 41:38:@23304.4]
  wire  _T_62147; // @[Switch.scala 41:52:@23306.4]
  wire  output_10_39; // @[Switch.scala 41:38:@23307.4]
  wire  _T_62150; // @[Switch.scala 41:52:@23309.4]
  wire  output_10_40; // @[Switch.scala 41:38:@23310.4]
  wire  _T_62153; // @[Switch.scala 41:52:@23312.4]
  wire  output_10_41; // @[Switch.scala 41:38:@23313.4]
  wire  _T_62156; // @[Switch.scala 41:52:@23315.4]
  wire  output_10_42; // @[Switch.scala 41:38:@23316.4]
  wire  _T_62159; // @[Switch.scala 41:52:@23318.4]
  wire  output_10_43; // @[Switch.scala 41:38:@23319.4]
  wire  _T_62162; // @[Switch.scala 41:52:@23321.4]
  wire  output_10_44; // @[Switch.scala 41:38:@23322.4]
  wire  _T_62165; // @[Switch.scala 41:52:@23324.4]
  wire  output_10_45; // @[Switch.scala 41:38:@23325.4]
  wire  _T_62168; // @[Switch.scala 41:52:@23327.4]
  wire  output_10_46; // @[Switch.scala 41:38:@23328.4]
  wire  _T_62171; // @[Switch.scala 41:52:@23330.4]
  wire  output_10_47; // @[Switch.scala 41:38:@23331.4]
  wire  _T_62174; // @[Switch.scala 41:52:@23333.4]
  wire  output_10_48; // @[Switch.scala 41:38:@23334.4]
  wire  _T_62177; // @[Switch.scala 41:52:@23336.4]
  wire  output_10_49; // @[Switch.scala 41:38:@23337.4]
  wire  _T_62180; // @[Switch.scala 41:52:@23339.4]
  wire  output_10_50; // @[Switch.scala 41:38:@23340.4]
  wire  _T_62183; // @[Switch.scala 41:52:@23342.4]
  wire  output_10_51; // @[Switch.scala 41:38:@23343.4]
  wire  _T_62186; // @[Switch.scala 41:52:@23345.4]
  wire  output_10_52; // @[Switch.scala 41:38:@23346.4]
  wire  _T_62189; // @[Switch.scala 41:52:@23348.4]
  wire  output_10_53; // @[Switch.scala 41:38:@23349.4]
  wire  _T_62192; // @[Switch.scala 41:52:@23351.4]
  wire  output_10_54; // @[Switch.scala 41:38:@23352.4]
  wire  _T_62195; // @[Switch.scala 41:52:@23354.4]
  wire  output_10_55; // @[Switch.scala 41:38:@23355.4]
  wire  _T_62198; // @[Switch.scala 41:52:@23357.4]
  wire  output_10_56; // @[Switch.scala 41:38:@23358.4]
  wire  _T_62201; // @[Switch.scala 41:52:@23360.4]
  wire  output_10_57; // @[Switch.scala 41:38:@23361.4]
  wire  _T_62204; // @[Switch.scala 41:52:@23363.4]
  wire  output_10_58; // @[Switch.scala 41:38:@23364.4]
  wire  _T_62207; // @[Switch.scala 41:52:@23366.4]
  wire  output_10_59; // @[Switch.scala 41:38:@23367.4]
  wire  _T_62210; // @[Switch.scala 41:52:@23369.4]
  wire  output_10_60; // @[Switch.scala 41:38:@23370.4]
  wire  _T_62213; // @[Switch.scala 41:52:@23372.4]
  wire  output_10_61; // @[Switch.scala 41:38:@23373.4]
  wire  _T_62216; // @[Switch.scala 41:52:@23375.4]
  wire  output_10_62; // @[Switch.scala 41:38:@23376.4]
  wire  _T_62219; // @[Switch.scala 41:52:@23378.4]
  wire  output_10_63; // @[Switch.scala 41:38:@23379.4]
  wire [7:0] _T_62227; // @[Switch.scala 43:31:@23387.4]
  wire [15:0] _T_62235; // @[Switch.scala 43:31:@23395.4]
  wire [7:0] _T_62242; // @[Switch.scala 43:31:@23402.4]
  wire [31:0] _T_62251; // @[Switch.scala 43:31:@23411.4]
  wire [7:0] _T_62258; // @[Switch.scala 43:31:@23418.4]
  wire [15:0] _T_62266; // @[Switch.scala 43:31:@23426.4]
  wire [7:0] _T_62273; // @[Switch.scala 43:31:@23433.4]
  wire [31:0] _T_62282; // @[Switch.scala 43:31:@23442.4]
  wire [63:0] _T_62283; // @[Switch.scala 43:31:@23443.4]
  wire  _T_62287; // @[Switch.scala 41:52:@23446.4]
  wire  output_11_0; // @[Switch.scala 41:38:@23447.4]
  wire  _T_62290; // @[Switch.scala 41:52:@23449.4]
  wire  output_11_1; // @[Switch.scala 41:38:@23450.4]
  wire  _T_62293; // @[Switch.scala 41:52:@23452.4]
  wire  output_11_2; // @[Switch.scala 41:38:@23453.4]
  wire  _T_62296; // @[Switch.scala 41:52:@23455.4]
  wire  output_11_3; // @[Switch.scala 41:38:@23456.4]
  wire  _T_62299; // @[Switch.scala 41:52:@23458.4]
  wire  output_11_4; // @[Switch.scala 41:38:@23459.4]
  wire  _T_62302; // @[Switch.scala 41:52:@23461.4]
  wire  output_11_5; // @[Switch.scala 41:38:@23462.4]
  wire  _T_62305; // @[Switch.scala 41:52:@23464.4]
  wire  output_11_6; // @[Switch.scala 41:38:@23465.4]
  wire  _T_62308; // @[Switch.scala 41:52:@23467.4]
  wire  output_11_7; // @[Switch.scala 41:38:@23468.4]
  wire  _T_62311; // @[Switch.scala 41:52:@23470.4]
  wire  output_11_8; // @[Switch.scala 41:38:@23471.4]
  wire  _T_62314; // @[Switch.scala 41:52:@23473.4]
  wire  output_11_9; // @[Switch.scala 41:38:@23474.4]
  wire  _T_62317; // @[Switch.scala 41:52:@23476.4]
  wire  output_11_10; // @[Switch.scala 41:38:@23477.4]
  wire  _T_62320; // @[Switch.scala 41:52:@23479.4]
  wire  output_11_11; // @[Switch.scala 41:38:@23480.4]
  wire  _T_62323; // @[Switch.scala 41:52:@23482.4]
  wire  output_11_12; // @[Switch.scala 41:38:@23483.4]
  wire  _T_62326; // @[Switch.scala 41:52:@23485.4]
  wire  output_11_13; // @[Switch.scala 41:38:@23486.4]
  wire  _T_62329; // @[Switch.scala 41:52:@23488.4]
  wire  output_11_14; // @[Switch.scala 41:38:@23489.4]
  wire  _T_62332; // @[Switch.scala 41:52:@23491.4]
  wire  output_11_15; // @[Switch.scala 41:38:@23492.4]
  wire  _T_62335; // @[Switch.scala 41:52:@23494.4]
  wire  output_11_16; // @[Switch.scala 41:38:@23495.4]
  wire  _T_62338; // @[Switch.scala 41:52:@23497.4]
  wire  output_11_17; // @[Switch.scala 41:38:@23498.4]
  wire  _T_62341; // @[Switch.scala 41:52:@23500.4]
  wire  output_11_18; // @[Switch.scala 41:38:@23501.4]
  wire  _T_62344; // @[Switch.scala 41:52:@23503.4]
  wire  output_11_19; // @[Switch.scala 41:38:@23504.4]
  wire  _T_62347; // @[Switch.scala 41:52:@23506.4]
  wire  output_11_20; // @[Switch.scala 41:38:@23507.4]
  wire  _T_62350; // @[Switch.scala 41:52:@23509.4]
  wire  output_11_21; // @[Switch.scala 41:38:@23510.4]
  wire  _T_62353; // @[Switch.scala 41:52:@23512.4]
  wire  output_11_22; // @[Switch.scala 41:38:@23513.4]
  wire  _T_62356; // @[Switch.scala 41:52:@23515.4]
  wire  output_11_23; // @[Switch.scala 41:38:@23516.4]
  wire  _T_62359; // @[Switch.scala 41:52:@23518.4]
  wire  output_11_24; // @[Switch.scala 41:38:@23519.4]
  wire  _T_62362; // @[Switch.scala 41:52:@23521.4]
  wire  output_11_25; // @[Switch.scala 41:38:@23522.4]
  wire  _T_62365; // @[Switch.scala 41:52:@23524.4]
  wire  output_11_26; // @[Switch.scala 41:38:@23525.4]
  wire  _T_62368; // @[Switch.scala 41:52:@23527.4]
  wire  output_11_27; // @[Switch.scala 41:38:@23528.4]
  wire  _T_62371; // @[Switch.scala 41:52:@23530.4]
  wire  output_11_28; // @[Switch.scala 41:38:@23531.4]
  wire  _T_62374; // @[Switch.scala 41:52:@23533.4]
  wire  output_11_29; // @[Switch.scala 41:38:@23534.4]
  wire  _T_62377; // @[Switch.scala 41:52:@23536.4]
  wire  output_11_30; // @[Switch.scala 41:38:@23537.4]
  wire  _T_62380; // @[Switch.scala 41:52:@23539.4]
  wire  output_11_31; // @[Switch.scala 41:38:@23540.4]
  wire  _T_62383; // @[Switch.scala 41:52:@23542.4]
  wire  output_11_32; // @[Switch.scala 41:38:@23543.4]
  wire  _T_62386; // @[Switch.scala 41:52:@23545.4]
  wire  output_11_33; // @[Switch.scala 41:38:@23546.4]
  wire  _T_62389; // @[Switch.scala 41:52:@23548.4]
  wire  output_11_34; // @[Switch.scala 41:38:@23549.4]
  wire  _T_62392; // @[Switch.scala 41:52:@23551.4]
  wire  output_11_35; // @[Switch.scala 41:38:@23552.4]
  wire  _T_62395; // @[Switch.scala 41:52:@23554.4]
  wire  output_11_36; // @[Switch.scala 41:38:@23555.4]
  wire  _T_62398; // @[Switch.scala 41:52:@23557.4]
  wire  output_11_37; // @[Switch.scala 41:38:@23558.4]
  wire  _T_62401; // @[Switch.scala 41:52:@23560.4]
  wire  output_11_38; // @[Switch.scala 41:38:@23561.4]
  wire  _T_62404; // @[Switch.scala 41:52:@23563.4]
  wire  output_11_39; // @[Switch.scala 41:38:@23564.4]
  wire  _T_62407; // @[Switch.scala 41:52:@23566.4]
  wire  output_11_40; // @[Switch.scala 41:38:@23567.4]
  wire  _T_62410; // @[Switch.scala 41:52:@23569.4]
  wire  output_11_41; // @[Switch.scala 41:38:@23570.4]
  wire  _T_62413; // @[Switch.scala 41:52:@23572.4]
  wire  output_11_42; // @[Switch.scala 41:38:@23573.4]
  wire  _T_62416; // @[Switch.scala 41:52:@23575.4]
  wire  output_11_43; // @[Switch.scala 41:38:@23576.4]
  wire  _T_62419; // @[Switch.scala 41:52:@23578.4]
  wire  output_11_44; // @[Switch.scala 41:38:@23579.4]
  wire  _T_62422; // @[Switch.scala 41:52:@23581.4]
  wire  output_11_45; // @[Switch.scala 41:38:@23582.4]
  wire  _T_62425; // @[Switch.scala 41:52:@23584.4]
  wire  output_11_46; // @[Switch.scala 41:38:@23585.4]
  wire  _T_62428; // @[Switch.scala 41:52:@23587.4]
  wire  output_11_47; // @[Switch.scala 41:38:@23588.4]
  wire  _T_62431; // @[Switch.scala 41:52:@23590.4]
  wire  output_11_48; // @[Switch.scala 41:38:@23591.4]
  wire  _T_62434; // @[Switch.scala 41:52:@23593.4]
  wire  output_11_49; // @[Switch.scala 41:38:@23594.4]
  wire  _T_62437; // @[Switch.scala 41:52:@23596.4]
  wire  output_11_50; // @[Switch.scala 41:38:@23597.4]
  wire  _T_62440; // @[Switch.scala 41:52:@23599.4]
  wire  output_11_51; // @[Switch.scala 41:38:@23600.4]
  wire  _T_62443; // @[Switch.scala 41:52:@23602.4]
  wire  output_11_52; // @[Switch.scala 41:38:@23603.4]
  wire  _T_62446; // @[Switch.scala 41:52:@23605.4]
  wire  output_11_53; // @[Switch.scala 41:38:@23606.4]
  wire  _T_62449; // @[Switch.scala 41:52:@23608.4]
  wire  output_11_54; // @[Switch.scala 41:38:@23609.4]
  wire  _T_62452; // @[Switch.scala 41:52:@23611.4]
  wire  output_11_55; // @[Switch.scala 41:38:@23612.4]
  wire  _T_62455; // @[Switch.scala 41:52:@23614.4]
  wire  output_11_56; // @[Switch.scala 41:38:@23615.4]
  wire  _T_62458; // @[Switch.scala 41:52:@23617.4]
  wire  output_11_57; // @[Switch.scala 41:38:@23618.4]
  wire  _T_62461; // @[Switch.scala 41:52:@23620.4]
  wire  output_11_58; // @[Switch.scala 41:38:@23621.4]
  wire  _T_62464; // @[Switch.scala 41:52:@23623.4]
  wire  output_11_59; // @[Switch.scala 41:38:@23624.4]
  wire  _T_62467; // @[Switch.scala 41:52:@23626.4]
  wire  output_11_60; // @[Switch.scala 41:38:@23627.4]
  wire  _T_62470; // @[Switch.scala 41:52:@23629.4]
  wire  output_11_61; // @[Switch.scala 41:38:@23630.4]
  wire  _T_62473; // @[Switch.scala 41:52:@23632.4]
  wire  output_11_62; // @[Switch.scala 41:38:@23633.4]
  wire  _T_62476; // @[Switch.scala 41:52:@23635.4]
  wire  output_11_63; // @[Switch.scala 41:38:@23636.4]
  wire [7:0] _T_62484; // @[Switch.scala 43:31:@23644.4]
  wire [15:0] _T_62492; // @[Switch.scala 43:31:@23652.4]
  wire [7:0] _T_62499; // @[Switch.scala 43:31:@23659.4]
  wire [31:0] _T_62508; // @[Switch.scala 43:31:@23668.4]
  wire [7:0] _T_62515; // @[Switch.scala 43:31:@23675.4]
  wire [15:0] _T_62523; // @[Switch.scala 43:31:@23683.4]
  wire [7:0] _T_62530; // @[Switch.scala 43:31:@23690.4]
  wire [31:0] _T_62539; // @[Switch.scala 43:31:@23699.4]
  wire [63:0] _T_62540; // @[Switch.scala 43:31:@23700.4]
  wire  _T_62544; // @[Switch.scala 41:52:@23703.4]
  wire  output_12_0; // @[Switch.scala 41:38:@23704.4]
  wire  _T_62547; // @[Switch.scala 41:52:@23706.4]
  wire  output_12_1; // @[Switch.scala 41:38:@23707.4]
  wire  _T_62550; // @[Switch.scala 41:52:@23709.4]
  wire  output_12_2; // @[Switch.scala 41:38:@23710.4]
  wire  _T_62553; // @[Switch.scala 41:52:@23712.4]
  wire  output_12_3; // @[Switch.scala 41:38:@23713.4]
  wire  _T_62556; // @[Switch.scala 41:52:@23715.4]
  wire  output_12_4; // @[Switch.scala 41:38:@23716.4]
  wire  _T_62559; // @[Switch.scala 41:52:@23718.4]
  wire  output_12_5; // @[Switch.scala 41:38:@23719.4]
  wire  _T_62562; // @[Switch.scala 41:52:@23721.4]
  wire  output_12_6; // @[Switch.scala 41:38:@23722.4]
  wire  _T_62565; // @[Switch.scala 41:52:@23724.4]
  wire  output_12_7; // @[Switch.scala 41:38:@23725.4]
  wire  _T_62568; // @[Switch.scala 41:52:@23727.4]
  wire  output_12_8; // @[Switch.scala 41:38:@23728.4]
  wire  _T_62571; // @[Switch.scala 41:52:@23730.4]
  wire  output_12_9; // @[Switch.scala 41:38:@23731.4]
  wire  _T_62574; // @[Switch.scala 41:52:@23733.4]
  wire  output_12_10; // @[Switch.scala 41:38:@23734.4]
  wire  _T_62577; // @[Switch.scala 41:52:@23736.4]
  wire  output_12_11; // @[Switch.scala 41:38:@23737.4]
  wire  _T_62580; // @[Switch.scala 41:52:@23739.4]
  wire  output_12_12; // @[Switch.scala 41:38:@23740.4]
  wire  _T_62583; // @[Switch.scala 41:52:@23742.4]
  wire  output_12_13; // @[Switch.scala 41:38:@23743.4]
  wire  _T_62586; // @[Switch.scala 41:52:@23745.4]
  wire  output_12_14; // @[Switch.scala 41:38:@23746.4]
  wire  _T_62589; // @[Switch.scala 41:52:@23748.4]
  wire  output_12_15; // @[Switch.scala 41:38:@23749.4]
  wire  _T_62592; // @[Switch.scala 41:52:@23751.4]
  wire  output_12_16; // @[Switch.scala 41:38:@23752.4]
  wire  _T_62595; // @[Switch.scala 41:52:@23754.4]
  wire  output_12_17; // @[Switch.scala 41:38:@23755.4]
  wire  _T_62598; // @[Switch.scala 41:52:@23757.4]
  wire  output_12_18; // @[Switch.scala 41:38:@23758.4]
  wire  _T_62601; // @[Switch.scala 41:52:@23760.4]
  wire  output_12_19; // @[Switch.scala 41:38:@23761.4]
  wire  _T_62604; // @[Switch.scala 41:52:@23763.4]
  wire  output_12_20; // @[Switch.scala 41:38:@23764.4]
  wire  _T_62607; // @[Switch.scala 41:52:@23766.4]
  wire  output_12_21; // @[Switch.scala 41:38:@23767.4]
  wire  _T_62610; // @[Switch.scala 41:52:@23769.4]
  wire  output_12_22; // @[Switch.scala 41:38:@23770.4]
  wire  _T_62613; // @[Switch.scala 41:52:@23772.4]
  wire  output_12_23; // @[Switch.scala 41:38:@23773.4]
  wire  _T_62616; // @[Switch.scala 41:52:@23775.4]
  wire  output_12_24; // @[Switch.scala 41:38:@23776.4]
  wire  _T_62619; // @[Switch.scala 41:52:@23778.4]
  wire  output_12_25; // @[Switch.scala 41:38:@23779.4]
  wire  _T_62622; // @[Switch.scala 41:52:@23781.4]
  wire  output_12_26; // @[Switch.scala 41:38:@23782.4]
  wire  _T_62625; // @[Switch.scala 41:52:@23784.4]
  wire  output_12_27; // @[Switch.scala 41:38:@23785.4]
  wire  _T_62628; // @[Switch.scala 41:52:@23787.4]
  wire  output_12_28; // @[Switch.scala 41:38:@23788.4]
  wire  _T_62631; // @[Switch.scala 41:52:@23790.4]
  wire  output_12_29; // @[Switch.scala 41:38:@23791.4]
  wire  _T_62634; // @[Switch.scala 41:52:@23793.4]
  wire  output_12_30; // @[Switch.scala 41:38:@23794.4]
  wire  _T_62637; // @[Switch.scala 41:52:@23796.4]
  wire  output_12_31; // @[Switch.scala 41:38:@23797.4]
  wire  _T_62640; // @[Switch.scala 41:52:@23799.4]
  wire  output_12_32; // @[Switch.scala 41:38:@23800.4]
  wire  _T_62643; // @[Switch.scala 41:52:@23802.4]
  wire  output_12_33; // @[Switch.scala 41:38:@23803.4]
  wire  _T_62646; // @[Switch.scala 41:52:@23805.4]
  wire  output_12_34; // @[Switch.scala 41:38:@23806.4]
  wire  _T_62649; // @[Switch.scala 41:52:@23808.4]
  wire  output_12_35; // @[Switch.scala 41:38:@23809.4]
  wire  _T_62652; // @[Switch.scala 41:52:@23811.4]
  wire  output_12_36; // @[Switch.scala 41:38:@23812.4]
  wire  _T_62655; // @[Switch.scala 41:52:@23814.4]
  wire  output_12_37; // @[Switch.scala 41:38:@23815.4]
  wire  _T_62658; // @[Switch.scala 41:52:@23817.4]
  wire  output_12_38; // @[Switch.scala 41:38:@23818.4]
  wire  _T_62661; // @[Switch.scala 41:52:@23820.4]
  wire  output_12_39; // @[Switch.scala 41:38:@23821.4]
  wire  _T_62664; // @[Switch.scala 41:52:@23823.4]
  wire  output_12_40; // @[Switch.scala 41:38:@23824.4]
  wire  _T_62667; // @[Switch.scala 41:52:@23826.4]
  wire  output_12_41; // @[Switch.scala 41:38:@23827.4]
  wire  _T_62670; // @[Switch.scala 41:52:@23829.4]
  wire  output_12_42; // @[Switch.scala 41:38:@23830.4]
  wire  _T_62673; // @[Switch.scala 41:52:@23832.4]
  wire  output_12_43; // @[Switch.scala 41:38:@23833.4]
  wire  _T_62676; // @[Switch.scala 41:52:@23835.4]
  wire  output_12_44; // @[Switch.scala 41:38:@23836.4]
  wire  _T_62679; // @[Switch.scala 41:52:@23838.4]
  wire  output_12_45; // @[Switch.scala 41:38:@23839.4]
  wire  _T_62682; // @[Switch.scala 41:52:@23841.4]
  wire  output_12_46; // @[Switch.scala 41:38:@23842.4]
  wire  _T_62685; // @[Switch.scala 41:52:@23844.4]
  wire  output_12_47; // @[Switch.scala 41:38:@23845.4]
  wire  _T_62688; // @[Switch.scala 41:52:@23847.4]
  wire  output_12_48; // @[Switch.scala 41:38:@23848.4]
  wire  _T_62691; // @[Switch.scala 41:52:@23850.4]
  wire  output_12_49; // @[Switch.scala 41:38:@23851.4]
  wire  _T_62694; // @[Switch.scala 41:52:@23853.4]
  wire  output_12_50; // @[Switch.scala 41:38:@23854.4]
  wire  _T_62697; // @[Switch.scala 41:52:@23856.4]
  wire  output_12_51; // @[Switch.scala 41:38:@23857.4]
  wire  _T_62700; // @[Switch.scala 41:52:@23859.4]
  wire  output_12_52; // @[Switch.scala 41:38:@23860.4]
  wire  _T_62703; // @[Switch.scala 41:52:@23862.4]
  wire  output_12_53; // @[Switch.scala 41:38:@23863.4]
  wire  _T_62706; // @[Switch.scala 41:52:@23865.4]
  wire  output_12_54; // @[Switch.scala 41:38:@23866.4]
  wire  _T_62709; // @[Switch.scala 41:52:@23868.4]
  wire  output_12_55; // @[Switch.scala 41:38:@23869.4]
  wire  _T_62712; // @[Switch.scala 41:52:@23871.4]
  wire  output_12_56; // @[Switch.scala 41:38:@23872.4]
  wire  _T_62715; // @[Switch.scala 41:52:@23874.4]
  wire  output_12_57; // @[Switch.scala 41:38:@23875.4]
  wire  _T_62718; // @[Switch.scala 41:52:@23877.4]
  wire  output_12_58; // @[Switch.scala 41:38:@23878.4]
  wire  _T_62721; // @[Switch.scala 41:52:@23880.4]
  wire  output_12_59; // @[Switch.scala 41:38:@23881.4]
  wire  _T_62724; // @[Switch.scala 41:52:@23883.4]
  wire  output_12_60; // @[Switch.scala 41:38:@23884.4]
  wire  _T_62727; // @[Switch.scala 41:52:@23886.4]
  wire  output_12_61; // @[Switch.scala 41:38:@23887.4]
  wire  _T_62730; // @[Switch.scala 41:52:@23889.4]
  wire  output_12_62; // @[Switch.scala 41:38:@23890.4]
  wire  _T_62733; // @[Switch.scala 41:52:@23892.4]
  wire  output_12_63; // @[Switch.scala 41:38:@23893.4]
  wire [7:0] _T_62741; // @[Switch.scala 43:31:@23901.4]
  wire [15:0] _T_62749; // @[Switch.scala 43:31:@23909.4]
  wire [7:0] _T_62756; // @[Switch.scala 43:31:@23916.4]
  wire [31:0] _T_62765; // @[Switch.scala 43:31:@23925.4]
  wire [7:0] _T_62772; // @[Switch.scala 43:31:@23932.4]
  wire [15:0] _T_62780; // @[Switch.scala 43:31:@23940.4]
  wire [7:0] _T_62787; // @[Switch.scala 43:31:@23947.4]
  wire [31:0] _T_62796; // @[Switch.scala 43:31:@23956.4]
  wire [63:0] _T_62797; // @[Switch.scala 43:31:@23957.4]
  wire  _T_62801; // @[Switch.scala 41:52:@23960.4]
  wire  output_13_0; // @[Switch.scala 41:38:@23961.4]
  wire  _T_62804; // @[Switch.scala 41:52:@23963.4]
  wire  output_13_1; // @[Switch.scala 41:38:@23964.4]
  wire  _T_62807; // @[Switch.scala 41:52:@23966.4]
  wire  output_13_2; // @[Switch.scala 41:38:@23967.4]
  wire  _T_62810; // @[Switch.scala 41:52:@23969.4]
  wire  output_13_3; // @[Switch.scala 41:38:@23970.4]
  wire  _T_62813; // @[Switch.scala 41:52:@23972.4]
  wire  output_13_4; // @[Switch.scala 41:38:@23973.4]
  wire  _T_62816; // @[Switch.scala 41:52:@23975.4]
  wire  output_13_5; // @[Switch.scala 41:38:@23976.4]
  wire  _T_62819; // @[Switch.scala 41:52:@23978.4]
  wire  output_13_6; // @[Switch.scala 41:38:@23979.4]
  wire  _T_62822; // @[Switch.scala 41:52:@23981.4]
  wire  output_13_7; // @[Switch.scala 41:38:@23982.4]
  wire  _T_62825; // @[Switch.scala 41:52:@23984.4]
  wire  output_13_8; // @[Switch.scala 41:38:@23985.4]
  wire  _T_62828; // @[Switch.scala 41:52:@23987.4]
  wire  output_13_9; // @[Switch.scala 41:38:@23988.4]
  wire  _T_62831; // @[Switch.scala 41:52:@23990.4]
  wire  output_13_10; // @[Switch.scala 41:38:@23991.4]
  wire  _T_62834; // @[Switch.scala 41:52:@23993.4]
  wire  output_13_11; // @[Switch.scala 41:38:@23994.4]
  wire  _T_62837; // @[Switch.scala 41:52:@23996.4]
  wire  output_13_12; // @[Switch.scala 41:38:@23997.4]
  wire  _T_62840; // @[Switch.scala 41:52:@23999.4]
  wire  output_13_13; // @[Switch.scala 41:38:@24000.4]
  wire  _T_62843; // @[Switch.scala 41:52:@24002.4]
  wire  output_13_14; // @[Switch.scala 41:38:@24003.4]
  wire  _T_62846; // @[Switch.scala 41:52:@24005.4]
  wire  output_13_15; // @[Switch.scala 41:38:@24006.4]
  wire  _T_62849; // @[Switch.scala 41:52:@24008.4]
  wire  output_13_16; // @[Switch.scala 41:38:@24009.4]
  wire  _T_62852; // @[Switch.scala 41:52:@24011.4]
  wire  output_13_17; // @[Switch.scala 41:38:@24012.4]
  wire  _T_62855; // @[Switch.scala 41:52:@24014.4]
  wire  output_13_18; // @[Switch.scala 41:38:@24015.4]
  wire  _T_62858; // @[Switch.scala 41:52:@24017.4]
  wire  output_13_19; // @[Switch.scala 41:38:@24018.4]
  wire  _T_62861; // @[Switch.scala 41:52:@24020.4]
  wire  output_13_20; // @[Switch.scala 41:38:@24021.4]
  wire  _T_62864; // @[Switch.scala 41:52:@24023.4]
  wire  output_13_21; // @[Switch.scala 41:38:@24024.4]
  wire  _T_62867; // @[Switch.scala 41:52:@24026.4]
  wire  output_13_22; // @[Switch.scala 41:38:@24027.4]
  wire  _T_62870; // @[Switch.scala 41:52:@24029.4]
  wire  output_13_23; // @[Switch.scala 41:38:@24030.4]
  wire  _T_62873; // @[Switch.scala 41:52:@24032.4]
  wire  output_13_24; // @[Switch.scala 41:38:@24033.4]
  wire  _T_62876; // @[Switch.scala 41:52:@24035.4]
  wire  output_13_25; // @[Switch.scala 41:38:@24036.4]
  wire  _T_62879; // @[Switch.scala 41:52:@24038.4]
  wire  output_13_26; // @[Switch.scala 41:38:@24039.4]
  wire  _T_62882; // @[Switch.scala 41:52:@24041.4]
  wire  output_13_27; // @[Switch.scala 41:38:@24042.4]
  wire  _T_62885; // @[Switch.scala 41:52:@24044.4]
  wire  output_13_28; // @[Switch.scala 41:38:@24045.4]
  wire  _T_62888; // @[Switch.scala 41:52:@24047.4]
  wire  output_13_29; // @[Switch.scala 41:38:@24048.4]
  wire  _T_62891; // @[Switch.scala 41:52:@24050.4]
  wire  output_13_30; // @[Switch.scala 41:38:@24051.4]
  wire  _T_62894; // @[Switch.scala 41:52:@24053.4]
  wire  output_13_31; // @[Switch.scala 41:38:@24054.4]
  wire  _T_62897; // @[Switch.scala 41:52:@24056.4]
  wire  output_13_32; // @[Switch.scala 41:38:@24057.4]
  wire  _T_62900; // @[Switch.scala 41:52:@24059.4]
  wire  output_13_33; // @[Switch.scala 41:38:@24060.4]
  wire  _T_62903; // @[Switch.scala 41:52:@24062.4]
  wire  output_13_34; // @[Switch.scala 41:38:@24063.4]
  wire  _T_62906; // @[Switch.scala 41:52:@24065.4]
  wire  output_13_35; // @[Switch.scala 41:38:@24066.4]
  wire  _T_62909; // @[Switch.scala 41:52:@24068.4]
  wire  output_13_36; // @[Switch.scala 41:38:@24069.4]
  wire  _T_62912; // @[Switch.scala 41:52:@24071.4]
  wire  output_13_37; // @[Switch.scala 41:38:@24072.4]
  wire  _T_62915; // @[Switch.scala 41:52:@24074.4]
  wire  output_13_38; // @[Switch.scala 41:38:@24075.4]
  wire  _T_62918; // @[Switch.scala 41:52:@24077.4]
  wire  output_13_39; // @[Switch.scala 41:38:@24078.4]
  wire  _T_62921; // @[Switch.scala 41:52:@24080.4]
  wire  output_13_40; // @[Switch.scala 41:38:@24081.4]
  wire  _T_62924; // @[Switch.scala 41:52:@24083.4]
  wire  output_13_41; // @[Switch.scala 41:38:@24084.4]
  wire  _T_62927; // @[Switch.scala 41:52:@24086.4]
  wire  output_13_42; // @[Switch.scala 41:38:@24087.4]
  wire  _T_62930; // @[Switch.scala 41:52:@24089.4]
  wire  output_13_43; // @[Switch.scala 41:38:@24090.4]
  wire  _T_62933; // @[Switch.scala 41:52:@24092.4]
  wire  output_13_44; // @[Switch.scala 41:38:@24093.4]
  wire  _T_62936; // @[Switch.scala 41:52:@24095.4]
  wire  output_13_45; // @[Switch.scala 41:38:@24096.4]
  wire  _T_62939; // @[Switch.scala 41:52:@24098.4]
  wire  output_13_46; // @[Switch.scala 41:38:@24099.4]
  wire  _T_62942; // @[Switch.scala 41:52:@24101.4]
  wire  output_13_47; // @[Switch.scala 41:38:@24102.4]
  wire  _T_62945; // @[Switch.scala 41:52:@24104.4]
  wire  output_13_48; // @[Switch.scala 41:38:@24105.4]
  wire  _T_62948; // @[Switch.scala 41:52:@24107.4]
  wire  output_13_49; // @[Switch.scala 41:38:@24108.4]
  wire  _T_62951; // @[Switch.scala 41:52:@24110.4]
  wire  output_13_50; // @[Switch.scala 41:38:@24111.4]
  wire  _T_62954; // @[Switch.scala 41:52:@24113.4]
  wire  output_13_51; // @[Switch.scala 41:38:@24114.4]
  wire  _T_62957; // @[Switch.scala 41:52:@24116.4]
  wire  output_13_52; // @[Switch.scala 41:38:@24117.4]
  wire  _T_62960; // @[Switch.scala 41:52:@24119.4]
  wire  output_13_53; // @[Switch.scala 41:38:@24120.4]
  wire  _T_62963; // @[Switch.scala 41:52:@24122.4]
  wire  output_13_54; // @[Switch.scala 41:38:@24123.4]
  wire  _T_62966; // @[Switch.scala 41:52:@24125.4]
  wire  output_13_55; // @[Switch.scala 41:38:@24126.4]
  wire  _T_62969; // @[Switch.scala 41:52:@24128.4]
  wire  output_13_56; // @[Switch.scala 41:38:@24129.4]
  wire  _T_62972; // @[Switch.scala 41:52:@24131.4]
  wire  output_13_57; // @[Switch.scala 41:38:@24132.4]
  wire  _T_62975; // @[Switch.scala 41:52:@24134.4]
  wire  output_13_58; // @[Switch.scala 41:38:@24135.4]
  wire  _T_62978; // @[Switch.scala 41:52:@24137.4]
  wire  output_13_59; // @[Switch.scala 41:38:@24138.4]
  wire  _T_62981; // @[Switch.scala 41:52:@24140.4]
  wire  output_13_60; // @[Switch.scala 41:38:@24141.4]
  wire  _T_62984; // @[Switch.scala 41:52:@24143.4]
  wire  output_13_61; // @[Switch.scala 41:38:@24144.4]
  wire  _T_62987; // @[Switch.scala 41:52:@24146.4]
  wire  output_13_62; // @[Switch.scala 41:38:@24147.4]
  wire  _T_62990; // @[Switch.scala 41:52:@24149.4]
  wire  output_13_63; // @[Switch.scala 41:38:@24150.4]
  wire [7:0] _T_62998; // @[Switch.scala 43:31:@24158.4]
  wire [15:0] _T_63006; // @[Switch.scala 43:31:@24166.4]
  wire [7:0] _T_63013; // @[Switch.scala 43:31:@24173.4]
  wire [31:0] _T_63022; // @[Switch.scala 43:31:@24182.4]
  wire [7:0] _T_63029; // @[Switch.scala 43:31:@24189.4]
  wire [15:0] _T_63037; // @[Switch.scala 43:31:@24197.4]
  wire [7:0] _T_63044; // @[Switch.scala 43:31:@24204.4]
  wire [31:0] _T_63053; // @[Switch.scala 43:31:@24213.4]
  wire [63:0] _T_63054; // @[Switch.scala 43:31:@24214.4]
  wire  _T_63058; // @[Switch.scala 41:52:@24217.4]
  wire  output_14_0; // @[Switch.scala 41:38:@24218.4]
  wire  _T_63061; // @[Switch.scala 41:52:@24220.4]
  wire  output_14_1; // @[Switch.scala 41:38:@24221.4]
  wire  _T_63064; // @[Switch.scala 41:52:@24223.4]
  wire  output_14_2; // @[Switch.scala 41:38:@24224.4]
  wire  _T_63067; // @[Switch.scala 41:52:@24226.4]
  wire  output_14_3; // @[Switch.scala 41:38:@24227.4]
  wire  _T_63070; // @[Switch.scala 41:52:@24229.4]
  wire  output_14_4; // @[Switch.scala 41:38:@24230.4]
  wire  _T_63073; // @[Switch.scala 41:52:@24232.4]
  wire  output_14_5; // @[Switch.scala 41:38:@24233.4]
  wire  _T_63076; // @[Switch.scala 41:52:@24235.4]
  wire  output_14_6; // @[Switch.scala 41:38:@24236.4]
  wire  _T_63079; // @[Switch.scala 41:52:@24238.4]
  wire  output_14_7; // @[Switch.scala 41:38:@24239.4]
  wire  _T_63082; // @[Switch.scala 41:52:@24241.4]
  wire  output_14_8; // @[Switch.scala 41:38:@24242.4]
  wire  _T_63085; // @[Switch.scala 41:52:@24244.4]
  wire  output_14_9; // @[Switch.scala 41:38:@24245.4]
  wire  _T_63088; // @[Switch.scala 41:52:@24247.4]
  wire  output_14_10; // @[Switch.scala 41:38:@24248.4]
  wire  _T_63091; // @[Switch.scala 41:52:@24250.4]
  wire  output_14_11; // @[Switch.scala 41:38:@24251.4]
  wire  _T_63094; // @[Switch.scala 41:52:@24253.4]
  wire  output_14_12; // @[Switch.scala 41:38:@24254.4]
  wire  _T_63097; // @[Switch.scala 41:52:@24256.4]
  wire  output_14_13; // @[Switch.scala 41:38:@24257.4]
  wire  _T_63100; // @[Switch.scala 41:52:@24259.4]
  wire  output_14_14; // @[Switch.scala 41:38:@24260.4]
  wire  _T_63103; // @[Switch.scala 41:52:@24262.4]
  wire  output_14_15; // @[Switch.scala 41:38:@24263.4]
  wire  _T_63106; // @[Switch.scala 41:52:@24265.4]
  wire  output_14_16; // @[Switch.scala 41:38:@24266.4]
  wire  _T_63109; // @[Switch.scala 41:52:@24268.4]
  wire  output_14_17; // @[Switch.scala 41:38:@24269.4]
  wire  _T_63112; // @[Switch.scala 41:52:@24271.4]
  wire  output_14_18; // @[Switch.scala 41:38:@24272.4]
  wire  _T_63115; // @[Switch.scala 41:52:@24274.4]
  wire  output_14_19; // @[Switch.scala 41:38:@24275.4]
  wire  _T_63118; // @[Switch.scala 41:52:@24277.4]
  wire  output_14_20; // @[Switch.scala 41:38:@24278.4]
  wire  _T_63121; // @[Switch.scala 41:52:@24280.4]
  wire  output_14_21; // @[Switch.scala 41:38:@24281.4]
  wire  _T_63124; // @[Switch.scala 41:52:@24283.4]
  wire  output_14_22; // @[Switch.scala 41:38:@24284.4]
  wire  _T_63127; // @[Switch.scala 41:52:@24286.4]
  wire  output_14_23; // @[Switch.scala 41:38:@24287.4]
  wire  _T_63130; // @[Switch.scala 41:52:@24289.4]
  wire  output_14_24; // @[Switch.scala 41:38:@24290.4]
  wire  _T_63133; // @[Switch.scala 41:52:@24292.4]
  wire  output_14_25; // @[Switch.scala 41:38:@24293.4]
  wire  _T_63136; // @[Switch.scala 41:52:@24295.4]
  wire  output_14_26; // @[Switch.scala 41:38:@24296.4]
  wire  _T_63139; // @[Switch.scala 41:52:@24298.4]
  wire  output_14_27; // @[Switch.scala 41:38:@24299.4]
  wire  _T_63142; // @[Switch.scala 41:52:@24301.4]
  wire  output_14_28; // @[Switch.scala 41:38:@24302.4]
  wire  _T_63145; // @[Switch.scala 41:52:@24304.4]
  wire  output_14_29; // @[Switch.scala 41:38:@24305.4]
  wire  _T_63148; // @[Switch.scala 41:52:@24307.4]
  wire  output_14_30; // @[Switch.scala 41:38:@24308.4]
  wire  _T_63151; // @[Switch.scala 41:52:@24310.4]
  wire  output_14_31; // @[Switch.scala 41:38:@24311.4]
  wire  _T_63154; // @[Switch.scala 41:52:@24313.4]
  wire  output_14_32; // @[Switch.scala 41:38:@24314.4]
  wire  _T_63157; // @[Switch.scala 41:52:@24316.4]
  wire  output_14_33; // @[Switch.scala 41:38:@24317.4]
  wire  _T_63160; // @[Switch.scala 41:52:@24319.4]
  wire  output_14_34; // @[Switch.scala 41:38:@24320.4]
  wire  _T_63163; // @[Switch.scala 41:52:@24322.4]
  wire  output_14_35; // @[Switch.scala 41:38:@24323.4]
  wire  _T_63166; // @[Switch.scala 41:52:@24325.4]
  wire  output_14_36; // @[Switch.scala 41:38:@24326.4]
  wire  _T_63169; // @[Switch.scala 41:52:@24328.4]
  wire  output_14_37; // @[Switch.scala 41:38:@24329.4]
  wire  _T_63172; // @[Switch.scala 41:52:@24331.4]
  wire  output_14_38; // @[Switch.scala 41:38:@24332.4]
  wire  _T_63175; // @[Switch.scala 41:52:@24334.4]
  wire  output_14_39; // @[Switch.scala 41:38:@24335.4]
  wire  _T_63178; // @[Switch.scala 41:52:@24337.4]
  wire  output_14_40; // @[Switch.scala 41:38:@24338.4]
  wire  _T_63181; // @[Switch.scala 41:52:@24340.4]
  wire  output_14_41; // @[Switch.scala 41:38:@24341.4]
  wire  _T_63184; // @[Switch.scala 41:52:@24343.4]
  wire  output_14_42; // @[Switch.scala 41:38:@24344.4]
  wire  _T_63187; // @[Switch.scala 41:52:@24346.4]
  wire  output_14_43; // @[Switch.scala 41:38:@24347.4]
  wire  _T_63190; // @[Switch.scala 41:52:@24349.4]
  wire  output_14_44; // @[Switch.scala 41:38:@24350.4]
  wire  _T_63193; // @[Switch.scala 41:52:@24352.4]
  wire  output_14_45; // @[Switch.scala 41:38:@24353.4]
  wire  _T_63196; // @[Switch.scala 41:52:@24355.4]
  wire  output_14_46; // @[Switch.scala 41:38:@24356.4]
  wire  _T_63199; // @[Switch.scala 41:52:@24358.4]
  wire  output_14_47; // @[Switch.scala 41:38:@24359.4]
  wire  _T_63202; // @[Switch.scala 41:52:@24361.4]
  wire  output_14_48; // @[Switch.scala 41:38:@24362.4]
  wire  _T_63205; // @[Switch.scala 41:52:@24364.4]
  wire  output_14_49; // @[Switch.scala 41:38:@24365.4]
  wire  _T_63208; // @[Switch.scala 41:52:@24367.4]
  wire  output_14_50; // @[Switch.scala 41:38:@24368.4]
  wire  _T_63211; // @[Switch.scala 41:52:@24370.4]
  wire  output_14_51; // @[Switch.scala 41:38:@24371.4]
  wire  _T_63214; // @[Switch.scala 41:52:@24373.4]
  wire  output_14_52; // @[Switch.scala 41:38:@24374.4]
  wire  _T_63217; // @[Switch.scala 41:52:@24376.4]
  wire  output_14_53; // @[Switch.scala 41:38:@24377.4]
  wire  _T_63220; // @[Switch.scala 41:52:@24379.4]
  wire  output_14_54; // @[Switch.scala 41:38:@24380.4]
  wire  _T_63223; // @[Switch.scala 41:52:@24382.4]
  wire  output_14_55; // @[Switch.scala 41:38:@24383.4]
  wire  _T_63226; // @[Switch.scala 41:52:@24385.4]
  wire  output_14_56; // @[Switch.scala 41:38:@24386.4]
  wire  _T_63229; // @[Switch.scala 41:52:@24388.4]
  wire  output_14_57; // @[Switch.scala 41:38:@24389.4]
  wire  _T_63232; // @[Switch.scala 41:52:@24391.4]
  wire  output_14_58; // @[Switch.scala 41:38:@24392.4]
  wire  _T_63235; // @[Switch.scala 41:52:@24394.4]
  wire  output_14_59; // @[Switch.scala 41:38:@24395.4]
  wire  _T_63238; // @[Switch.scala 41:52:@24397.4]
  wire  output_14_60; // @[Switch.scala 41:38:@24398.4]
  wire  _T_63241; // @[Switch.scala 41:52:@24400.4]
  wire  output_14_61; // @[Switch.scala 41:38:@24401.4]
  wire  _T_63244; // @[Switch.scala 41:52:@24403.4]
  wire  output_14_62; // @[Switch.scala 41:38:@24404.4]
  wire  _T_63247; // @[Switch.scala 41:52:@24406.4]
  wire  output_14_63; // @[Switch.scala 41:38:@24407.4]
  wire [7:0] _T_63255; // @[Switch.scala 43:31:@24415.4]
  wire [15:0] _T_63263; // @[Switch.scala 43:31:@24423.4]
  wire [7:0] _T_63270; // @[Switch.scala 43:31:@24430.4]
  wire [31:0] _T_63279; // @[Switch.scala 43:31:@24439.4]
  wire [7:0] _T_63286; // @[Switch.scala 43:31:@24446.4]
  wire [15:0] _T_63294; // @[Switch.scala 43:31:@24454.4]
  wire [7:0] _T_63301; // @[Switch.scala 43:31:@24461.4]
  wire [31:0] _T_63310; // @[Switch.scala 43:31:@24470.4]
  wire [63:0] _T_63311; // @[Switch.scala 43:31:@24471.4]
  wire  _T_63315; // @[Switch.scala 41:52:@24474.4]
  wire  output_15_0; // @[Switch.scala 41:38:@24475.4]
  wire  _T_63318; // @[Switch.scala 41:52:@24477.4]
  wire  output_15_1; // @[Switch.scala 41:38:@24478.4]
  wire  _T_63321; // @[Switch.scala 41:52:@24480.4]
  wire  output_15_2; // @[Switch.scala 41:38:@24481.4]
  wire  _T_63324; // @[Switch.scala 41:52:@24483.4]
  wire  output_15_3; // @[Switch.scala 41:38:@24484.4]
  wire  _T_63327; // @[Switch.scala 41:52:@24486.4]
  wire  output_15_4; // @[Switch.scala 41:38:@24487.4]
  wire  _T_63330; // @[Switch.scala 41:52:@24489.4]
  wire  output_15_5; // @[Switch.scala 41:38:@24490.4]
  wire  _T_63333; // @[Switch.scala 41:52:@24492.4]
  wire  output_15_6; // @[Switch.scala 41:38:@24493.4]
  wire  _T_63336; // @[Switch.scala 41:52:@24495.4]
  wire  output_15_7; // @[Switch.scala 41:38:@24496.4]
  wire  _T_63339; // @[Switch.scala 41:52:@24498.4]
  wire  output_15_8; // @[Switch.scala 41:38:@24499.4]
  wire  _T_63342; // @[Switch.scala 41:52:@24501.4]
  wire  output_15_9; // @[Switch.scala 41:38:@24502.4]
  wire  _T_63345; // @[Switch.scala 41:52:@24504.4]
  wire  output_15_10; // @[Switch.scala 41:38:@24505.4]
  wire  _T_63348; // @[Switch.scala 41:52:@24507.4]
  wire  output_15_11; // @[Switch.scala 41:38:@24508.4]
  wire  _T_63351; // @[Switch.scala 41:52:@24510.4]
  wire  output_15_12; // @[Switch.scala 41:38:@24511.4]
  wire  _T_63354; // @[Switch.scala 41:52:@24513.4]
  wire  output_15_13; // @[Switch.scala 41:38:@24514.4]
  wire  _T_63357; // @[Switch.scala 41:52:@24516.4]
  wire  output_15_14; // @[Switch.scala 41:38:@24517.4]
  wire  _T_63360; // @[Switch.scala 41:52:@24519.4]
  wire  output_15_15; // @[Switch.scala 41:38:@24520.4]
  wire  _T_63363; // @[Switch.scala 41:52:@24522.4]
  wire  output_15_16; // @[Switch.scala 41:38:@24523.4]
  wire  _T_63366; // @[Switch.scala 41:52:@24525.4]
  wire  output_15_17; // @[Switch.scala 41:38:@24526.4]
  wire  _T_63369; // @[Switch.scala 41:52:@24528.4]
  wire  output_15_18; // @[Switch.scala 41:38:@24529.4]
  wire  _T_63372; // @[Switch.scala 41:52:@24531.4]
  wire  output_15_19; // @[Switch.scala 41:38:@24532.4]
  wire  _T_63375; // @[Switch.scala 41:52:@24534.4]
  wire  output_15_20; // @[Switch.scala 41:38:@24535.4]
  wire  _T_63378; // @[Switch.scala 41:52:@24537.4]
  wire  output_15_21; // @[Switch.scala 41:38:@24538.4]
  wire  _T_63381; // @[Switch.scala 41:52:@24540.4]
  wire  output_15_22; // @[Switch.scala 41:38:@24541.4]
  wire  _T_63384; // @[Switch.scala 41:52:@24543.4]
  wire  output_15_23; // @[Switch.scala 41:38:@24544.4]
  wire  _T_63387; // @[Switch.scala 41:52:@24546.4]
  wire  output_15_24; // @[Switch.scala 41:38:@24547.4]
  wire  _T_63390; // @[Switch.scala 41:52:@24549.4]
  wire  output_15_25; // @[Switch.scala 41:38:@24550.4]
  wire  _T_63393; // @[Switch.scala 41:52:@24552.4]
  wire  output_15_26; // @[Switch.scala 41:38:@24553.4]
  wire  _T_63396; // @[Switch.scala 41:52:@24555.4]
  wire  output_15_27; // @[Switch.scala 41:38:@24556.4]
  wire  _T_63399; // @[Switch.scala 41:52:@24558.4]
  wire  output_15_28; // @[Switch.scala 41:38:@24559.4]
  wire  _T_63402; // @[Switch.scala 41:52:@24561.4]
  wire  output_15_29; // @[Switch.scala 41:38:@24562.4]
  wire  _T_63405; // @[Switch.scala 41:52:@24564.4]
  wire  output_15_30; // @[Switch.scala 41:38:@24565.4]
  wire  _T_63408; // @[Switch.scala 41:52:@24567.4]
  wire  output_15_31; // @[Switch.scala 41:38:@24568.4]
  wire  _T_63411; // @[Switch.scala 41:52:@24570.4]
  wire  output_15_32; // @[Switch.scala 41:38:@24571.4]
  wire  _T_63414; // @[Switch.scala 41:52:@24573.4]
  wire  output_15_33; // @[Switch.scala 41:38:@24574.4]
  wire  _T_63417; // @[Switch.scala 41:52:@24576.4]
  wire  output_15_34; // @[Switch.scala 41:38:@24577.4]
  wire  _T_63420; // @[Switch.scala 41:52:@24579.4]
  wire  output_15_35; // @[Switch.scala 41:38:@24580.4]
  wire  _T_63423; // @[Switch.scala 41:52:@24582.4]
  wire  output_15_36; // @[Switch.scala 41:38:@24583.4]
  wire  _T_63426; // @[Switch.scala 41:52:@24585.4]
  wire  output_15_37; // @[Switch.scala 41:38:@24586.4]
  wire  _T_63429; // @[Switch.scala 41:52:@24588.4]
  wire  output_15_38; // @[Switch.scala 41:38:@24589.4]
  wire  _T_63432; // @[Switch.scala 41:52:@24591.4]
  wire  output_15_39; // @[Switch.scala 41:38:@24592.4]
  wire  _T_63435; // @[Switch.scala 41:52:@24594.4]
  wire  output_15_40; // @[Switch.scala 41:38:@24595.4]
  wire  _T_63438; // @[Switch.scala 41:52:@24597.4]
  wire  output_15_41; // @[Switch.scala 41:38:@24598.4]
  wire  _T_63441; // @[Switch.scala 41:52:@24600.4]
  wire  output_15_42; // @[Switch.scala 41:38:@24601.4]
  wire  _T_63444; // @[Switch.scala 41:52:@24603.4]
  wire  output_15_43; // @[Switch.scala 41:38:@24604.4]
  wire  _T_63447; // @[Switch.scala 41:52:@24606.4]
  wire  output_15_44; // @[Switch.scala 41:38:@24607.4]
  wire  _T_63450; // @[Switch.scala 41:52:@24609.4]
  wire  output_15_45; // @[Switch.scala 41:38:@24610.4]
  wire  _T_63453; // @[Switch.scala 41:52:@24612.4]
  wire  output_15_46; // @[Switch.scala 41:38:@24613.4]
  wire  _T_63456; // @[Switch.scala 41:52:@24615.4]
  wire  output_15_47; // @[Switch.scala 41:38:@24616.4]
  wire  _T_63459; // @[Switch.scala 41:52:@24618.4]
  wire  output_15_48; // @[Switch.scala 41:38:@24619.4]
  wire  _T_63462; // @[Switch.scala 41:52:@24621.4]
  wire  output_15_49; // @[Switch.scala 41:38:@24622.4]
  wire  _T_63465; // @[Switch.scala 41:52:@24624.4]
  wire  output_15_50; // @[Switch.scala 41:38:@24625.4]
  wire  _T_63468; // @[Switch.scala 41:52:@24627.4]
  wire  output_15_51; // @[Switch.scala 41:38:@24628.4]
  wire  _T_63471; // @[Switch.scala 41:52:@24630.4]
  wire  output_15_52; // @[Switch.scala 41:38:@24631.4]
  wire  _T_63474; // @[Switch.scala 41:52:@24633.4]
  wire  output_15_53; // @[Switch.scala 41:38:@24634.4]
  wire  _T_63477; // @[Switch.scala 41:52:@24636.4]
  wire  output_15_54; // @[Switch.scala 41:38:@24637.4]
  wire  _T_63480; // @[Switch.scala 41:52:@24639.4]
  wire  output_15_55; // @[Switch.scala 41:38:@24640.4]
  wire  _T_63483; // @[Switch.scala 41:52:@24642.4]
  wire  output_15_56; // @[Switch.scala 41:38:@24643.4]
  wire  _T_63486; // @[Switch.scala 41:52:@24645.4]
  wire  output_15_57; // @[Switch.scala 41:38:@24646.4]
  wire  _T_63489; // @[Switch.scala 41:52:@24648.4]
  wire  output_15_58; // @[Switch.scala 41:38:@24649.4]
  wire  _T_63492; // @[Switch.scala 41:52:@24651.4]
  wire  output_15_59; // @[Switch.scala 41:38:@24652.4]
  wire  _T_63495; // @[Switch.scala 41:52:@24654.4]
  wire  output_15_60; // @[Switch.scala 41:38:@24655.4]
  wire  _T_63498; // @[Switch.scala 41:52:@24657.4]
  wire  output_15_61; // @[Switch.scala 41:38:@24658.4]
  wire  _T_63501; // @[Switch.scala 41:52:@24660.4]
  wire  output_15_62; // @[Switch.scala 41:38:@24661.4]
  wire  _T_63504; // @[Switch.scala 41:52:@24663.4]
  wire  output_15_63; // @[Switch.scala 41:38:@24664.4]
  wire [7:0] _T_63512; // @[Switch.scala 43:31:@24672.4]
  wire [15:0] _T_63520; // @[Switch.scala 43:31:@24680.4]
  wire [7:0] _T_63527; // @[Switch.scala 43:31:@24687.4]
  wire [31:0] _T_63536; // @[Switch.scala 43:31:@24696.4]
  wire [7:0] _T_63543; // @[Switch.scala 43:31:@24703.4]
  wire [15:0] _T_63551; // @[Switch.scala 43:31:@24711.4]
  wire [7:0] _T_63558; // @[Switch.scala 43:31:@24718.4]
  wire [31:0] _T_63567; // @[Switch.scala 43:31:@24727.4]
  wire [63:0] _T_63568; // @[Switch.scala 43:31:@24728.4]
  wire  _T_63572; // @[Switch.scala 41:52:@24731.4]
  wire  output_16_0; // @[Switch.scala 41:38:@24732.4]
  wire  _T_63575; // @[Switch.scala 41:52:@24734.4]
  wire  output_16_1; // @[Switch.scala 41:38:@24735.4]
  wire  _T_63578; // @[Switch.scala 41:52:@24737.4]
  wire  output_16_2; // @[Switch.scala 41:38:@24738.4]
  wire  _T_63581; // @[Switch.scala 41:52:@24740.4]
  wire  output_16_3; // @[Switch.scala 41:38:@24741.4]
  wire  _T_63584; // @[Switch.scala 41:52:@24743.4]
  wire  output_16_4; // @[Switch.scala 41:38:@24744.4]
  wire  _T_63587; // @[Switch.scala 41:52:@24746.4]
  wire  output_16_5; // @[Switch.scala 41:38:@24747.4]
  wire  _T_63590; // @[Switch.scala 41:52:@24749.4]
  wire  output_16_6; // @[Switch.scala 41:38:@24750.4]
  wire  _T_63593; // @[Switch.scala 41:52:@24752.4]
  wire  output_16_7; // @[Switch.scala 41:38:@24753.4]
  wire  _T_63596; // @[Switch.scala 41:52:@24755.4]
  wire  output_16_8; // @[Switch.scala 41:38:@24756.4]
  wire  _T_63599; // @[Switch.scala 41:52:@24758.4]
  wire  output_16_9; // @[Switch.scala 41:38:@24759.4]
  wire  _T_63602; // @[Switch.scala 41:52:@24761.4]
  wire  output_16_10; // @[Switch.scala 41:38:@24762.4]
  wire  _T_63605; // @[Switch.scala 41:52:@24764.4]
  wire  output_16_11; // @[Switch.scala 41:38:@24765.4]
  wire  _T_63608; // @[Switch.scala 41:52:@24767.4]
  wire  output_16_12; // @[Switch.scala 41:38:@24768.4]
  wire  _T_63611; // @[Switch.scala 41:52:@24770.4]
  wire  output_16_13; // @[Switch.scala 41:38:@24771.4]
  wire  _T_63614; // @[Switch.scala 41:52:@24773.4]
  wire  output_16_14; // @[Switch.scala 41:38:@24774.4]
  wire  _T_63617; // @[Switch.scala 41:52:@24776.4]
  wire  output_16_15; // @[Switch.scala 41:38:@24777.4]
  wire  _T_63620; // @[Switch.scala 41:52:@24779.4]
  wire  output_16_16; // @[Switch.scala 41:38:@24780.4]
  wire  _T_63623; // @[Switch.scala 41:52:@24782.4]
  wire  output_16_17; // @[Switch.scala 41:38:@24783.4]
  wire  _T_63626; // @[Switch.scala 41:52:@24785.4]
  wire  output_16_18; // @[Switch.scala 41:38:@24786.4]
  wire  _T_63629; // @[Switch.scala 41:52:@24788.4]
  wire  output_16_19; // @[Switch.scala 41:38:@24789.4]
  wire  _T_63632; // @[Switch.scala 41:52:@24791.4]
  wire  output_16_20; // @[Switch.scala 41:38:@24792.4]
  wire  _T_63635; // @[Switch.scala 41:52:@24794.4]
  wire  output_16_21; // @[Switch.scala 41:38:@24795.4]
  wire  _T_63638; // @[Switch.scala 41:52:@24797.4]
  wire  output_16_22; // @[Switch.scala 41:38:@24798.4]
  wire  _T_63641; // @[Switch.scala 41:52:@24800.4]
  wire  output_16_23; // @[Switch.scala 41:38:@24801.4]
  wire  _T_63644; // @[Switch.scala 41:52:@24803.4]
  wire  output_16_24; // @[Switch.scala 41:38:@24804.4]
  wire  _T_63647; // @[Switch.scala 41:52:@24806.4]
  wire  output_16_25; // @[Switch.scala 41:38:@24807.4]
  wire  _T_63650; // @[Switch.scala 41:52:@24809.4]
  wire  output_16_26; // @[Switch.scala 41:38:@24810.4]
  wire  _T_63653; // @[Switch.scala 41:52:@24812.4]
  wire  output_16_27; // @[Switch.scala 41:38:@24813.4]
  wire  _T_63656; // @[Switch.scala 41:52:@24815.4]
  wire  output_16_28; // @[Switch.scala 41:38:@24816.4]
  wire  _T_63659; // @[Switch.scala 41:52:@24818.4]
  wire  output_16_29; // @[Switch.scala 41:38:@24819.4]
  wire  _T_63662; // @[Switch.scala 41:52:@24821.4]
  wire  output_16_30; // @[Switch.scala 41:38:@24822.4]
  wire  _T_63665; // @[Switch.scala 41:52:@24824.4]
  wire  output_16_31; // @[Switch.scala 41:38:@24825.4]
  wire  _T_63668; // @[Switch.scala 41:52:@24827.4]
  wire  output_16_32; // @[Switch.scala 41:38:@24828.4]
  wire  _T_63671; // @[Switch.scala 41:52:@24830.4]
  wire  output_16_33; // @[Switch.scala 41:38:@24831.4]
  wire  _T_63674; // @[Switch.scala 41:52:@24833.4]
  wire  output_16_34; // @[Switch.scala 41:38:@24834.4]
  wire  _T_63677; // @[Switch.scala 41:52:@24836.4]
  wire  output_16_35; // @[Switch.scala 41:38:@24837.4]
  wire  _T_63680; // @[Switch.scala 41:52:@24839.4]
  wire  output_16_36; // @[Switch.scala 41:38:@24840.4]
  wire  _T_63683; // @[Switch.scala 41:52:@24842.4]
  wire  output_16_37; // @[Switch.scala 41:38:@24843.4]
  wire  _T_63686; // @[Switch.scala 41:52:@24845.4]
  wire  output_16_38; // @[Switch.scala 41:38:@24846.4]
  wire  _T_63689; // @[Switch.scala 41:52:@24848.4]
  wire  output_16_39; // @[Switch.scala 41:38:@24849.4]
  wire  _T_63692; // @[Switch.scala 41:52:@24851.4]
  wire  output_16_40; // @[Switch.scala 41:38:@24852.4]
  wire  _T_63695; // @[Switch.scala 41:52:@24854.4]
  wire  output_16_41; // @[Switch.scala 41:38:@24855.4]
  wire  _T_63698; // @[Switch.scala 41:52:@24857.4]
  wire  output_16_42; // @[Switch.scala 41:38:@24858.4]
  wire  _T_63701; // @[Switch.scala 41:52:@24860.4]
  wire  output_16_43; // @[Switch.scala 41:38:@24861.4]
  wire  _T_63704; // @[Switch.scala 41:52:@24863.4]
  wire  output_16_44; // @[Switch.scala 41:38:@24864.4]
  wire  _T_63707; // @[Switch.scala 41:52:@24866.4]
  wire  output_16_45; // @[Switch.scala 41:38:@24867.4]
  wire  _T_63710; // @[Switch.scala 41:52:@24869.4]
  wire  output_16_46; // @[Switch.scala 41:38:@24870.4]
  wire  _T_63713; // @[Switch.scala 41:52:@24872.4]
  wire  output_16_47; // @[Switch.scala 41:38:@24873.4]
  wire  _T_63716; // @[Switch.scala 41:52:@24875.4]
  wire  output_16_48; // @[Switch.scala 41:38:@24876.4]
  wire  _T_63719; // @[Switch.scala 41:52:@24878.4]
  wire  output_16_49; // @[Switch.scala 41:38:@24879.4]
  wire  _T_63722; // @[Switch.scala 41:52:@24881.4]
  wire  output_16_50; // @[Switch.scala 41:38:@24882.4]
  wire  _T_63725; // @[Switch.scala 41:52:@24884.4]
  wire  output_16_51; // @[Switch.scala 41:38:@24885.4]
  wire  _T_63728; // @[Switch.scala 41:52:@24887.4]
  wire  output_16_52; // @[Switch.scala 41:38:@24888.4]
  wire  _T_63731; // @[Switch.scala 41:52:@24890.4]
  wire  output_16_53; // @[Switch.scala 41:38:@24891.4]
  wire  _T_63734; // @[Switch.scala 41:52:@24893.4]
  wire  output_16_54; // @[Switch.scala 41:38:@24894.4]
  wire  _T_63737; // @[Switch.scala 41:52:@24896.4]
  wire  output_16_55; // @[Switch.scala 41:38:@24897.4]
  wire  _T_63740; // @[Switch.scala 41:52:@24899.4]
  wire  output_16_56; // @[Switch.scala 41:38:@24900.4]
  wire  _T_63743; // @[Switch.scala 41:52:@24902.4]
  wire  output_16_57; // @[Switch.scala 41:38:@24903.4]
  wire  _T_63746; // @[Switch.scala 41:52:@24905.4]
  wire  output_16_58; // @[Switch.scala 41:38:@24906.4]
  wire  _T_63749; // @[Switch.scala 41:52:@24908.4]
  wire  output_16_59; // @[Switch.scala 41:38:@24909.4]
  wire  _T_63752; // @[Switch.scala 41:52:@24911.4]
  wire  output_16_60; // @[Switch.scala 41:38:@24912.4]
  wire  _T_63755; // @[Switch.scala 41:52:@24914.4]
  wire  output_16_61; // @[Switch.scala 41:38:@24915.4]
  wire  _T_63758; // @[Switch.scala 41:52:@24917.4]
  wire  output_16_62; // @[Switch.scala 41:38:@24918.4]
  wire  _T_63761; // @[Switch.scala 41:52:@24920.4]
  wire  output_16_63; // @[Switch.scala 41:38:@24921.4]
  wire [7:0] _T_63769; // @[Switch.scala 43:31:@24929.4]
  wire [15:0] _T_63777; // @[Switch.scala 43:31:@24937.4]
  wire [7:0] _T_63784; // @[Switch.scala 43:31:@24944.4]
  wire [31:0] _T_63793; // @[Switch.scala 43:31:@24953.4]
  wire [7:0] _T_63800; // @[Switch.scala 43:31:@24960.4]
  wire [15:0] _T_63808; // @[Switch.scala 43:31:@24968.4]
  wire [7:0] _T_63815; // @[Switch.scala 43:31:@24975.4]
  wire [31:0] _T_63824; // @[Switch.scala 43:31:@24984.4]
  wire [63:0] _T_63825; // @[Switch.scala 43:31:@24985.4]
  wire  _T_63829; // @[Switch.scala 41:52:@24988.4]
  wire  output_17_0; // @[Switch.scala 41:38:@24989.4]
  wire  _T_63832; // @[Switch.scala 41:52:@24991.4]
  wire  output_17_1; // @[Switch.scala 41:38:@24992.4]
  wire  _T_63835; // @[Switch.scala 41:52:@24994.4]
  wire  output_17_2; // @[Switch.scala 41:38:@24995.4]
  wire  _T_63838; // @[Switch.scala 41:52:@24997.4]
  wire  output_17_3; // @[Switch.scala 41:38:@24998.4]
  wire  _T_63841; // @[Switch.scala 41:52:@25000.4]
  wire  output_17_4; // @[Switch.scala 41:38:@25001.4]
  wire  _T_63844; // @[Switch.scala 41:52:@25003.4]
  wire  output_17_5; // @[Switch.scala 41:38:@25004.4]
  wire  _T_63847; // @[Switch.scala 41:52:@25006.4]
  wire  output_17_6; // @[Switch.scala 41:38:@25007.4]
  wire  _T_63850; // @[Switch.scala 41:52:@25009.4]
  wire  output_17_7; // @[Switch.scala 41:38:@25010.4]
  wire  _T_63853; // @[Switch.scala 41:52:@25012.4]
  wire  output_17_8; // @[Switch.scala 41:38:@25013.4]
  wire  _T_63856; // @[Switch.scala 41:52:@25015.4]
  wire  output_17_9; // @[Switch.scala 41:38:@25016.4]
  wire  _T_63859; // @[Switch.scala 41:52:@25018.4]
  wire  output_17_10; // @[Switch.scala 41:38:@25019.4]
  wire  _T_63862; // @[Switch.scala 41:52:@25021.4]
  wire  output_17_11; // @[Switch.scala 41:38:@25022.4]
  wire  _T_63865; // @[Switch.scala 41:52:@25024.4]
  wire  output_17_12; // @[Switch.scala 41:38:@25025.4]
  wire  _T_63868; // @[Switch.scala 41:52:@25027.4]
  wire  output_17_13; // @[Switch.scala 41:38:@25028.4]
  wire  _T_63871; // @[Switch.scala 41:52:@25030.4]
  wire  output_17_14; // @[Switch.scala 41:38:@25031.4]
  wire  _T_63874; // @[Switch.scala 41:52:@25033.4]
  wire  output_17_15; // @[Switch.scala 41:38:@25034.4]
  wire  _T_63877; // @[Switch.scala 41:52:@25036.4]
  wire  output_17_16; // @[Switch.scala 41:38:@25037.4]
  wire  _T_63880; // @[Switch.scala 41:52:@25039.4]
  wire  output_17_17; // @[Switch.scala 41:38:@25040.4]
  wire  _T_63883; // @[Switch.scala 41:52:@25042.4]
  wire  output_17_18; // @[Switch.scala 41:38:@25043.4]
  wire  _T_63886; // @[Switch.scala 41:52:@25045.4]
  wire  output_17_19; // @[Switch.scala 41:38:@25046.4]
  wire  _T_63889; // @[Switch.scala 41:52:@25048.4]
  wire  output_17_20; // @[Switch.scala 41:38:@25049.4]
  wire  _T_63892; // @[Switch.scala 41:52:@25051.4]
  wire  output_17_21; // @[Switch.scala 41:38:@25052.4]
  wire  _T_63895; // @[Switch.scala 41:52:@25054.4]
  wire  output_17_22; // @[Switch.scala 41:38:@25055.4]
  wire  _T_63898; // @[Switch.scala 41:52:@25057.4]
  wire  output_17_23; // @[Switch.scala 41:38:@25058.4]
  wire  _T_63901; // @[Switch.scala 41:52:@25060.4]
  wire  output_17_24; // @[Switch.scala 41:38:@25061.4]
  wire  _T_63904; // @[Switch.scala 41:52:@25063.4]
  wire  output_17_25; // @[Switch.scala 41:38:@25064.4]
  wire  _T_63907; // @[Switch.scala 41:52:@25066.4]
  wire  output_17_26; // @[Switch.scala 41:38:@25067.4]
  wire  _T_63910; // @[Switch.scala 41:52:@25069.4]
  wire  output_17_27; // @[Switch.scala 41:38:@25070.4]
  wire  _T_63913; // @[Switch.scala 41:52:@25072.4]
  wire  output_17_28; // @[Switch.scala 41:38:@25073.4]
  wire  _T_63916; // @[Switch.scala 41:52:@25075.4]
  wire  output_17_29; // @[Switch.scala 41:38:@25076.4]
  wire  _T_63919; // @[Switch.scala 41:52:@25078.4]
  wire  output_17_30; // @[Switch.scala 41:38:@25079.4]
  wire  _T_63922; // @[Switch.scala 41:52:@25081.4]
  wire  output_17_31; // @[Switch.scala 41:38:@25082.4]
  wire  _T_63925; // @[Switch.scala 41:52:@25084.4]
  wire  output_17_32; // @[Switch.scala 41:38:@25085.4]
  wire  _T_63928; // @[Switch.scala 41:52:@25087.4]
  wire  output_17_33; // @[Switch.scala 41:38:@25088.4]
  wire  _T_63931; // @[Switch.scala 41:52:@25090.4]
  wire  output_17_34; // @[Switch.scala 41:38:@25091.4]
  wire  _T_63934; // @[Switch.scala 41:52:@25093.4]
  wire  output_17_35; // @[Switch.scala 41:38:@25094.4]
  wire  _T_63937; // @[Switch.scala 41:52:@25096.4]
  wire  output_17_36; // @[Switch.scala 41:38:@25097.4]
  wire  _T_63940; // @[Switch.scala 41:52:@25099.4]
  wire  output_17_37; // @[Switch.scala 41:38:@25100.4]
  wire  _T_63943; // @[Switch.scala 41:52:@25102.4]
  wire  output_17_38; // @[Switch.scala 41:38:@25103.4]
  wire  _T_63946; // @[Switch.scala 41:52:@25105.4]
  wire  output_17_39; // @[Switch.scala 41:38:@25106.4]
  wire  _T_63949; // @[Switch.scala 41:52:@25108.4]
  wire  output_17_40; // @[Switch.scala 41:38:@25109.4]
  wire  _T_63952; // @[Switch.scala 41:52:@25111.4]
  wire  output_17_41; // @[Switch.scala 41:38:@25112.4]
  wire  _T_63955; // @[Switch.scala 41:52:@25114.4]
  wire  output_17_42; // @[Switch.scala 41:38:@25115.4]
  wire  _T_63958; // @[Switch.scala 41:52:@25117.4]
  wire  output_17_43; // @[Switch.scala 41:38:@25118.4]
  wire  _T_63961; // @[Switch.scala 41:52:@25120.4]
  wire  output_17_44; // @[Switch.scala 41:38:@25121.4]
  wire  _T_63964; // @[Switch.scala 41:52:@25123.4]
  wire  output_17_45; // @[Switch.scala 41:38:@25124.4]
  wire  _T_63967; // @[Switch.scala 41:52:@25126.4]
  wire  output_17_46; // @[Switch.scala 41:38:@25127.4]
  wire  _T_63970; // @[Switch.scala 41:52:@25129.4]
  wire  output_17_47; // @[Switch.scala 41:38:@25130.4]
  wire  _T_63973; // @[Switch.scala 41:52:@25132.4]
  wire  output_17_48; // @[Switch.scala 41:38:@25133.4]
  wire  _T_63976; // @[Switch.scala 41:52:@25135.4]
  wire  output_17_49; // @[Switch.scala 41:38:@25136.4]
  wire  _T_63979; // @[Switch.scala 41:52:@25138.4]
  wire  output_17_50; // @[Switch.scala 41:38:@25139.4]
  wire  _T_63982; // @[Switch.scala 41:52:@25141.4]
  wire  output_17_51; // @[Switch.scala 41:38:@25142.4]
  wire  _T_63985; // @[Switch.scala 41:52:@25144.4]
  wire  output_17_52; // @[Switch.scala 41:38:@25145.4]
  wire  _T_63988; // @[Switch.scala 41:52:@25147.4]
  wire  output_17_53; // @[Switch.scala 41:38:@25148.4]
  wire  _T_63991; // @[Switch.scala 41:52:@25150.4]
  wire  output_17_54; // @[Switch.scala 41:38:@25151.4]
  wire  _T_63994; // @[Switch.scala 41:52:@25153.4]
  wire  output_17_55; // @[Switch.scala 41:38:@25154.4]
  wire  _T_63997; // @[Switch.scala 41:52:@25156.4]
  wire  output_17_56; // @[Switch.scala 41:38:@25157.4]
  wire  _T_64000; // @[Switch.scala 41:52:@25159.4]
  wire  output_17_57; // @[Switch.scala 41:38:@25160.4]
  wire  _T_64003; // @[Switch.scala 41:52:@25162.4]
  wire  output_17_58; // @[Switch.scala 41:38:@25163.4]
  wire  _T_64006; // @[Switch.scala 41:52:@25165.4]
  wire  output_17_59; // @[Switch.scala 41:38:@25166.4]
  wire  _T_64009; // @[Switch.scala 41:52:@25168.4]
  wire  output_17_60; // @[Switch.scala 41:38:@25169.4]
  wire  _T_64012; // @[Switch.scala 41:52:@25171.4]
  wire  output_17_61; // @[Switch.scala 41:38:@25172.4]
  wire  _T_64015; // @[Switch.scala 41:52:@25174.4]
  wire  output_17_62; // @[Switch.scala 41:38:@25175.4]
  wire  _T_64018; // @[Switch.scala 41:52:@25177.4]
  wire  output_17_63; // @[Switch.scala 41:38:@25178.4]
  wire [7:0] _T_64026; // @[Switch.scala 43:31:@25186.4]
  wire [15:0] _T_64034; // @[Switch.scala 43:31:@25194.4]
  wire [7:0] _T_64041; // @[Switch.scala 43:31:@25201.4]
  wire [31:0] _T_64050; // @[Switch.scala 43:31:@25210.4]
  wire [7:0] _T_64057; // @[Switch.scala 43:31:@25217.4]
  wire [15:0] _T_64065; // @[Switch.scala 43:31:@25225.4]
  wire [7:0] _T_64072; // @[Switch.scala 43:31:@25232.4]
  wire [31:0] _T_64081; // @[Switch.scala 43:31:@25241.4]
  wire [63:0] _T_64082; // @[Switch.scala 43:31:@25242.4]
  wire  _T_64086; // @[Switch.scala 41:52:@25245.4]
  wire  output_18_0; // @[Switch.scala 41:38:@25246.4]
  wire  _T_64089; // @[Switch.scala 41:52:@25248.4]
  wire  output_18_1; // @[Switch.scala 41:38:@25249.4]
  wire  _T_64092; // @[Switch.scala 41:52:@25251.4]
  wire  output_18_2; // @[Switch.scala 41:38:@25252.4]
  wire  _T_64095; // @[Switch.scala 41:52:@25254.4]
  wire  output_18_3; // @[Switch.scala 41:38:@25255.4]
  wire  _T_64098; // @[Switch.scala 41:52:@25257.4]
  wire  output_18_4; // @[Switch.scala 41:38:@25258.4]
  wire  _T_64101; // @[Switch.scala 41:52:@25260.4]
  wire  output_18_5; // @[Switch.scala 41:38:@25261.4]
  wire  _T_64104; // @[Switch.scala 41:52:@25263.4]
  wire  output_18_6; // @[Switch.scala 41:38:@25264.4]
  wire  _T_64107; // @[Switch.scala 41:52:@25266.4]
  wire  output_18_7; // @[Switch.scala 41:38:@25267.4]
  wire  _T_64110; // @[Switch.scala 41:52:@25269.4]
  wire  output_18_8; // @[Switch.scala 41:38:@25270.4]
  wire  _T_64113; // @[Switch.scala 41:52:@25272.4]
  wire  output_18_9; // @[Switch.scala 41:38:@25273.4]
  wire  _T_64116; // @[Switch.scala 41:52:@25275.4]
  wire  output_18_10; // @[Switch.scala 41:38:@25276.4]
  wire  _T_64119; // @[Switch.scala 41:52:@25278.4]
  wire  output_18_11; // @[Switch.scala 41:38:@25279.4]
  wire  _T_64122; // @[Switch.scala 41:52:@25281.4]
  wire  output_18_12; // @[Switch.scala 41:38:@25282.4]
  wire  _T_64125; // @[Switch.scala 41:52:@25284.4]
  wire  output_18_13; // @[Switch.scala 41:38:@25285.4]
  wire  _T_64128; // @[Switch.scala 41:52:@25287.4]
  wire  output_18_14; // @[Switch.scala 41:38:@25288.4]
  wire  _T_64131; // @[Switch.scala 41:52:@25290.4]
  wire  output_18_15; // @[Switch.scala 41:38:@25291.4]
  wire  _T_64134; // @[Switch.scala 41:52:@25293.4]
  wire  output_18_16; // @[Switch.scala 41:38:@25294.4]
  wire  _T_64137; // @[Switch.scala 41:52:@25296.4]
  wire  output_18_17; // @[Switch.scala 41:38:@25297.4]
  wire  _T_64140; // @[Switch.scala 41:52:@25299.4]
  wire  output_18_18; // @[Switch.scala 41:38:@25300.4]
  wire  _T_64143; // @[Switch.scala 41:52:@25302.4]
  wire  output_18_19; // @[Switch.scala 41:38:@25303.4]
  wire  _T_64146; // @[Switch.scala 41:52:@25305.4]
  wire  output_18_20; // @[Switch.scala 41:38:@25306.4]
  wire  _T_64149; // @[Switch.scala 41:52:@25308.4]
  wire  output_18_21; // @[Switch.scala 41:38:@25309.4]
  wire  _T_64152; // @[Switch.scala 41:52:@25311.4]
  wire  output_18_22; // @[Switch.scala 41:38:@25312.4]
  wire  _T_64155; // @[Switch.scala 41:52:@25314.4]
  wire  output_18_23; // @[Switch.scala 41:38:@25315.4]
  wire  _T_64158; // @[Switch.scala 41:52:@25317.4]
  wire  output_18_24; // @[Switch.scala 41:38:@25318.4]
  wire  _T_64161; // @[Switch.scala 41:52:@25320.4]
  wire  output_18_25; // @[Switch.scala 41:38:@25321.4]
  wire  _T_64164; // @[Switch.scala 41:52:@25323.4]
  wire  output_18_26; // @[Switch.scala 41:38:@25324.4]
  wire  _T_64167; // @[Switch.scala 41:52:@25326.4]
  wire  output_18_27; // @[Switch.scala 41:38:@25327.4]
  wire  _T_64170; // @[Switch.scala 41:52:@25329.4]
  wire  output_18_28; // @[Switch.scala 41:38:@25330.4]
  wire  _T_64173; // @[Switch.scala 41:52:@25332.4]
  wire  output_18_29; // @[Switch.scala 41:38:@25333.4]
  wire  _T_64176; // @[Switch.scala 41:52:@25335.4]
  wire  output_18_30; // @[Switch.scala 41:38:@25336.4]
  wire  _T_64179; // @[Switch.scala 41:52:@25338.4]
  wire  output_18_31; // @[Switch.scala 41:38:@25339.4]
  wire  _T_64182; // @[Switch.scala 41:52:@25341.4]
  wire  output_18_32; // @[Switch.scala 41:38:@25342.4]
  wire  _T_64185; // @[Switch.scala 41:52:@25344.4]
  wire  output_18_33; // @[Switch.scala 41:38:@25345.4]
  wire  _T_64188; // @[Switch.scala 41:52:@25347.4]
  wire  output_18_34; // @[Switch.scala 41:38:@25348.4]
  wire  _T_64191; // @[Switch.scala 41:52:@25350.4]
  wire  output_18_35; // @[Switch.scala 41:38:@25351.4]
  wire  _T_64194; // @[Switch.scala 41:52:@25353.4]
  wire  output_18_36; // @[Switch.scala 41:38:@25354.4]
  wire  _T_64197; // @[Switch.scala 41:52:@25356.4]
  wire  output_18_37; // @[Switch.scala 41:38:@25357.4]
  wire  _T_64200; // @[Switch.scala 41:52:@25359.4]
  wire  output_18_38; // @[Switch.scala 41:38:@25360.4]
  wire  _T_64203; // @[Switch.scala 41:52:@25362.4]
  wire  output_18_39; // @[Switch.scala 41:38:@25363.4]
  wire  _T_64206; // @[Switch.scala 41:52:@25365.4]
  wire  output_18_40; // @[Switch.scala 41:38:@25366.4]
  wire  _T_64209; // @[Switch.scala 41:52:@25368.4]
  wire  output_18_41; // @[Switch.scala 41:38:@25369.4]
  wire  _T_64212; // @[Switch.scala 41:52:@25371.4]
  wire  output_18_42; // @[Switch.scala 41:38:@25372.4]
  wire  _T_64215; // @[Switch.scala 41:52:@25374.4]
  wire  output_18_43; // @[Switch.scala 41:38:@25375.4]
  wire  _T_64218; // @[Switch.scala 41:52:@25377.4]
  wire  output_18_44; // @[Switch.scala 41:38:@25378.4]
  wire  _T_64221; // @[Switch.scala 41:52:@25380.4]
  wire  output_18_45; // @[Switch.scala 41:38:@25381.4]
  wire  _T_64224; // @[Switch.scala 41:52:@25383.4]
  wire  output_18_46; // @[Switch.scala 41:38:@25384.4]
  wire  _T_64227; // @[Switch.scala 41:52:@25386.4]
  wire  output_18_47; // @[Switch.scala 41:38:@25387.4]
  wire  _T_64230; // @[Switch.scala 41:52:@25389.4]
  wire  output_18_48; // @[Switch.scala 41:38:@25390.4]
  wire  _T_64233; // @[Switch.scala 41:52:@25392.4]
  wire  output_18_49; // @[Switch.scala 41:38:@25393.4]
  wire  _T_64236; // @[Switch.scala 41:52:@25395.4]
  wire  output_18_50; // @[Switch.scala 41:38:@25396.4]
  wire  _T_64239; // @[Switch.scala 41:52:@25398.4]
  wire  output_18_51; // @[Switch.scala 41:38:@25399.4]
  wire  _T_64242; // @[Switch.scala 41:52:@25401.4]
  wire  output_18_52; // @[Switch.scala 41:38:@25402.4]
  wire  _T_64245; // @[Switch.scala 41:52:@25404.4]
  wire  output_18_53; // @[Switch.scala 41:38:@25405.4]
  wire  _T_64248; // @[Switch.scala 41:52:@25407.4]
  wire  output_18_54; // @[Switch.scala 41:38:@25408.4]
  wire  _T_64251; // @[Switch.scala 41:52:@25410.4]
  wire  output_18_55; // @[Switch.scala 41:38:@25411.4]
  wire  _T_64254; // @[Switch.scala 41:52:@25413.4]
  wire  output_18_56; // @[Switch.scala 41:38:@25414.4]
  wire  _T_64257; // @[Switch.scala 41:52:@25416.4]
  wire  output_18_57; // @[Switch.scala 41:38:@25417.4]
  wire  _T_64260; // @[Switch.scala 41:52:@25419.4]
  wire  output_18_58; // @[Switch.scala 41:38:@25420.4]
  wire  _T_64263; // @[Switch.scala 41:52:@25422.4]
  wire  output_18_59; // @[Switch.scala 41:38:@25423.4]
  wire  _T_64266; // @[Switch.scala 41:52:@25425.4]
  wire  output_18_60; // @[Switch.scala 41:38:@25426.4]
  wire  _T_64269; // @[Switch.scala 41:52:@25428.4]
  wire  output_18_61; // @[Switch.scala 41:38:@25429.4]
  wire  _T_64272; // @[Switch.scala 41:52:@25431.4]
  wire  output_18_62; // @[Switch.scala 41:38:@25432.4]
  wire  _T_64275; // @[Switch.scala 41:52:@25434.4]
  wire  output_18_63; // @[Switch.scala 41:38:@25435.4]
  wire [7:0] _T_64283; // @[Switch.scala 43:31:@25443.4]
  wire [15:0] _T_64291; // @[Switch.scala 43:31:@25451.4]
  wire [7:0] _T_64298; // @[Switch.scala 43:31:@25458.4]
  wire [31:0] _T_64307; // @[Switch.scala 43:31:@25467.4]
  wire [7:0] _T_64314; // @[Switch.scala 43:31:@25474.4]
  wire [15:0] _T_64322; // @[Switch.scala 43:31:@25482.4]
  wire [7:0] _T_64329; // @[Switch.scala 43:31:@25489.4]
  wire [31:0] _T_64338; // @[Switch.scala 43:31:@25498.4]
  wire [63:0] _T_64339; // @[Switch.scala 43:31:@25499.4]
  wire  _T_64343; // @[Switch.scala 41:52:@25502.4]
  wire  output_19_0; // @[Switch.scala 41:38:@25503.4]
  wire  _T_64346; // @[Switch.scala 41:52:@25505.4]
  wire  output_19_1; // @[Switch.scala 41:38:@25506.4]
  wire  _T_64349; // @[Switch.scala 41:52:@25508.4]
  wire  output_19_2; // @[Switch.scala 41:38:@25509.4]
  wire  _T_64352; // @[Switch.scala 41:52:@25511.4]
  wire  output_19_3; // @[Switch.scala 41:38:@25512.4]
  wire  _T_64355; // @[Switch.scala 41:52:@25514.4]
  wire  output_19_4; // @[Switch.scala 41:38:@25515.4]
  wire  _T_64358; // @[Switch.scala 41:52:@25517.4]
  wire  output_19_5; // @[Switch.scala 41:38:@25518.4]
  wire  _T_64361; // @[Switch.scala 41:52:@25520.4]
  wire  output_19_6; // @[Switch.scala 41:38:@25521.4]
  wire  _T_64364; // @[Switch.scala 41:52:@25523.4]
  wire  output_19_7; // @[Switch.scala 41:38:@25524.4]
  wire  _T_64367; // @[Switch.scala 41:52:@25526.4]
  wire  output_19_8; // @[Switch.scala 41:38:@25527.4]
  wire  _T_64370; // @[Switch.scala 41:52:@25529.4]
  wire  output_19_9; // @[Switch.scala 41:38:@25530.4]
  wire  _T_64373; // @[Switch.scala 41:52:@25532.4]
  wire  output_19_10; // @[Switch.scala 41:38:@25533.4]
  wire  _T_64376; // @[Switch.scala 41:52:@25535.4]
  wire  output_19_11; // @[Switch.scala 41:38:@25536.4]
  wire  _T_64379; // @[Switch.scala 41:52:@25538.4]
  wire  output_19_12; // @[Switch.scala 41:38:@25539.4]
  wire  _T_64382; // @[Switch.scala 41:52:@25541.4]
  wire  output_19_13; // @[Switch.scala 41:38:@25542.4]
  wire  _T_64385; // @[Switch.scala 41:52:@25544.4]
  wire  output_19_14; // @[Switch.scala 41:38:@25545.4]
  wire  _T_64388; // @[Switch.scala 41:52:@25547.4]
  wire  output_19_15; // @[Switch.scala 41:38:@25548.4]
  wire  _T_64391; // @[Switch.scala 41:52:@25550.4]
  wire  output_19_16; // @[Switch.scala 41:38:@25551.4]
  wire  _T_64394; // @[Switch.scala 41:52:@25553.4]
  wire  output_19_17; // @[Switch.scala 41:38:@25554.4]
  wire  _T_64397; // @[Switch.scala 41:52:@25556.4]
  wire  output_19_18; // @[Switch.scala 41:38:@25557.4]
  wire  _T_64400; // @[Switch.scala 41:52:@25559.4]
  wire  output_19_19; // @[Switch.scala 41:38:@25560.4]
  wire  _T_64403; // @[Switch.scala 41:52:@25562.4]
  wire  output_19_20; // @[Switch.scala 41:38:@25563.4]
  wire  _T_64406; // @[Switch.scala 41:52:@25565.4]
  wire  output_19_21; // @[Switch.scala 41:38:@25566.4]
  wire  _T_64409; // @[Switch.scala 41:52:@25568.4]
  wire  output_19_22; // @[Switch.scala 41:38:@25569.4]
  wire  _T_64412; // @[Switch.scala 41:52:@25571.4]
  wire  output_19_23; // @[Switch.scala 41:38:@25572.4]
  wire  _T_64415; // @[Switch.scala 41:52:@25574.4]
  wire  output_19_24; // @[Switch.scala 41:38:@25575.4]
  wire  _T_64418; // @[Switch.scala 41:52:@25577.4]
  wire  output_19_25; // @[Switch.scala 41:38:@25578.4]
  wire  _T_64421; // @[Switch.scala 41:52:@25580.4]
  wire  output_19_26; // @[Switch.scala 41:38:@25581.4]
  wire  _T_64424; // @[Switch.scala 41:52:@25583.4]
  wire  output_19_27; // @[Switch.scala 41:38:@25584.4]
  wire  _T_64427; // @[Switch.scala 41:52:@25586.4]
  wire  output_19_28; // @[Switch.scala 41:38:@25587.4]
  wire  _T_64430; // @[Switch.scala 41:52:@25589.4]
  wire  output_19_29; // @[Switch.scala 41:38:@25590.4]
  wire  _T_64433; // @[Switch.scala 41:52:@25592.4]
  wire  output_19_30; // @[Switch.scala 41:38:@25593.4]
  wire  _T_64436; // @[Switch.scala 41:52:@25595.4]
  wire  output_19_31; // @[Switch.scala 41:38:@25596.4]
  wire  _T_64439; // @[Switch.scala 41:52:@25598.4]
  wire  output_19_32; // @[Switch.scala 41:38:@25599.4]
  wire  _T_64442; // @[Switch.scala 41:52:@25601.4]
  wire  output_19_33; // @[Switch.scala 41:38:@25602.4]
  wire  _T_64445; // @[Switch.scala 41:52:@25604.4]
  wire  output_19_34; // @[Switch.scala 41:38:@25605.4]
  wire  _T_64448; // @[Switch.scala 41:52:@25607.4]
  wire  output_19_35; // @[Switch.scala 41:38:@25608.4]
  wire  _T_64451; // @[Switch.scala 41:52:@25610.4]
  wire  output_19_36; // @[Switch.scala 41:38:@25611.4]
  wire  _T_64454; // @[Switch.scala 41:52:@25613.4]
  wire  output_19_37; // @[Switch.scala 41:38:@25614.4]
  wire  _T_64457; // @[Switch.scala 41:52:@25616.4]
  wire  output_19_38; // @[Switch.scala 41:38:@25617.4]
  wire  _T_64460; // @[Switch.scala 41:52:@25619.4]
  wire  output_19_39; // @[Switch.scala 41:38:@25620.4]
  wire  _T_64463; // @[Switch.scala 41:52:@25622.4]
  wire  output_19_40; // @[Switch.scala 41:38:@25623.4]
  wire  _T_64466; // @[Switch.scala 41:52:@25625.4]
  wire  output_19_41; // @[Switch.scala 41:38:@25626.4]
  wire  _T_64469; // @[Switch.scala 41:52:@25628.4]
  wire  output_19_42; // @[Switch.scala 41:38:@25629.4]
  wire  _T_64472; // @[Switch.scala 41:52:@25631.4]
  wire  output_19_43; // @[Switch.scala 41:38:@25632.4]
  wire  _T_64475; // @[Switch.scala 41:52:@25634.4]
  wire  output_19_44; // @[Switch.scala 41:38:@25635.4]
  wire  _T_64478; // @[Switch.scala 41:52:@25637.4]
  wire  output_19_45; // @[Switch.scala 41:38:@25638.4]
  wire  _T_64481; // @[Switch.scala 41:52:@25640.4]
  wire  output_19_46; // @[Switch.scala 41:38:@25641.4]
  wire  _T_64484; // @[Switch.scala 41:52:@25643.4]
  wire  output_19_47; // @[Switch.scala 41:38:@25644.4]
  wire  _T_64487; // @[Switch.scala 41:52:@25646.4]
  wire  output_19_48; // @[Switch.scala 41:38:@25647.4]
  wire  _T_64490; // @[Switch.scala 41:52:@25649.4]
  wire  output_19_49; // @[Switch.scala 41:38:@25650.4]
  wire  _T_64493; // @[Switch.scala 41:52:@25652.4]
  wire  output_19_50; // @[Switch.scala 41:38:@25653.4]
  wire  _T_64496; // @[Switch.scala 41:52:@25655.4]
  wire  output_19_51; // @[Switch.scala 41:38:@25656.4]
  wire  _T_64499; // @[Switch.scala 41:52:@25658.4]
  wire  output_19_52; // @[Switch.scala 41:38:@25659.4]
  wire  _T_64502; // @[Switch.scala 41:52:@25661.4]
  wire  output_19_53; // @[Switch.scala 41:38:@25662.4]
  wire  _T_64505; // @[Switch.scala 41:52:@25664.4]
  wire  output_19_54; // @[Switch.scala 41:38:@25665.4]
  wire  _T_64508; // @[Switch.scala 41:52:@25667.4]
  wire  output_19_55; // @[Switch.scala 41:38:@25668.4]
  wire  _T_64511; // @[Switch.scala 41:52:@25670.4]
  wire  output_19_56; // @[Switch.scala 41:38:@25671.4]
  wire  _T_64514; // @[Switch.scala 41:52:@25673.4]
  wire  output_19_57; // @[Switch.scala 41:38:@25674.4]
  wire  _T_64517; // @[Switch.scala 41:52:@25676.4]
  wire  output_19_58; // @[Switch.scala 41:38:@25677.4]
  wire  _T_64520; // @[Switch.scala 41:52:@25679.4]
  wire  output_19_59; // @[Switch.scala 41:38:@25680.4]
  wire  _T_64523; // @[Switch.scala 41:52:@25682.4]
  wire  output_19_60; // @[Switch.scala 41:38:@25683.4]
  wire  _T_64526; // @[Switch.scala 41:52:@25685.4]
  wire  output_19_61; // @[Switch.scala 41:38:@25686.4]
  wire  _T_64529; // @[Switch.scala 41:52:@25688.4]
  wire  output_19_62; // @[Switch.scala 41:38:@25689.4]
  wire  _T_64532; // @[Switch.scala 41:52:@25691.4]
  wire  output_19_63; // @[Switch.scala 41:38:@25692.4]
  wire [7:0] _T_64540; // @[Switch.scala 43:31:@25700.4]
  wire [15:0] _T_64548; // @[Switch.scala 43:31:@25708.4]
  wire [7:0] _T_64555; // @[Switch.scala 43:31:@25715.4]
  wire [31:0] _T_64564; // @[Switch.scala 43:31:@25724.4]
  wire [7:0] _T_64571; // @[Switch.scala 43:31:@25731.4]
  wire [15:0] _T_64579; // @[Switch.scala 43:31:@25739.4]
  wire [7:0] _T_64586; // @[Switch.scala 43:31:@25746.4]
  wire [31:0] _T_64595; // @[Switch.scala 43:31:@25755.4]
  wire [63:0] _T_64596; // @[Switch.scala 43:31:@25756.4]
  wire  _T_64600; // @[Switch.scala 41:52:@25759.4]
  wire  output_20_0; // @[Switch.scala 41:38:@25760.4]
  wire  _T_64603; // @[Switch.scala 41:52:@25762.4]
  wire  output_20_1; // @[Switch.scala 41:38:@25763.4]
  wire  _T_64606; // @[Switch.scala 41:52:@25765.4]
  wire  output_20_2; // @[Switch.scala 41:38:@25766.4]
  wire  _T_64609; // @[Switch.scala 41:52:@25768.4]
  wire  output_20_3; // @[Switch.scala 41:38:@25769.4]
  wire  _T_64612; // @[Switch.scala 41:52:@25771.4]
  wire  output_20_4; // @[Switch.scala 41:38:@25772.4]
  wire  _T_64615; // @[Switch.scala 41:52:@25774.4]
  wire  output_20_5; // @[Switch.scala 41:38:@25775.4]
  wire  _T_64618; // @[Switch.scala 41:52:@25777.4]
  wire  output_20_6; // @[Switch.scala 41:38:@25778.4]
  wire  _T_64621; // @[Switch.scala 41:52:@25780.4]
  wire  output_20_7; // @[Switch.scala 41:38:@25781.4]
  wire  _T_64624; // @[Switch.scala 41:52:@25783.4]
  wire  output_20_8; // @[Switch.scala 41:38:@25784.4]
  wire  _T_64627; // @[Switch.scala 41:52:@25786.4]
  wire  output_20_9; // @[Switch.scala 41:38:@25787.4]
  wire  _T_64630; // @[Switch.scala 41:52:@25789.4]
  wire  output_20_10; // @[Switch.scala 41:38:@25790.4]
  wire  _T_64633; // @[Switch.scala 41:52:@25792.4]
  wire  output_20_11; // @[Switch.scala 41:38:@25793.4]
  wire  _T_64636; // @[Switch.scala 41:52:@25795.4]
  wire  output_20_12; // @[Switch.scala 41:38:@25796.4]
  wire  _T_64639; // @[Switch.scala 41:52:@25798.4]
  wire  output_20_13; // @[Switch.scala 41:38:@25799.4]
  wire  _T_64642; // @[Switch.scala 41:52:@25801.4]
  wire  output_20_14; // @[Switch.scala 41:38:@25802.4]
  wire  _T_64645; // @[Switch.scala 41:52:@25804.4]
  wire  output_20_15; // @[Switch.scala 41:38:@25805.4]
  wire  _T_64648; // @[Switch.scala 41:52:@25807.4]
  wire  output_20_16; // @[Switch.scala 41:38:@25808.4]
  wire  _T_64651; // @[Switch.scala 41:52:@25810.4]
  wire  output_20_17; // @[Switch.scala 41:38:@25811.4]
  wire  _T_64654; // @[Switch.scala 41:52:@25813.4]
  wire  output_20_18; // @[Switch.scala 41:38:@25814.4]
  wire  _T_64657; // @[Switch.scala 41:52:@25816.4]
  wire  output_20_19; // @[Switch.scala 41:38:@25817.4]
  wire  _T_64660; // @[Switch.scala 41:52:@25819.4]
  wire  output_20_20; // @[Switch.scala 41:38:@25820.4]
  wire  _T_64663; // @[Switch.scala 41:52:@25822.4]
  wire  output_20_21; // @[Switch.scala 41:38:@25823.4]
  wire  _T_64666; // @[Switch.scala 41:52:@25825.4]
  wire  output_20_22; // @[Switch.scala 41:38:@25826.4]
  wire  _T_64669; // @[Switch.scala 41:52:@25828.4]
  wire  output_20_23; // @[Switch.scala 41:38:@25829.4]
  wire  _T_64672; // @[Switch.scala 41:52:@25831.4]
  wire  output_20_24; // @[Switch.scala 41:38:@25832.4]
  wire  _T_64675; // @[Switch.scala 41:52:@25834.4]
  wire  output_20_25; // @[Switch.scala 41:38:@25835.4]
  wire  _T_64678; // @[Switch.scala 41:52:@25837.4]
  wire  output_20_26; // @[Switch.scala 41:38:@25838.4]
  wire  _T_64681; // @[Switch.scala 41:52:@25840.4]
  wire  output_20_27; // @[Switch.scala 41:38:@25841.4]
  wire  _T_64684; // @[Switch.scala 41:52:@25843.4]
  wire  output_20_28; // @[Switch.scala 41:38:@25844.4]
  wire  _T_64687; // @[Switch.scala 41:52:@25846.4]
  wire  output_20_29; // @[Switch.scala 41:38:@25847.4]
  wire  _T_64690; // @[Switch.scala 41:52:@25849.4]
  wire  output_20_30; // @[Switch.scala 41:38:@25850.4]
  wire  _T_64693; // @[Switch.scala 41:52:@25852.4]
  wire  output_20_31; // @[Switch.scala 41:38:@25853.4]
  wire  _T_64696; // @[Switch.scala 41:52:@25855.4]
  wire  output_20_32; // @[Switch.scala 41:38:@25856.4]
  wire  _T_64699; // @[Switch.scala 41:52:@25858.4]
  wire  output_20_33; // @[Switch.scala 41:38:@25859.4]
  wire  _T_64702; // @[Switch.scala 41:52:@25861.4]
  wire  output_20_34; // @[Switch.scala 41:38:@25862.4]
  wire  _T_64705; // @[Switch.scala 41:52:@25864.4]
  wire  output_20_35; // @[Switch.scala 41:38:@25865.4]
  wire  _T_64708; // @[Switch.scala 41:52:@25867.4]
  wire  output_20_36; // @[Switch.scala 41:38:@25868.4]
  wire  _T_64711; // @[Switch.scala 41:52:@25870.4]
  wire  output_20_37; // @[Switch.scala 41:38:@25871.4]
  wire  _T_64714; // @[Switch.scala 41:52:@25873.4]
  wire  output_20_38; // @[Switch.scala 41:38:@25874.4]
  wire  _T_64717; // @[Switch.scala 41:52:@25876.4]
  wire  output_20_39; // @[Switch.scala 41:38:@25877.4]
  wire  _T_64720; // @[Switch.scala 41:52:@25879.4]
  wire  output_20_40; // @[Switch.scala 41:38:@25880.4]
  wire  _T_64723; // @[Switch.scala 41:52:@25882.4]
  wire  output_20_41; // @[Switch.scala 41:38:@25883.4]
  wire  _T_64726; // @[Switch.scala 41:52:@25885.4]
  wire  output_20_42; // @[Switch.scala 41:38:@25886.4]
  wire  _T_64729; // @[Switch.scala 41:52:@25888.4]
  wire  output_20_43; // @[Switch.scala 41:38:@25889.4]
  wire  _T_64732; // @[Switch.scala 41:52:@25891.4]
  wire  output_20_44; // @[Switch.scala 41:38:@25892.4]
  wire  _T_64735; // @[Switch.scala 41:52:@25894.4]
  wire  output_20_45; // @[Switch.scala 41:38:@25895.4]
  wire  _T_64738; // @[Switch.scala 41:52:@25897.4]
  wire  output_20_46; // @[Switch.scala 41:38:@25898.4]
  wire  _T_64741; // @[Switch.scala 41:52:@25900.4]
  wire  output_20_47; // @[Switch.scala 41:38:@25901.4]
  wire  _T_64744; // @[Switch.scala 41:52:@25903.4]
  wire  output_20_48; // @[Switch.scala 41:38:@25904.4]
  wire  _T_64747; // @[Switch.scala 41:52:@25906.4]
  wire  output_20_49; // @[Switch.scala 41:38:@25907.4]
  wire  _T_64750; // @[Switch.scala 41:52:@25909.4]
  wire  output_20_50; // @[Switch.scala 41:38:@25910.4]
  wire  _T_64753; // @[Switch.scala 41:52:@25912.4]
  wire  output_20_51; // @[Switch.scala 41:38:@25913.4]
  wire  _T_64756; // @[Switch.scala 41:52:@25915.4]
  wire  output_20_52; // @[Switch.scala 41:38:@25916.4]
  wire  _T_64759; // @[Switch.scala 41:52:@25918.4]
  wire  output_20_53; // @[Switch.scala 41:38:@25919.4]
  wire  _T_64762; // @[Switch.scala 41:52:@25921.4]
  wire  output_20_54; // @[Switch.scala 41:38:@25922.4]
  wire  _T_64765; // @[Switch.scala 41:52:@25924.4]
  wire  output_20_55; // @[Switch.scala 41:38:@25925.4]
  wire  _T_64768; // @[Switch.scala 41:52:@25927.4]
  wire  output_20_56; // @[Switch.scala 41:38:@25928.4]
  wire  _T_64771; // @[Switch.scala 41:52:@25930.4]
  wire  output_20_57; // @[Switch.scala 41:38:@25931.4]
  wire  _T_64774; // @[Switch.scala 41:52:@25933.4]
  wire  output_20_58; // @[Switch.scala 41:38:@25934.4]
  wire  _T_64777; // @[Switch.scala 41:52:@25936.4]
  wire  output_20_59; // @[Switch.scala 41:38:@25937.4]
  wire  _T_64780; // @[Switch.scala 41:52:@25939.4]
  wire  output_20_60; // @[Switch.scala 41:38:@25940.4]
  wire  _T_64783; // @[Switch.scala 41:52:@25942.4]
  wire  output_20_61; // @[Switch.scala 41:38:@25943.4]
  wire  _T_64786; // @[Switch.scala 41:52:@25945.4]
  wire  output_20_62; // @[Switch.scala 41:38:@25946.4]
  wire  _T_64789; // @[Switch.scala 41:52:@25948.4]
  wire  output_20_63; // @[Switch.scala 41:38:@25949.4]
  wire [7:0] _T_64797; // @[Switch.scala 43:31:@25957.4]
  wire [15:0] _T_64805; // @[Switch.scala 43:31:@25965.4]
  wire [7:0] _T_64812; // @[Switch.scala 43:31:@25972.4]
  wire [31:0] _T_64821; // @[Switch.scala 43:31:@25981.4]
  wire [7:0] _T_64828; // @[Switch.scala 43:31:@25988.4]
  wire [15:0] _T_64836; // @[Switch.scala 43:31:@25996.4]
  wire [7:0] _T_64843; // @[Switch.scala 43:31:@26003.4]
  wire [31:0] _T_64852; // @[Switch.scala 43:31:@26012.4]
  wire [63:0] _T_64853; // @[Switch.scala 43:31:@26013.4]
  wire  _T_64857; // @[Switch.scala 41:52:@26016.4]
  wire  output_21_0; // @[Switch.scala 41:38:@26017.4]
  wire  _T_64860; // @[Switch.scala 41:52:@26019.4]
  wire  output_21_1; // @[Switch.scala 41:38:@26020.4]
  wire  _T_64863; // @[Switch.scala 41:52:@26022.4]
  wire  output_21_2; // @[Switch.scala 41:38:@26023.4]
  wire  _T_64866; // @[Switch.scala 41:52:@26025.4]
  wire  output_21_3; // @[Switch.scala 41:38:@26026.4]
  wire  _T_64869; // @[Switch.scala 41:52:@26028.4]
  wire  output_21_4; // @[Switch.scala 41:38:@26029.4]
  wire  _T_64872; // @[Switch.scala 41:52:@26031.4]
  wire  output_21_5; // @[Switch.scala 41:38:@26032.4]
  wire  _T_64875; // @[Switch.scala 41:52:@26034.4]
  wire  output_21_6; // @[Switch.scala 41:38:@26035.4]
  wire  _T_64878; // @[Switch.scala 41:52:@26037.4]
  wire  output_21_7; // @[Switch.scala 41:38:@26038.4]
  wire  _T_64881; // @[Switch.scala 41:52:@26040.4]
  wire  output_21_8; // @[Switch.scala 41:38:@26041.4]
  wire  _T_64884; // @[Switch.scala 41:52:@26043.4]
  wire  output_21_9; // @[Switch.scala 41:38:@26044.4]
  wire  _T_64887; // @[Switch.scala 41:52:@26046.4]
  wire  output_21_10; // @[Switch.scala 41:38:@26047.4]
  wire  _T_64890; // @[Switch.scala 41:52:@26049.4]
  wire  output_21_11; // @[Switch.scala 41:38:@26050.4]
  wire  _T_64893; // @[Switch.scala 41:52:@26052.4]
  wire  output_21_12; // @[Switch.scala 41:38:@26053.4]
  wire  _T_64896; // @[Switch.scala 41:52:@26055.4]
  wire  output_21_13; // @[Switch.scala 41:38:@26056.4]
  wire  _T_64899; // @[Switch.scala 41:52:@26058.4]
  wire  output_21_14; // @[Switch.scala 41:38:@26059.4]
  wire  _T_64902; // @[Switch.scala 41:52:@26061.4]
  wire  output_21_15; // @[Switch.scala 41:38:@26062.4]
  wire  _T_64905; // @[Switch.scala 41:52:@26064.4]
  wire  output_21_16; // @[Switch.scala 41:38:@26065.4]
  wire  _T_64908; // @[Switch.scala 41:52:@26067.4]
  wire  output_21_17; // @[Switch.scala 41:38:@26068.4]
  wire  _T_64911; // @[Switch.scala 41:52:@26070.4]
  wire  output_21_18; // @[Switch.scala 41:38:@26071.4]
  wire  _T_64914; // @[Switch.scala 41:52:@26073.4]
  wire  output_21_19; // @[Switch.scala 41:38:@26074.4]
  wire  _T_64917; // @[Switch.scala 41:52:@26076.4]
  wire  output_21_20; // @[Switch.scala 41:38:@26077.4]
  wire  _T_64920; // @[Switch.scala 41:52:@26079.4]
  wire  output_21_21; // @[Switch.scala 41:38:@26080.4]
  wire  _T_64923; // @[Switch.scala 41:52:@26082.4]
  wire  output_21_22; // @[Switch.scala 41:38:@26083.4]
  wire  _T_64926; // @[Switch.scala 41:52:@26085.4]
  wire  output_21_23; // @[Switch.scala 41:38:@26086.4]
  wire  _T_64929; // @[Switch.scala 41:52:@26088.4]
  wire  output_21_24; // @[Switch.scala 41:38:@26089.4]
  wire  _T_64932; // @[Switch.scala 41:52:@26091.4]
  wire  output_21_25; // @[Switch.scala 41:38:@26092.4]
  wire  _T_64935; // @[Switch.scala 41:52:@26094.4]
  wire  output_21_26; // @[Switch.scala 41:38:@26095.4]
  wire  _T_64938; // @[Switch.scala 41:52:@26097.4]
  wire  output_21_27; // @[Switch.scala 41:38:@26098.4]
  wire  _T_64941; // @[Switch.scala 41:52:@26100.4]
  wire  output_21_28; // @[Switch.scala 41:38:@26101.4]
  wire  _T_64944; // @[Switch.scala 41:52:@26103.4]
  wire  output_21_29; // @[Switch.scala 41:38:@26104.4]
  wire  _T_64947; // @[Switch.scala 41:52:@26106.4]
  wire  output_21_30; // @[Switch.scala 41:38:@26107.4]
  wire  _T_64950; // @[Switch.scala 41:52:@26109.4]
  wire  output_21_31; // @[Switch.scala 41:38:@26110.4]
  wire  _T_64953; // @[Switch.scala 41:52:@26112.4]
  wire  output_21_32; // @[Switch.scala 41:38:@26113.4]
  wire  _T_64956; // @[Switch.scala 41:52:@26115.4]
  wire  output_21_33; // @[Switch.scala 41:38:@26116.4]
  wire  _T_64959; // @[Switch.scala 41:52:@26118.4]
  wire  output_21_34; // @[Switch.scala 41:38:@26119.4]
  wire  _T_64962; // @[Switch.scala 41:52:@26121.4]
  wire  output_21_35; // @[Switch.scala 41:38:@26122.4]
  wire  _T_64965; // @[Switch.scala 41:52:@26124.4]
  wire  output_21_36; // @[Switch.scala 41:38:@26125.4]
  wire  _T_64968; // @[Switch.scala 41:52:@26127.4]
  wire  output_21_37; // @[Switch.scala 41:38:@26128.4]
  wire  _T_64971; // @[Switch.scala 41:52:@26130.4]
  wire  output_21_38; // @[Switch.scala 41:38:@26131.4]
  wire  _T_64974; // @[Switch.scala 41:52:@26133.4]
  wire  output_21_39; // @[Switch.scala 41:38:@26134.4]
  wire  _T_64977; // @[Switch.scala 41:52:@26136.4]
  wire  output_21_40; // @[Switch.scala 41:38:@26137.4]
  wire  _T_64980; // @[Switch.scala 41:52:@26139.4]
  wire  output_21_41; // @[Switch.scala 41:38:@26140.4]
  wire  _T_64983; // @[Switch.scala 41:52:@26142.4]
  wire  output_21_42; // @[Switch.scala 41:38:@26143.4]
  wire  _T_64986; // @[Switch.scala 41:52:@26145.4]
  wire  output_21_43; // @[Switch.scala 41:38:@26146.4]
  wire  _T_64989; // @[Switch.scala 41:52:@26148.4]
  wire  output_21_44; // @[Switch.scala 41:38:@26149.4]
  wire  _T_64992; // @[Switch.scala 41:52:@26151.4]
  wire  output_21_45; // @[Switch.scala 41:38:@26152.4]
  wire  _T_64995; // @[Switch.scala 41:52:@26154.4]
  wire  output_21_46; // @[Switch.scala 41:38:@26155.4]
  wire  _T_64998; // @[Switch.scala 41:52:@26157.4]
  wire  output_21_47; // @[Switch.scala 41:38:@26158.4]
  wire  _T_65001; // @[Switch.scala 41:52:@26160.4]
  wire  output_21_48; // @[Switch.scala 41:38:@26161.4]
  wire  _T_65004; // @[Switch.scala 41:52:@26163.4]
  wire  output_21_49; // @[Switch.scala 41:38:@26164.4]
  wire  _T_65007; // @[Switch.scala 41:52:@26166.4]
  wire  output_21_50; // @[Switch.scala 41:38:@26167.4]
  wire  _T_65010; // @[Switch.scala 41:52:@26169.4]
  wire  output_21_51; // @[Switch.scala 41:38:@26170.4]
  wire  _T_65013; // @[Switch.scala 41:52:@26172.4]
  wire  output_21_52; // @[Switch.scala 41:38:@26173.4]
  wire  _T_65016; // @[Switch.scala 41:52:@26175.4]
  wire  output_21_53; // @[Switch.scala 41:38:@26176.4]
  wire  _T_65019; // @[Switch.scala 41:52:@26178.4]
  wire  output_21_54; // @[Switch.scala 41:38:@26179.4]
  wire  _T_65022; // @[Switch.scala 41:52:@26181.4]
  wire  output_21_55; // @[Switch.scala 41:38:@26182.4]
  wire  _T_65025; // @[Switch.scala 41:52:@26184.4]
  wire  output_21_56; // @[Switch.scala 41:38:@26185.4]
  wire  _T_65028; // @[Switch.scala 41:52:@26187.4]
  wire  output_21_57; // @[Switch.scala 41:38:@26188.4]
  wire  _T_65031; // @[Switch.scala 41:52:@26190.4]
  wire  output_21_58; // @[Switch.scala 41:38:@26191.4]
  wire  _T_65034; // @[Switch.scala 41:52:@26193.4]
  wire  output_21_59; // @[Switch.scala 41:38:@26194.4]
  wire  _T_65037; // @[Switch.scala 41:52:@26196.4]
  wire  output_21_60; // @[Switch.scala 41:38:@26197.4]
  wire  _T_65040; // @[Switch.scala 41:52:@26199.4]
  wire  output_21_61; // @[Switch.scala 41:38:@26200.4]
  wire  _T_65043; // @[Switch.scala 41:52:@26202.4]
  wire  output_21_62; // @[Switch.scala 41:38:@26203.4]
  wire  _T_65046; // @[Switch.scala 41:52:@26205.4]
  wire  output_21_63; // @[Switch.scala 41:38:@26206.4]
  wire [7:0] _T_65054; // @[Switch.scala 43:31:@26214.4]
  wire [15:0] _T_65062; // @[Switch.scala 43:31:@26222.4]
  wire [7:0] _T_65069; // @[Switch.scala 43:31:@26229.4]
  wire [31:0] _T_65078; // @[Switch.scala 43:31:@26238.4]
  wire [7:0] _T_65085; // @[Switch.scala 43:31:@26245.4]
  wire [15:0] _T_65093; // @[Switch.scala 43:31:@26253.4]
  wire [7:0] _T_65100; // @[Switch.scala 43:31:@26260.4]
  wire [31:0] _T_65109; // @[Switch.scala 43:31:@26269.4]
  wire [63:0] _T_65110; // @[Switch.scala 43:31:@26270.4]
  wire  _T_65114; // @[Switch.scala 41:52:@26273.4]
  wire  output_22_0; // @[Switch.scala 41:38:@26274.4]
  wire  _T_65117; // @[Switch.scala 41:52:@26276.4]
  wire  output_22_1; // @[Switch.scala 41:38:@26277.4]
  wire  _T_65120; // @[Switch.scala 41:52:@26279.4]
  wire  output_22_2; // @[Switch.scala 41:38:@26280.4]
  wire  _T_65123; // @[Switch.scala 41:52:@26282.4]
  wire  output_22_3; // @[Switch.scala 41:38:@26283.4]
  wire  _T_65126; // @[Switch.scala 41:52:@26285.4]
  wire  output_22_4; // @[Switch.scala 41:38:@26286.4]
  wire  _T_65129; // @[Switch.scala 41:52:@26288.4]
  wire  output_22_5; // @[Switch.scala 41:38:@26289.4]
  wire  _T_65132; // @[Switch.scala 41:52:@26291.4]
  wire  output_22_6; // @[Switch.scala 41:38:@26292.4]
  wire  _T_65135; // @[Switch.scala 41:52:@26294.4]
  wire  output_22_7; // @[Switch.scala 41:38:@26295.4]
  wire  _T_65138; // @[Switch.scala 41:52:@26297.4]
  wire  output_22_8; // @[Switch.scala 41:38:@26298.4]
  wire  _T_65141; // @[Switch.scala 41:52:@26300.4]
  wire  output_22_9; // @[Switch.scala 41:38:@26301.4]
  wire  _T_65144; // @[Switch.scala 41:52:@26303.4]
  wire  output_22_10; // @[Switch.scala 41:38:@26304.4]
  wire  _T_65147; // @[Switch.scala 41:52:@26306.4]
  wire  output_22_11; // @[Switch.scala 41:38:@26307.4]
  wire  _T_65150; // @[Switch.scala 41:52:@26309.4]
  wire  output_22_12; // @[Switch.scala 41:38:@26310.4]
  wire  _T_65153; // @[Switch.scala 41:52:@26312.4]
  wire  output_22_13; // @[Switch.scala 41:38:@26313.4]
  wire  _T_65156; // @[Switch.scala 41:52:@26315.4]
  wire  output_22_14; // @[Switch.scala 41:38:@26316.4]
  wire  _T_65159; // @[Switch.scala 41:52:@26318.4]
  wire  output_22_15; // @[Switch.scala 41:38:@26319.4]
  wire  _T_65162; // @[Switch.scala 41:52:@26321.4]
  wire  output_22_16; // @[Switch.scala 41:38:@26322.4]
  wire  _T_65165; // @[Switch.scala 41:52:@26324.4]
  wire  output_22_17; // @[Switch.scala 41:38:@26325.4]
  wire  _T_65168; // @[Switch.scala 41:52:@26327.4]
  wire  output_22_18; // @[Switch.scala 41:38:@26328.4]
  wire  _T_65171; // @[Switch.scala 41:52:@26330.4]
  wire  output_22_19; // @[Switch.scala 41:38:@26331.4]
  wire  _T_65174; // @[Switch.scala 41:52:@26333.4]
  wire  output_22_20; // @[Switch.scala 41:38:@26334.4]
  wire  _T_65177; // @[Switch.scala 41:52:@26336.4]
  wire  output_22_21; // @[Switch.scala 41:38:@26337.4]
  wire  _T_65180; // @[Switch.scala 41:52:@26339.4]
  wire  output_22_22; // @[Switch.scala 41:38:@26340.4]
  wire  _T_65183; // @[Switch.scala 41:52:@26342.4]
  wire  output_22_23; // @[Switch.scala 41:38:@26343.4]
  wire  _T_65186; // @[Switch.scala 41:52:@26345.4]
  wire  output_22_24; // @[Switch.scala 41:38:@26346.4]
  wire  _T_65189; // @[Switch.scala 41:52:@26348.4]
  wire  output_22_25; // @[Switch.scala 41:38:@26349.4]
  wire  _T_65192; // @[Switch.scala 41:52:@26351.4]
  wire  output_22_26; // @[Switch.scala 41:38:@26352.4]
  wire  _T_65195; // @[Switch.scala 41:52:@26354.4]
  wire  output_22_27; // @[Switch.scala 41:38:@26355.4]
  wire  _T_65198; // @[Switch.scala 41:52:@26357.4]
  wire  output_22_28; // @[Switch.scala 41:38:@26358.4]
  wire  _T_65201; // @[Switch.scala 41:52:@26360.4]
  wire  output_22_29; // @[Switch.scala 41:38:@26361.4]
  wire  _T_65204; // @[Switch.scala 41:52:@26363.4]
  wire  output_22_30; // @[Switch.scala 41:38:@26364.4]
  wire  _T_65207; // @[Switch.scala 41:52:@26366.4]
  wire  output_22_31; // @[Switch.scala 41:38:@26367.4]
  wire  _T_65210; // @[Switch.scala 41:52:@26369.4]
  wire  output_22_32; // @[Switch.scala 41:38:@26370.4]
  wire  _T_65213; // @[Switch.scala 41:52:@26372.4]
  wire  output_22_33; // @[Switch.scala 41:38:@26373.4]
  wire  _T_65216; // @[Switch.scala 41:52:@26375.4]
  wire  output_22_34; // @[Switch.scala 41:38:@26376.4]
  wire  _T_65219; // @[Switch.scala 41:52:@26378.4]
  wire  output_22_35; // @[Switch.scala 41:38:@26379.4]
  wire  _T_65222; // @[Switch.scala 41:52:@26381.4]
  wire  output_22_36; // @[Switch.scala 41:38:@26382.4]
  wire  _T_65225; // @[Switch.scala 41:52:@26384.4]
  wire  output_22_37; // @[Switch.scala 41:38:@26385.4]
  wire  _T_65228; // @[Switch.scala 41:52:@26387.4]
  wire  output_22_38; // @[Switch.scala 41:38:@26388.4]
  wire  _T_65231; // @[Switch.scala 41:52:@26390.4]
  wire  output_22_39; // @[Switch.scala 41:38:@26391.4]
  wire  _T_65234; // @[Switch.scala 41:52:@26393.4]
  wire  output_22_40; // @[Switch.scala 41:38:@26394.4]
  wire  _T_65237; // @[Switch.scala 41:52:@26396.4]
  wire  output_22_41; // @[Switch.scala 41:38:@26397.4]
  wire  _T_65240; // @[Switch.scala 41:52:@26399.4]
  wire  output_22_42; // @[Switch.scala 41:38:@26400.4]
  wire  _T_65243; // @[Switch.scala 41:52:@26402.4]
  wire  output_22_43; // @[Switch.scala 41:38:@26403.4]
  wire  _T_65246; // @[Switch.scala 41:52:@26405.4]
  wire  output_22_44; // @[Switch.scala 41:38:@26406.4]
  wire  _T_65249; // @[Switch.scala 41:52:@26408.4]
  wire  output_22_45; // @[Switch.scala 41:38:@26409.4]
  wire  _T_65252; // @[Switch.scala 41:52:@26411.4]
  wire  output_22_46; // @[Switch.scala 41:38:@26412.4]
  wire  _T_65255; // @[Switch.scala 41:52:@26414.4]
  wire  output_22_47; // @[Switch.scala 41:38:@26415.4]
  wire  _T_65258; // @[Switch.scala 41:52:@26417.4]
  wire  output_22_48; // @[Switch.scala 41:38:@26418.4]
  wire  _T_65261; // @[Switch.scala 41:52:@26420.4]
  wire  output_22_49; // @[Switch.scala 41:38:@26421.4]
  wire  _T_65264; // @[Switch.scala 41:52:@26423.4]
  wire  output_22_50; // @[Switch.scala 41:38:@26424.4]
  wire  _T_65267; // @[Switch.scala 41:52:@26426.4]
  wire  output_22_51; // @[Switch.scala 41:38:@26427.4]
  wire  _T_65270; // @[Switch.scala 41:52:@26429.4]
  wire  output_22_52; // @[Switch.scala 41:38:@26430.4]
  wire  _T_65273; // @[Switch.scala 41:52:@26432.4]
  wire  output_22_53; // @[Switch.scala 41:38:@26433.4]
  wire  _T_65276; // @[Switch.scala 41:52:@26435.4]
  wire  output_22_54; // @[Switch.scala 41:38:@26436.4]
  wire  _T_65279; // @[Switch.scala 41:52:@26438.4]
  wire  output_22_55; // @[Switch.scala 41:38:@26439.4]
  wire  _T_65282; // @[Switch.scala 41:52:@26441.4]
  wire  output_22_56; // @[Switch.scala 41:38:@26442.4]
  wire  _T_65285; // @[Switch.scala 41:52:@26444.4]
  wire  output_22_57; // @[Switch.scala 41:38:@26445.4]
  wire  _T_65288; // @[Switch.scala 41:52:@26447.4]
  wire  output_22_58; // @[Switch.scala 41:38:@26448.4]
  wire  _T_65291; // @[Switch.scala 41:52:@26450.4]
  wire  output_22_59; // @[Switch.scala 41:38:@26451.4]
  wire  _T_65294; // @[Switch.scala 41:52:@26453.4]
  wire  output_22_60; // @[Switch.scala 41:38:@26454.4]
  wire  _T_65297; // @[Switch.scala 41:52:@26456.4]
  wire  output_22_61; // @[Switch.scala 41:38:@26457.4]
  wire  _T_65300; // @[Switch.scala 41:52:@26459.4]
  wire  output_22_62; // @[Switch.scala 41:38:@26460.4]
  wire  _T_65303; // @[Switch.scala 41:52:@26462.4]
  wire  output_22_63; // @[Switch.scala 41:38:@26463.4]
  wire [7:0] _T_65311; // @[Switch.scala 43:31:@26471.4]
  wire [15:0] _T_65319; // @[Switch.scala 43:31:@26479.4]
  wire [7:0] _T_65326; // @[Switch.scala 43:31:@26486.4]
  wire [31:0] _T_65335; // @[Switch.scala 43:31:@26495.4]
  wire [7:0] _T_65342; // @[Switch.scala 43:31:@26502.4]
  wire [15:0] _T_65350; // @[Switch.scala 43:31:@26510.4]
  wire [7:0] _T_65357; // @[Switch.scala 43:31:@26517.4]
  wire [31:0] _T_65366; // @[Switch.scala 43:31:@26526.4]
  wire [63:0] _T_65367; // @[Switch.scala 43:31:@26527.4]
  wire  _T_65371; // @[Switch.scala 41:52:@26530.4]
  wire  output_23_0; // @[Switch.scala 41:38:@26531.4]
  wire  _T_65374; // @[Switch.scala 41:52:@26533.4]
  wire  output_23_1; // @[Switch.scala 41:38:@26534.4]
  wire  _T_65377; // @[Switch.scala 41:52:@26536.4]
  wire  output_23_2; // @[Switch.scala 41:38:@26537.4]
  wire  _T_65380; // @[Switch.scala 41:52:@26539.4]
  wire  output_23_3; // @[Switch.scala 41:38:@26540.4]
  wire  _T_65383; // @[Switch.scala 41:52:@26542.4]
  wire  output_23_4; // @[Switch.scala 41:38:@26543.4]
  wire  _T_65386; // @[Switch.scala 41:52:@26545.4]
  wire  output_23_5; // @[Switch.scala 41:38:@26546.4]
  wire  _T_65389; // @[Switch.scala 41:52:@26548.4]
  wire  output_23_6; // @[Switch.scala 41:38:@26549.4]
  wire  _T_65392; // @[Switch.scala 41:52:@26551.4]
  wire  output_23_7; // @[Switch.scala 41:38:@26552.4]
  wire  _T_65395; // @[Switch.scala 41:52:@26554.4]
  wire  output_23_8; // @[Switch.scala 41:38:@26555.4]
  wire  _T_65398; // @[Switch.scala 41:52:@26557.4]
  wire  output_23_9; // @[Switch.scala 41:38:@26558.4]
  wire  _T_65401; // @[Switch.scala 41:52:@26560.4]
  wire  output_23_10; // @[Switch.scala 41:38:@26561.4]
  wire  _T_65404; // @[Switch.scala 41:52:@26563.4]
  wire  output_23_11; // @[Switch.scala 41:38:@26564.4]
  wire  _T_65407; // @[Switch.scala 41:52:@26566.4]
  wire  output_23_12; // @[Switch.scala 41:38:@26567.4]
  wire  _T_65410; // @[Switch.scala 41:52:@26569.4]
  wire  output_23_13; // @[Switch.scala 41:38:@26570.4]
  wire  _T_65413; // @[Switch.scala 41:52:@26572.4]
  wire  output_23_14; // @[Switch.scala 41:38:@26573.4]
  wire  _T_65416; // @[Switch.scala 41:52:@26575.4]
  wire  output_23_15; // @[Switch.scala 41:38:@26576.4]
  wire  _T_65419; // @[Switch.scala 41:52:@26578.4]
  wire  output_23_16; // @[Switch.scala 41:38:@26579.4]
  wire  _T_65422; // @[Switch.scala 41:52:@26581.4]
  wire  output_23_17; // @[Switch.scala 41:38:@26582.4]
  wire  _T_65425; // @[Switch.scala 41:52:@26584.4]
  wire  output_23_18; // @[Switch.scala 41:38:@26585.4]
  wire  _T_65428; // @[Switch.scala 41:52:@26587.4]
  wire  output_23_19; // @[Switch.scala 41:38:@26588.4]
  wire  _T_65431; // @[Switch.scala 41:52:@26590.4]
  wire  output_23_20; // @[Switch.scala 41:38:@26591.4]
  wire  _T_65434; // @[Switch.scala 41:52:@26593.4]
  wire  output_23_21; // @[Switch.scala 41:38:@26594.4]
  wire  _T_65437; // @[Switch.scala 41:52:@26596.4]
  wire  output_23_22; // @[Switch.scala 41:38:@26597.4]
  wire  _T_65440; // @[Switch.scala 41:52:@26599.4]
  wire  output_23_23; // @[Switch.scala 41:38:@26600.4]
  wire  _T_65443; // @[Switch.scala 41:52:@26602.4]
  wire  output_23_24; // @[Switch.scala 41:38:@26603.4]
  wire  _T_65446; // @[Switch.scala 41:52:@26605.4]
  wire  output_23_25; // @[Switch.scala 41:38:@26606.4]
  wire  _T_65449; // @[Switch.scala 41:52:@26608.4]
  wire  output_23_26; // @[Switch.scala 41:38:@26609.4]
  wire  _T_65452; // @[Switch.scala 41:52:@26611.4]
  wire  output_23_27; // @[Switch.scala 41:38:@26612.4]
  wire  _T_65455; // @[Switch.scala 41:52:@26614.4]
  wire  output_23_28; // @[Switch.scala 41:38:@26615.4]
  wire  _T_65458; // @[Switch.scala 41:52:@26617.4]
  wire  output_23_29; // @[Switch.scala 41:38:@26618.4]
  wire  _T_65461; // @[Switch.scala 41:52:@26620.4]
  wire  output_23_30; // @[Switch.scala 41:38:@26621.4]
  wire  _T_65464; // @[Switch.scala 41:52:@26623.4]
  wire  output_23_31; // @[Switch.scala 41:38:@26624.4]
  wire  _T_65467; // @[Switch.scala 41:52:@26626.4]
  wire  output_23_32; // @[Switch.scala 41:38:@26627.4]
  wire  _T_65470; // @[Switch.scala 41:52:@26629.4]
  wire  output_23_33; // @[Switch.scala 41:38:@26630.4]
  wire  _T_65473; // @[Switch.scala 41:52:@26632.4]
  wire  output_23_34; // @[Switch.scala 41:38:@26633.4]
  wire  _T_65476; // @[Switch.scala 41:52:@26635.4]
  wire  output_23_35; // @[Switch.scala 41:38:@26636.4]
  wire  _T_65479; // @[Switch.scala 41:52:@26638.4]
  wire  output_23_36; // @[Switch.scala 41:38:@26639.4]
  wire  _T_65482; // @[Switch.scala 41:52:@26641.4]
  wire  output_23_37; // @[Switch.scala 41:38:@26642.4]
  wire  _T_65485; // @[Switch.scala 41:52:@26644.4]
  wire  output_23_38; // @[Switch.scala 41:38:@26645.4]
  wire  _T_65488; // @[Switch.scala 41:52:@26647.4]
  wire  output_23_39; // @[Switch.scala 41:38:@26648.4]
  wire  _T_65491; // @[Switch.scala 41:52:@26650.4]
  wire  output_23_40; // @[Switch.scala 41:38:@26651.4]
  wire  _T_65494; // @[Switch.scala 41:52:@26653.4]
  wire  output_23_41; // @[Switch.scala 41:38:@26654.4]
  wire  _T_65497; // @[Switch.scala 41:52:@26656.4]
  wire  output_23_42; // @[Switch.scala 41:38:@26657.4]
  wire  _T_65500; // @[Switch.scala 41:52:@26659.4]
  wire  output_23_43; // @[Switch.scala 41:38:@26660.4]
  wire  _T_65503; // @[Switch.scala 41:52:@26662.4]
  wire  output_23_44; // @[Switch.scala 41:38:@26663.4]
  wire  _T_65506; // @[Switch.scala 41:52:@26665.4]
  wire  output_23_45; // @[Switch.scala 41:38:@26666.4]
  wire  _T_65509; // @[Switch.scala 41:52:@26668.4]
  wire  output_23_46; // @[Switch.scala 41:38:@26669.4]
  wire  _T_65512; // @[Switch.scala 41:52:@26671.4]
  wire  output_23_47; // @[Switch.scala 41:38:@26672.4]
  wire  _T_65515; // @[Switch.scala 41:52:@26674.4]
  wire  output_23_48; // @[Switch.scala 41:38:@26675.4]
  wire  _T_65518; // @[Switch.scala 41:52:@26677.4]
  wire  output_23_49; // @[Switch.scala 41:38:@26678.4]
  wire  _T_65521; // @[Switch.scala 41:52:@26680.4]
  wire  output_23_50; // @[Switch.scala 41:38:@26681.4]
  wire  _T_65524; // @[Switch.scala 41:52:@26683.4]
  wire  output_23_51; // @[Switch.scala 41:38:@26684.4]
  wire  _T_65527; // @[Switch.scala 41:52:@26686.4]
  wire  output_23_52; // @[Switch.scala 41:38:@26687.4]
  wire  _T_65530; // @[Switch.scala 41:52:@26689.4]
  wire  output_23_53; // @[Switch.scala 41:38:@26690.4]
  wire  _T_65533; // @[Switch.scala 41:52:@26692.4]
  wire  output_23_54; // @[Switch.scala 41:38:@26693.4]
  wire  _T_65536; // @[Switch.scala 41:52:@26695.4]
  wire  output_23_55; // @[Switch.scala 41:38:@26696.4]
  wire  _T_65539; // @[Switch.scala 41:52:@26698.4]
  wire  output_23_56; // @[Switch.scala 41:38:@26699.4]
  wire  _T_65542; // @[Switch.scala 41:52:@26701.4]
  wire  output_23_57; // @[Switch.scala 41:38:@26702.4]
  wire  _T_65545; // @[Switch.scala 41:52:@26704.4]
  wire  output_23_58; // @[Switch.scala 41:38:@26705.4]
  wire  _T_65548; // @[Switch.scala 41:52:@26707.4]
  wire  output_23_59; // @[Switch.scala 41:38:@26708.4]
  wire  _T_65551; // @[Switch.scala 41:52:@26710.4]
  wire  output_23_60; // @[Switch.scala 41:38:@26711.4]
  wire  _T_65554; // @[Switch.scala 41:52:@26713.4]
  wire  output_23_61; // @[Switch.scala 41:38:@26714.4]
  wire  _T_65557; // @[Switch.scala 41:52:@26716.4]
  wire  output_23_62; // @[Switch.scala 41:38:@26717.4]
  wire  _T_65560; // @[Switch.scala 41:52:@26719.4]
  wire  output_23_63; // @[Switch.scala 41:38:@26720.4]
  wire [7:0] _T_65568; // @[Switch.scala 43:31:@26728.4]
  wire [15:0] _T_65576; // @[Switch.scala 43:31:@26736.4]
  wire [7:0] _T_65583; // @[Switch.scala 43:31:@26743.4]
  wire [31:0] _T_65592; // @[Switch.scala 43:31:@26752.4]
  wire [7:0] _T_65599; // @[Switch.scala 43:31:@26759.4]
  wire [15:0] _T_65607; // @[Switch.scala 43:31:@26767.4]
  wire [7:0] _T_65614; // @[Switch.scala 43:31:@26774.4]
  wire [31:0] _T_65623; // @[Switch.scala 43:31:@26783.4]
  wire [63:0] _T_65624; // @[Switch.scala 43:31:@26784.4]
  wire  _T_65628; // @[Switch.scala 41:52:@26787.4]
  wire  output_24_0; // @[Switch.scala 41:38:@26788.4]
  wire  _T_65631; // @[Switch.scala 41:52:@26790.4]
  wire  output_24_1; // @[Switch.scala 41:38:@26791.4]
  wire  _T_65634; // @[Switch.scala 41:52:@26793.4]
  wire  output_24_2; // @[Switch.scala 41:38:@26794.4]
  wire  _T_65637; // @[Switch.scala 41:52:@26796.4]
  wire  output_24_3; // @[Switch.scala 41:38:@26797.4]
  wire  _T_65640; // @[Switch.scala 41:52:@26799.4]
  wire  output_24_4; // @[Switch.scala 41:38:@26800.4]
  wire  _T_65643; // @[Switch.scala 41:52:@26802.4]
  wire  output_24_5; // @[Switch.scala 41:38:@26803.4]
  wire  _T_65646; // @[Switch.scala 41:52:@26805.4]
  wire  output_24_6; // @[Switch.scala 41:38:@26806.4]
  wire  _T_65649; // @[Switch.scala 41:52:@26808.4]
  wire  output_24_7; // @[Switch.scala 41:38:@26809.4]
  wire  _T_65652; // @[Switch.scala 41:52:@26811.4]
  wire  output_24_8; // @[Switch.scala 41:38:@26812.4]
  wire  _T_65655; // @[Switch.scala 41:52:@26814.4]
  wire  output_24_9; // @[Switch.scala 41:38:@26815.4]
  wire  _T_65658; // @[Switch.scala 41:52:@26817.4]
  wire  output_24_10; // @[Switch.scala 41:38:@26818.4]
  wire  _T_65661; // @[Switch.scala 41:52:@26820.4]
  wire  output_24_11; // @[Switch.scala 41:38:@26821.4]
  wire  _T_65664; // @[Switch.scala 41:52:@26823.4]
  wire  output_24_12; // @[Switch.scala 41:38:@26824.4]
  wire  _T_65667; // @[Switch.scala 41:52:@26826.4]
  wire  output_24_13; // @[Switch.scala 41:38:@26827.4]
  wire  _T_65670; // @[Switch.scala 41:52:@26829.4]
  wire  output_24_14; // @[Switch.scala 41:38:@26830.4]
  wire  _T_65673; // @[Switch.scala 41:52:@26832.4]
  wire  output_24_15; // @[Switch.scala 41:38:@26833.4]
  wire  _T_65676; // @[Switch.scala 41:52:@26835.4]
  wire  output_24_16; // @[Switch.scala 41:38:@26836.4]
  wire  _T_65679; // @[Switch.scala 41:52:@26838.4]
  wire  output_24_17; // @[Switch.scala 41:38:@26839.4]
  wire  _T_65682; // @[Switch.scala 41:52:@26841.4]
  wire  output_24_18; // @[Switch.scala 41:38:@26842.4]
  wire  _T_65685; // @[Switch.scala 41:52:@26844.4]
  wire  output_24_19; // @[Switch.scala 41:38:@26845.4]
  wire  _T_65688; // @[Switch.scala 41:52:@26847.4]
  wire  output_24_20; // @[Switch.scala 41:38:@26848.4]
  wire  _T_65691; // @[Switch.scala 41:52:@26850.4]
  wire  output_24_21; // @[Switch.scala 41:38:@26851.4]
  wire  _T_65694; // @[Switch.scala 41:52:@26853.4]
  wire  output_24_22; // @[Switch.scala 41:38:@26854.4]
  wire  _T_65697; // @[Switch.scala 41:52:@26856.4]
  wire  output_24_23; // @[Switch.scala 41:38:@26857.4]
  wire  _T_65700; // @[Switch.scala 41:52:@26859.4]
  wire  output_24_24; // @[Switch.scala 41:38:@26860.4]
  wire  _T_65703; // @[Switch.scala 41:52:@26862.4]
  wire  output_24_25; // @[Switch.scala 41:38:@26863.4]
  wire  _T_65706; // @[Switch.scala 41:52:@26865.4]
  wire  output_24_26; // @[Switch.scala 41:38:@26866.4]
  wire  _T_65709; // @[Switch.scala 41:52:@26868.4]
  wire  output_24_27; // @[Switch.scala 41:38:@26869.4]
  wire  _T_65712; // @[Switch.scala 41:52:@26871.4]
  wire  output_24_28; // @[Switch.scala 41:38:@26872.4]
  wire  _T_65715; // @[Switch.scala 41:52:@26874.4]
  wire  output_24_29; // @[Switch.scala 41:38:@26875.4]
  wire  _T_65718; // @[Switch.scala 41:52:@26877.4]
  wire  output_24_30; // @[Switch.scala 41:38:@26878.4]
  wire  _T_65721; // @[Switch.scala 41:52:@26880.4]
  wire  output_24_31; // @[Switch.scala 41:38:@26881.4]
  wire  _T_65724; // @[Switch.scala 41:52:@26883.4]
  wire  output_24_32; // @[Switch.scala 41:38:@26884.4]
  wire  _T_65727; // @[Switch.scala 41:52:@26886.4]
  wire  output_24_33; // @[Switch.scala 41:38:@26887.4]
  wire  _T_65730; // @[Switch.scala 41:52:@26889.4]
  wire  output_24_34; // @[Switch.scala 41:38:@26890.4]
  wire  _T_65733; // @[Switch.scala 41:52:@26892.4]
  wire  output_24_35; // @[Switch.scala 41:38:@26893.4]
  wire  _T_65736; // @[Switch.scala 41:52:@26895.4]
  wire  output_24_36; // @[Switch.scala 41:38:@26896.4]
  wire  _T_65739; // @[Switch.scala 41:52:@26898.4]
  wire  output_24_37; // @[Switch.scala 41:38:@26899.4]
  wire  _T_65742; // @[Switch.scala 41:52:@26901.4]
  wire  output_24_38; // @[Switch.scala 41:38:@26902.4]
  wire  _T_65745; // @[Switch.scala 41:52:@26904.4]
  wire  output_24_39; // @[Switch.scala 41:38:@26905.4]
  wire  _T_65748; // @[Switch.scala 41:52:@26907.4]
  wire  output_24_40; // @[Switch.scala 41:38:@26908.4]
  wire  _T_65751; // @[Switch.scala 41:52:@26910.4]
  wire  output_24_41; // @[Switch.scala 41:38:@26911.4]
  wire  _T_65754; // @[Switch.scala 41:52:@26913.4]
  wire  output_24_42; // @[Switch.scala 41:38:@26914.4]
  wire  _T_65757; // @[Switch.scala 41:52:@26916.4]
  wire  output_24_43; // @[Switch.scala 41:38:@26917.4]
  wire  _T_65760; // @[Switch.scala 41:52:@26919.4]
  wire  output_24_44; // @[Switch.scala 41:38:@26920.4]
  wire  _T_65763; // @[Switch.scala 41:52:@26922.4]
  wire  output_24_45; // @[Switch.scala 41:38:@26923.4]
  wire  _T_65766; // @[Switch.scala 41:52:@26925.4]
  wire  output_24_46; // @[Switch.scala 41:38:@26926.4]
  wire  _T_65769; // @[Switch.scala 41:52:@26928.4]
  wire  output_24_47; // @[Switch.scala 41:38:@26929.4]
  wire  _T_65772; // @[Switch.scala 41:52:@26931.4]
  wire  output_24_48; // @[Switch.scala 41:38:@26932.4]
  wire  _T_65775; // @[Switch.scala 41:52:@26934.4]
  wire  output_24_49; // @[Switch.scala 41:38:@26935.4]
  wire  _T_65778; // @[Switch.scala 41:52:@26937.4]
  wire  output_24_50; // @[Switch.scala 41:38:@26938.4]
  wire  _T_65781; // @[Switch.scala 41:52:@26940.4]
  wire  output_24_51; // @[Switch.scala 41:38:@26941.4]
  wire  _T_65784; // @[Switch.scala 41:52:@26943.4]
  wire  output_24_52; // @[Switch.scala 41:38:@26944.4]
  wire  _T_65787; // @[Switch.scala 41:52:@26946.4]
  wire  output_24_53; // @[Switch.scala 41:38:@26947.4]
  wire  _T_65790; // @[Switch.scala 41:52:@26949.4]
  wire  output_24_54; // @[Switch.scala 41:38:@26950.4]
  wire  _T_65793; // @[Switch.scala 41:52:@26952.4]
  wire  output_24_55; // @[Switch.scala 41:38:@26953.4]
  wire  _T_65796; // @[Switch.scala 41:52:@26955.4]
  wire  output_24_56; // @[Switch.scala 41:38:@26956.4]
  wire  _T_65799; // @[Switch.scala 41:52:@26958.4]
  wire  output_24_57; // @[Switch.scala 41:38:@26959.4]
  wire  _T_65802; // @[Switch.scala 41:52:@26961.4]
  wire  output_24_58; // @[Switch.scala 41:38:@26962.4]
  wire  _T_65805; // @[Switch.scala 41:52:@26964.4]
  wire  output_24_59; // @[Switch.scala 41:38:@26965.4]
  wire  _T_65808; // @[Switch.scala 41:52:@26967.4]
  wire  output_24_60; // @[Switch.scala 41:38:@26968.4]
  wire  _T_65811; // @[Switch.scala 41:52:@26970.4]
  wire  output_24_61; // @[Switch.scala 41:38:@26971.4]
  wire  _T_65814; // @[Switch.scala 41:52:@26973.4]
  wire  output_24_62; // @[Switch.scala 41:38:@26974.4]
  wire  _T_65817; // @[Switch.scala 41:52:@26976.4]
  wire  output_24_63; // @[Switch.scala 41:38:@26977.4]
  wire [7:0] _T_65825; // @[Switch.scala 43:31:@26985.4]
  wire [15:0] _T_65833; // @[Switch.scala 43:31:@26993.4]
  wire [7:0] _T_65840; // @[Switch.scala 43:31:@27000.4]
  wire [31:0] _T_65849; // @[Switch.scala 43:31:@27009.4]
  wire [7:0] _T_65856; // @[Switch.scala 43:31:@27016.4]
  wire [15:0] _T_65864; // @[Switch.scala 43:31:@27024.4]
  wire [7:0] _T_65871; // @[Switch.scala 43:31:@27031.4]
  wire [31:0] _T_65880; // @[Switch.scala 43:31:@27040.4]
  wire [63:0] _T_65881; // @[Switch.scala 43:31:@27041.4]
  wire  _T_65885; // @[Switch.scala 41:52:@27044.4]
  wire  output_25_0; // @[Switch.scala 41:38:@27045.4]
  wire  _T_65888; // @[Switch.scala 41:52:@27047.4]
  wire  output_25_1; // @[Switch.scala 41:38:@27048.4]
  wire  _T_65891; // @[Switch.scala 41:52:@27050.4]
  wire  output_25_2; // @[Switch.scala 41:38:@27051.4]
  wire  _T_65894; // @[Switch.scala 41:52:@27053.4]
  wire  output_25_3; // @[Switch.scala 41:38:@27054.4]
  wire  _T_65897; // @[Switch.scala 41:52:@27056.4]
  wire  output_25_4; // @[Switch.scala 41:38:@27057.4]
  wire  _T_65900; // @[Switch.scala 41:52:@27059.4]
  wire  output_25_5; // @[Switch.scala 41:38:@27060.4]
  wire  _T_65903; // @[Switch.scala 41:52:@27062.4]
  wire  output_25_6; // @[Switch.scala 41:38:@27063.4]
  wire  _T_65906; // @[Switch.scala 41:52:@27065.4]
  wire  output_25_7; // @[Switch.scala 41:38:@27066.4]
  wire  _T_65909; // @[Switch.scala 41:52:@27068.4]
  wire  output_25_8; // @[Switch.scala 41:38:@27069.4]
  wire  _T_65912; // @[Switch.scala 41:52:@27071.4]
  wire  output_25_9; // @[Switch.scala 41:38:@27072.4]
  wire  _T_65915; // @[Switch.scala 41:52:@27074.4]
  wire  output_25_10; // @[Switch.scala 41:38:@27075.4]
  wire  _T_65918; // @[Switch.scala 41:52:@27077.4]
  wire  output_25_11; // @[Switch.scala 41:38:@27078.4]
  wire  _T_65921; // @[Switch.scala 41:52:@27080.4]
  wire  output_25_12; // @[Switch.scala 41:38:@27081.4]
  wire  _T_65924; // @[Switch.scala 41:52:@27083.4]
  wire  output_25_13; // @[Switch.scala 41:38:@27084.4]
  wire  _T_65927; // @[Switch.scala 41:52:@27086.4]
  wire  output_25_14; // @[Switch.scala 41:38:@27087.4]
  wire  _T_65930; // @[Switch.scala 41:52:@27089.4]
  wire  output_25_15; // @[Switch.scala 41:38:@27090.4]
  wire  _T_65933; // @[Switch.scala 41:52:@27092.4]
  wire  output_25_16; // @[Switch.scala 41:38:@27093.4]
  wire  _T_65936; // @[Switch.scala 41:52:@27095.4]
  wire  output_25_17; // @[Switch.scala 41:38:@27096.4]
  wire  _T_65939; // @[Switch.scala 41:52:@27098.4]
  wire  output_25_18; // @[Switch.scala 41:38:@27099.4]
  wire  _T_65942; // @[Switch.scala 41:52:@27101.4]
  wire  output_25_19; // @[Switch.scala 41:38:@27102.4]
  wire  _T_65945; // @[Switch.scala 41:52:@27104.4]
  wire  output_25_20; // @[Switch.scala 41:38:@27105.4]
  wire  _T_65948; // @[Switch.scala 41:52:@27107.4]
  wire  output_25_21; // @[Switch.scala 41:38:@27108.4]
  wire  _T_65951; // @[Switch.scala 41:52:@27110.4]
  wire  output_25_22; // @[Switch.scala 41:38:@27111.4]
  wire  _T_65954; // @[Switch.scala 41:52:@27113.4]
  wire  output_25_23; // @[Switch.scala 41:38:@27114.4]
  wire  _T_65957; // @[Switch.scala 41:52:@27116.4]
  wire  output_25_24; // @[Switch.scala 41:38:@27117.4]
  wire  _T_65960; // @[Switch.scala 41:52:@27119.4]
  wire  output_25_25; // @[Switch.scala 41:38:@27120.4]
  wire  _T_65963; // @[Switch.scala 41:52:@27122.4]
  wire  output_25_26; // @[Switch.scala 41:38:@27123.4]
  wire  _T_65966; // @[Switch.scala 41:52:@27125.4]
  wire  output_25_27; // @[Switch.scala 41:38:@27126.4]
  wire  _T_65969; // @[Switch.scala 41:52:@27128.4]
  wire  output_25_28; // @[Switch.scala 41:38:@27129.4]
  wire  _T_65972; // @[Switch.scala 41:52:@27131.4]
  wire  output_25_29; // @[Switch.scala 41:38:@27132.4]
  wire  _T_65975; // @[Switch.scala 41:52:@27134.4]
  wire  output_25_30; // @[Switch.scala 41:38:@27135.4]
  wire  _T_65978; // @[Switch.scala 41:52:@27137.4]
  wire  output_25_31; // @[Switch.scala 41:38:@27138.4]
  wire  _T_65981; // @[Switch.scala 41:52:@27140.4]
  wire  output_25_32; // @[Switch.scala 41:38:@27141.4]
  wire  _T_65984; // @[Switch.scala 41:52:@27143.4]
  wire  output_25_33; // @[Switch.scala 41:38:@27144.4]
  wire  _T_65987; // @[Switch.scala 41:52:@27146.4]
  wire  output_25_34; // @[Switch.scala 41:38:@27147.4]
  wire  _T_65990; // @[Switch.scala 41:52:@27149.4]
  wire  output_25_35; // @[Switch.scala 41:38:@27150.4]
  wire  _T_65993; // @[Switch.scala 41:52:@27152.4]
  wire  output_25_36; // @[Switch.scala 41:38:@27153.4]
  wire  _T_65996; // @[Switch.scala 41:52:@27155.4]
  wire  output_25_37; // @[Switch.scala 41:38:@27156.4]
  wire  _T_65999; // @[Switch.scala 41:52:@27158.4]
  wire  output_25_38; // @[Switch.scala 41:38:@27159.4]
  wire  _T_66002; // @[Switch.scala 41:52:@27161.4]
  wire  output_25_39; // @[Switch.scala 41:38:@27162.4]
  wire  _T_66005; // @[Switch.scala 41:52:@27164.4]
  wire  output_25_40; // @[Switch.scala 41:38:@27165.4]
  wire  _T_66008; // @[Switch.scala 41:52:@27167.4]
  wire  output_25_41; // @[Switch.scala 41:38:@27168.4]
  wire  _T_66011; // @[Switch.scala 41:52:@27170.4]
  wire  output_25_42; // @[Switch.scala 41:38:@27171.4]
  wire  _T_66014; // @[Switch.scala 41:52:@27173.4]
  wire  output_25_43; // @[Switch.scala 41:38:@27174.4]
  wire  _T_66017; // @[Switch.scala 41:52:@27176.4]
  wire  output_25_44; // @[Switch.scala 41:38:@27177.4]
  wire  _T_66020; // @[Switch.scala 41:52:@27179.4]
  wire  output_25_45; // @[Switch.scala 41:38:@27180.4]
  wire  _T_66023; // @[Switch.scala 41:52:@27182.4]
  wire  output_25_46; // @[Switch.scala 41:38:@27183.4]
  wire  _T_66026; // @[Switch.scala 41:52:@27185.4]
  wire  output_25_47; // @[Switch.scala 41:38:@27186.4]
  wire  _T_66029; // @[Switch.scala 41:52:@27188.4]
  wire  output_25_48; // @[Switch.scala 41:38:@27189.4]
  wire  _T_66032; // @[Switch.scala 41:52:@27191.4]
  wire  output_25_49; // @[Switch.scala 41:38:@27192.4]
  wire  _T_66035; // @[Switch.scala 41:52:@27194.4]
  wire  output_25_50; // @[Switch.scala 41:38:@27195.4]
  wire  _T_66038; // @[Switch.scala 41:52:@27197.4]
  wire  output_25_51; // @[Switch.scala 41:38:@27198.4]
  wire  _T_66041; // @[Switch.scala 41:52:@27200.4]
  wire  output_25_52; // @[Switch.scala 41:38:@27201.4]
  wire  _T_66044; // @[Switch.scala 41:52:@27203.4]
  wire  output_25_53; // @[Switch.scala 41:38:@27204.4]
  wire  _T_66047; // @[Switch.scala 41:52:@27206.4]
  wire  output_25_54; // @[Switch.scala 41:38:@27207.4]
  wire  _T_66050; // @[Switch.scala 41:52:@27209.4]
  wire  output_25_55; // @[Switch.scala 41:38:@27210.4]
  wire  _T_66053; // @[Switch.scala 41:52:@27212.4]
  wire  output_25_56; // @[Switch.scala 41:38:@27213.4]
  wire  _T_66056; // @[Switch.scala 41:52:@27215.4]
  wire  output_25_57; // @[Switch.scala 41:38:@27216.4]
  wire  _T_66059; // @[Switch.scala 41:52:@27218.4]
  wire  output_25_58; // @[Switch.scala 41:38:@27219.4]
  wire  _T_66062; // @[Switch.scala 41:52:@27221.4]
  wire  output_25_59; // @[Switch.scala 41:38:@27222.4]
  wire  _T_66065; // @[Switch.scala 41:52:@27224.4]
  wire  output_25_60; // @[Switch.scala 41:38:@27225.4]
  wire  _T_66068; // @[Switch.scala 41:52:@27227.4]
  wire  output_25_61; // @[Switch.scala 41:38:@27228.4]
  wire  _T_66071; // @[Switch.scala 41:52:@27230.4]
  wire  output_25_62; // @[Switch.scala 41:38:@27231.4]
  wire  _T_66074; // @[Switch.scala 41:52:@27233.4]
  wire  output_25_63; // @[Switch.scala 41:38:@27234.4]
  wire [7:0] _T_66082; // @[Switch.scala 43:31:@27242.4]
  wire [15:0] _T_66090; // @[Switch.scala 43:31:@27250.4]
  wire [7:0] _T_66097; // @[Switch.scala 43:31:@27257.4]
  wire [31:0] _T_66106; // @[Switch.scala 43:31:@27266.4]
  wire [7:0] _T_66113; // @[Switch.scala 43:31:@27273.4]
  wire [15:0] _T_66121; // @[Switch.scala 43:31:@27281.4]
  wire [7:0] _T_66128; // @[Switch.scala 43:31:@27288.4]
  wire [31:0] _T_66137; // @[Switch.scala 43:31:@27297.4]
  wire [63:0] _T_66138; // @[Switch.scala 43:31:@27298.4]
  wire  _T_66142; // @[Switch.scala 41:52:@27301.4]
  wire  output_26_0; // @[Switch.scala 41:38:@27302.4]
  wire  _T_66145; // @[Switch.scala 41:52:@27304.4]
  wire  output_26_1; // @[Switch.scala 41:38:@27305.4]
  wire  _T_66148; // @[Switch.scala 41:52:@27307.4]
  wire  output_26_2; // @[Switch.scala 41:38:@27308.4]
  wire  _T_66151; // @[Switch.scala 41:52:@27310.4]
  wire  output_26_3; // @[Switch.scala 41:38:@27311.4]
  wire  _T_66154; // @[Switch.scala 41:52:@27313.4]
  wire  output_26_4; // @[Switch.scala 41:38:@27314.4]
  wire  _T_66157; // @[Switch.scala 41:52:@27316.4]
  wire  output_26_5; // @[Switch.scala 41:38:@27317.4]
  wire  _T_66160; // @[Switch.scala 41:52:@27319.4]
  wire  output_26_6; // @[Switch.scala 41:38:@27320.4]
  wire  _T_66163; // @[Switch.scala 41:52:@27322.4]
  wire  output_26_7; // @[Switch.scala 41:38:@27323.4]
  wire  _T_66166; // @[Switch.scala 41:52:@27325.4]
  wire  output_26_8; // @[Switch.scala 41:38:@27326.4]
  wire  _T_66169; // @[Switch.scala 41:52:@27328.4]
  wire  output_26_9; // @[Switch.scala 41:38:@27329.4]
  wire  _T_66172; // @[Switch.scala 41:52:@27331.4]
  wire  output_26_10; // @[Switch.scala 41:38:@27332.4]
  wire  _T_66175; // @[Switch.scala 41:52:@27334.4]
  wire  output_26_11; // @[Switch.scala 41:38:@27335.4]
  wire  _T_66178; // @[Switch.scala 41:52:@27337.4]
  wire  output_26_12; // @[Switch.scala 41:38:@27338.4]
  wire  _T_66181; // @[Switch.scala 41:52:@27340.4]
  wire  output_26_13; // @[Switch.scala 41:38:@27341.4]
  wire  _T_66184; // @[Switch.scala 41:52:@27343.4]
  wire  output_26_14; // @[Switch.scala 41:38:@27344.4]
  wire  _T_66187; // @[Switch.scala 41:52:@27346.4]
  wire  output_26_15; // @[Switch.scala 41:38:@27347.4]
  wire  _T_66190; // @[Switch.scala 41:52:@27349.4]
  wire  output_26_16; // @[Switch.scala 41:38:@27350.4]
  wire  _T_66193; // @[Switch.scala 41:52:@27352.4]
  wire  output_26_17; // @[Switch.scala 41:38:@27353.4]
  wire  _T_66196; // @[Switch.scala 41:52:@27355.4]
  wire  output_26_18; // @[Switch.scala 41:38:@27356.4]
  wire  _T_66199; // @[Switch.scala 41:52:@27358.4]
  wire  output_26_19; // @[Switch.scala 41:38:@27359.4]
  wire  _T_66202; // @[Switch.scala 41:52:@27361.4]
  wire  output_26_20; // @[Switch.scala 41:38:@27362.4]
  wire  _T_66205; // @[Switch.scala 41:52:@27364.4]
  wire  output_26_21; // @[Switch.scala 41:38:@27365.4]
  wire  _T_66208; // @[Switch.scala 41:52:@27367.4]
  wire  output_26_22; // @[Switch.scala 41:38:@27368.4]
  wire  _T_66211; // @[Switch.scala 41:52:@27370.4]
  wire  output_26_23; // @[Switch.scala 41:38:@27371.4]
  wire  _T_66214; // @[Switch.scala 41:52:@27373.4]
  wire  output_26_24; // @[Switch.scala 41:38:@27374.4]
  wire  _T_66217; // @[Switch.scala 41:52:@27376.4]
  wire  output_26_25; // @[Switch.scala 41:38:@27377.4]
  wire  _T_66220; // @[Switch.scala 41:52:@27379.4]
  wire  output_26_26; // @[Switch.scala 41:38:@27380.4]
  wire  _T_66223; // @[Switch.scala 41:52:@27382.4]
  wire  output_26_27; // @[Switch.scala 41:38:@27383.4]
  wire  _T_66226; // @[Switch.scala 41:52:@27385.4]
  wire  output_26_28; // @[Switch.scala 41:38:@27386.4]
  wire  _T_66229; // @[Switch.scala 41:52:@27388.4]
  wire  output_26_29; // @[Switch.scala 41:38:@27389.4]
  wire  _T_66232; // @[Switch.scala 41:52:@27391.4]
  wire  output_26_30; // @[Switch.scala 41:38:@27392.4]
  wire  _T_66235; // @[Switch.scala 41:52:@27394.4]
  wire  output_26_31; // @[Switch.scala 41:38:@27395.4]
  wire  _T_66238; // @[Switch.scala 41:52:@27397.4]
  wire  output_26_32; // @[Switch.scala 41:38:@27398.4]
  wire  _T_66241; // @[Switch.scala 41:52:@27400.4]
  wire  output_26_33; // @[Switch.scala 41:38:@27401.4]
  wire  _T_66244; // @[Switch.scala 41:52:@27403.4]
  wire  output_26_34; // @[Switch.scala 41:38:@27404.4]
  wire  _T_66247; // @[Switch.scala 41:52:@27406.4]
  wire  output_26_35; // @[Switch.scala 41:38:@27407.4]
  wire  _T_66250; // @[Switch.scala 41:52:@27409.4]
  wire  output_26_36; // @[Switch.scala 41:38:@27410.4]
  wire  _T_66253; // @[Switch.scala 41:52:@27412.4]
  wire  output_26_37; // @[Switch.scala 41:38:@27413.4]
  wire  _T_66256; // @[Switch.scala 41:52:@27415.4]
  wire  output_26_38; // @[Switch.scala 41:38:@27416.4]
  wire  _T_66259; // @[Switch.scala 41:52:@27418.4]
  wire  output_26_39; // @[Switch.scala 41:38:@27419.4]
  wire  _T_66262; // @[Switch.scala 41:52:@27421.4]
  wire  output_26_40; // @[Switch.scala 41:38:@27422.4]
  wire  _T_66265; // @[Switch.scala 41:52:@27424.4]
  wire  output_26_41; // @[Switch.scala 41:38:@27425.4]
  wire  _T_66268; // @[Switch.scala 41:52:@27427.4]
  wire  output_26_42; // @[Switch.scala 41:38:@27428.4]
  wire  _T_66271; // @[Switch.scala 41:52:@27430.4]
  wire  output_26_43; // @[Switch.scala 41:38:@27431.4]
  wire  _T_66274; // @[Switch.scala 41:52:@27433.4]
  wire  output_26_44; // @[Switch.scala 41:38:@27434.4]
  wire  _T_66277; // @[Switch.scala 41:52:@27436.4]
  wire  output_26_45; // @[Switch.scala 41:38:@27437.4]
  wire  _T_66280; // @[Switch.scala 41:52:@27439.4]
  wire  output_26_46; // @[Switch.scala 41:38:@27440.4]
  wire  _T_66283; // @[Switch.scala 41:52:@27442.4]
  wire  output_26_47; // @[Switch.scala 41:38:@27443.4]
  wire  _T_66286; // @[Switch.scala 41:52:@27445.4]
  wire  output_26_48; // @[Switch.scala 41:38:@27446.4]
  wire  _T_66289; // @[Switch.scala 41:52:@27448.4]
  wire  output_26_49; // @[Switch.scala 41:38:@27449.4]
  wire  _T_66292; // @[Switch.scala 41:52:@27451.4]
  wire  output_26_50; // @[Switch.scala 41:38:@27452.4]
  wire  _T_66295; // @[Switch.scala 41:52:@27454.4]
  wire  output_26_51; // @[Switch.scala 41:38:@27455.4]
  wire  _T_66298; // @[Switch.scala 41:52:@27457.4]
  wire  output_26_52; // @[Switch.scala 41:38:@27458.4]
  wire  _T_66301; // @[Switch.scala 41:52:@27460.4]
  wire  output_26_53; // @[Switch.scala 41:38:@27461.4]
  wire  _T_66304; // @[Switch.scala 41:52:@27463.4]
  wire  output_26_54; // @[Switch.scala 41:38:@27464.4]
  wire  _T_66307; // @[Switch.scala 41:52:@27466.4]
  wire  output_26_55; // @[Switch.scala 41:38:@27467.4]
  wire  _T_66310; // @[Switch.scala 41:52:@27469.4]
  wire  output_26_56; // @[Switch.scala 41:38:@27470.4]
  wire  _T_66313; // @[Switch.scala 41:52:@27472.4]
  wire  output_26_57; // @[Switch.scala 41:38:@27473.4]
  wire  _T_66316; // @[Switch.scala 41:52:@27475.4]
  wire  output_26_58; // @[Switch.scala 41:38:@27476.4]
  wire  _T_66319; // @[Switch.scala 41:52:@27478.4]
  wire  output_26_59; // @[Switch.scala 41:38:@27479.4]
  wire  _T_66322; // @[Switch.scala 41:52:@27481.4]
  wire  output_26_60; // @[Switch.scala 41:38:@27482.4]
  wire  _T_66325; // @[Switch.scala 41:52:@27484.4]
  wire  output_26_61; // @[Switch.scala 41:38:@27485.4]
  wire  _T_66328; // @[Switch.scala 41:52:@27487.4]
  wire  output_26_62; // @[Switch.scala 41:38:@27488.4]
  wire  _T_66331; // @[Switch.scala 41:52:@27490.4]
  wire  output_26_63; // @[Switch.scala 41:38:@27491.4]
  wire [7:0] _T_66339; // @[Switch.scala 43:31:@27499.4]
  wire [15:0] _T_66347; // @[Switch.scala 43:31:@27507.4]
  wire [7:0] _T_66354; // @[Switch.scala 43:31:@27514.4]
  wire [31:0] _T_66363; // @[Switch.scala 43:31:@27523.4]
  wire [7:0] _T_66370; // @[Switch.scala 43:31:@27530.4]
  wire [15:0] _T_66378; // @[Switch.scala 43:31:@27538.4]
  wire [7:0] _T_66385; // @[Switch.scala 43:31:@27545.4]
  wire [31:0] _T_66394; // @[Switch.scala 43:31:@27554.4]
  wire [63:0] _T_66395; // @[Switch.scala 43:31:@27555.4]
  wire  _T_66399; // @[Switch.scala 41:52:@27558.4]
  wire  output_27_0; // @[Switch.scala 41:38:@27559.4]
  wire  _T_66402; // @[Switch.scala 41:52:@27561.4]
  wire  output_27_1; // @[Switch.scala 41:38:@27562.4]
  wire  _T_66405; // @[Switch.scala 41:52:@27564.4]
  wire  output_27_2; // @[Switch.scala 41:38:@27565.4]
  wire  _T_66408; // @[Switch.scala 41:52:@27567.4]
  wire  output_27_3; // @[Switch.scala 41:38:@27568.4]
  wire  _T_66411; // @[Switch.scala 41:52:@27570.4]
  wire  output_27_4; // @[Switch.scala 41:38:@27571.4]
  wire  _T_66414; // @[Switch.scala 41:52:@27573.4]
  wire  output_27_5; // @[Switch.scala 41:38:@27574.4]
  wire  _T_66417; // @[Switch.scala 41:52:@27576.4]
  wire  output_27_6; // @[Switch.scala 41:38:@27577.4]
  wire  _T_66420; // @[Switch.scala 41:52:@27579.4]
  wire  output_27_7; // @[Switch.scala 41:38:@27580.4]
  wire  _T_66423; // @[Switch.scala 41:52:@27582.4]
  wire  output_27_8; // @[Switch.scala 41:38:@27583.4]
  wire  _T_66426; // @[Switch.scala 41:52:@27585.4]
  wire  output_27_9; // @[Switch.scala 41:38:@27586.4]
  wire  _T_66429; // @[Switch.scala 41:52:@27588.4]
  wire  output_27_10; // @[Switch.scala 41:38:@27589.4]
  wire  _T_66432; // @[Switch.scala 41:52:@27591.4]
  wire  output_27_11; // @[Switch.scala 41:38:@27592.4]
  wire  _T_66435; // @[Switch.scala 41:52:@27594.4]
  wire  output_27_12; // @[Switch.scala 41:38:@27595.4]
  wire  _T_66438; // @[Switch.scala 41:52:@27597.4]
  wire  output_27_13; // @[Switch.scala 41:38:@27598.4]
  wire  _T_66441; // @[Switch.scala 41:52:@27600.4]
  wire  output_27_14; // @[Switch.scala 41:38:@27601.4]
  wire  _T_66444; // @[Switch.scala 41:52:@27603.4]
  wire  output_27_15; // @[Switch.scala 41:38:@27604.4]
  wire  _T_66447; // @[Switch.scala 41:52:@27606.4]
  wire  output_27_16; // @[Switch.scala 41:38:@27607.4]
  wire  _T_66450; // @[Switch.scala 41:52:@27609.4]
  wire  output_27_17; // @[Switch.scala 41:38:@27610.4]
  wire  _T_66453; // @[Switch.scala 41:52:@27612.4]
  wire  output_27_18; // @[Switch.scala 41:38:@27613.4]
  wire  _T_66456; // @[Switch.scala 41:52:@27615.4]
  wire  output_27_19; // @[Switch.scala 41:38:@27616.4]
  wire  _T_66459; // @[Switch.scala 41:52:@27618.4]
  wire  output_27_20; // @[Switch.scala 41:38:@27619.4]
  wire  _T_66462; // @[Switch.scala 41:52:@27621.4]
  wire  output_27_21; // @[Switch.scala 41:38:@27622.4]
  wire  _T_66465; // @[Switch.scala 41:52:@27624.4]
  wire  output_27_22; // @[Switch.scala 41:38:@27625.4]
  wire  _T_66468; // @[Switch.scala 41:52:@27627.4]
  wire  output_27_23; // @[Switch.scala 41:38:@27628.4]
  wire  _T_66471; // @[Switch.scala 41:52:@27630.4]
  wire  output_27_24; // @[Switch.scala 41:38:@27631.4]
  wire  _T_66474; // @[Switch.scala 41:52:@27633.4]
  wire  output_27_25; // @[Switch.scala 41:38:@27634.4]
  wire  _T_66477; // @[Switch.scala 41:52:@27636.4]
  wire  output_27_26; // @[Switch.scala 41:38:@27637.4]
  wire  _T_66480; // @[Switch.scala 41:52:@27639.4]
  wire  output_27_27; // @[Switch.scala 41:38:@27640.4]
  wire  _T_66483; // @[Switch.scala 41:52:@27642.4]
  wire  output_27_28; // @[Switch.scala 41:38:@27643.4]
  wire  _T_66486; // @[Switch.scala 41:52:@27645.4]
  wire  output_27_29; // @[Switch.scala 41:38:@27646.4]
  wire  _T_66489; // @[Switch.scala 41:52:@27648.4]
  wire  output_27_30; // @[Switch.scala 41:38:@27649.4]
  wire  _T_66492; // @[Switch.scala 41:52:@27651.4]
  wire  output_27_31; // @[Switch.scala 41:38:@27652.4]
  wire  _T_66495; // @[Switch.scala 41:52:@27654.4]
  wire  output_27_32; // @[Switch.scala 41:38:@27655.4]
  wire  _T_66498; // @[Switch.scala 41:52:@27657.4]
  wire  output_27_33; // @[Switch.scala 41:38:@27658.4]
  wire  _T_66501; // @[Switch.scala 41:52:@27660.4]
  wire  output_27_34; // @[Switch.scala 41:38:@27661.4]
  wire  _T_66504; // @[Switch.scala 41:52:@27663.4]
  wire  output_27_35; // @[Switch.scala 41:38:@27664.4]
  wire  _T_66507; // @[Switch.scala 41:52:@27666.4]
  wire  output_27_36; // @[Switch.scala 41:38:@27667.4]
  wire  _T_66510; // @[Switch.scala 41:52:@27669.4]
  wire  output_27_37; // @[Switch.scala 41:38:@27670.4]
  wire  _T_66513; // @[Switch.scala 41:52:@27672.4]
  wire  output_27_38; // @[Switch.scala 41:38:@27673.4]
  wire  _T_66516; // @[Switch.scala 41:52:@27675.4]
  wire  output_27_39; // @[Switch.scala 41:38:@27676.4]
  wire  _T_66519; // @[Switch.scala 41:52:@27678.4]
  wire  output_27_40; // @[Switch.scala 41:38:@27679.4]
  wire  _T_66522; // @[Switch.scala 41:52:@27681.4]
  wire  output_27_41; // @[Switch.scala 41:38:@27682.4]
  wire  _T_66525; // @[Switch.scala 41:52:@27684.4]
  wire  output_27_42; // @[Switch.scala 41:38:@27685.4]
  wire  _T_66528; // @[Switch.scala 41:52:@27687.4]
  wire  output_27_43; // @[Switch.scala 41:38:@27688.4]
  wire  _T_66531; // @[Switch.scala 41:52:@27690.4]
  wire  output_27_44; // @[Switch.scala 41:38:@27691.4]
  wire  _T_66534; // @[Switch.scala 41:52:@27693.4]
  wire  output_27_45; // @[Switch.scala 41:38:@27694.4]
  wire  _T_66537; // @[Switch.scala 41:52:@27696.4]
  wire  output_27_46; // @[Switch.scala 41:38:@27697.4]
  wire  _T_66540; // @[Switch.scala 41:52:@27699.4]
  wire  output_27_47; // @[Switch.scala 41:38:@27700.4]
  wire  _T_66543; // @[Switch.scala 41:52:@27702.4]
  wire  output_27_48; // @[Switch.scala 41:38:@27703.4]
  wire  _T_66546; // @[Switch.scala 41:52:@27705.4]
  wire  output_27_49; // @[Switch.scala 41:38:@27706.4]
  wire  _T_66549; // @[Switch.scala 41:52:@27708.4]
  wire  output_27_50; // @[Switch.scala 41:38:@27709.4]
  wire  _T_66552; // @[Switch.scala 41:52:@27711.4]
  wire  output_27_51; // @[Switch.scala 41:38:@27712.4]
  wire  _T_66555; // @[Switch.scala 41:52:@27714.4]
  wire  output_27_52; // @[Switch.scala 41:38:@27715.4]
  wire  _T_66558; // @[Switch.scala 41:52:@27717.4]
  wire  output_27_53; // @[Switch.scala 41:38:@27718.4]
  wire  _T_66561; // @[Switch.scala 41:52:@27720.4]
  wire  output_27_54; // @[Switch.scala 41:38:@27721.4]
  wire  _T_66564; // @[Switch.scala 41:52:@27723.4]
  wire  output_27_55; // @[Switch.scala 41:38:@27724.4]
  wire  _T_66567; // @[Switch.scala 41:52:@27726.4]
  wire  output_27_56; // @[Switch.scala 41:38:@27727.4]
  wire  _T_66570; // @[Switch.scala 41:52:@27729.4]
  wire  output_27_57; // @[Switch.scala 41:38:@27730.4]
  wire  _T_66573; // @[Switch.scala 41:52:@27732.4]
  wire  output_27_58; // @[Switch.scala 41:38:@27733.4]
  wire  _T_66576; // @[Switch.scala 41:52:@27735.4]
  wire  output_27_59; // @[Switch.scala 41:38:@27736.4]
  wire  _T_66579; // @[Switch.scala 41:52:@27738.4]
  wire  output_27_60; // @[Switch.scala 41:38:@27739.4]
  wire  _T_66582; // @[Switch.scala 41:52:@27741.4]
  wire  output_27_61; // @[Switch.scala 41:38:@27742.4]
  wire  _T_66585; // @[Switch.scala 41:52:@27744.4]
  wire  output_27_62; // @[Switch.scala 41:38:@27745.4]
  wire  _T_66588; // @[Switch.scala 41:52:@27747.4]
  wire  output_27_63; // @[Switch.scala 41:38:@27748.4]
  wire [7:0] _T_66596; // @[Switch.scala 43:31:@27756.4]
  wire [15:0] _T_66604; // @[Switch.scala 43:31:@27764.4]
  wire [7:0] _T_66611; // @[Switch.scala 43:31:@27771.4]
  wire [31:0] _T_66620; // @[Switch.scala 43:31:@27780.4]
  wire [7:0] _T_66627; // @[Switch.scala 43:31:@27787.4]
  wire [15:0] _T_66635; // @[Switch.scala 43:31:@27795.4]
  wire [7:0] _T_66642; // @[Switch.scala 43:31:@27802.4]
  wire [31:0] _T_66651; // @[Switch.scala 43:31:@27811.4]
  wire [63:0] _T_66652; // @[Switch.scala 43:31:@27812.4]
  wire  _T_66656; // @[Switch.scala 41:52:@27815.4]
  wire  output_28_0; // @[Switch.scala 41:38:@27816.4]
  wire  _T_66659; // @[Switch.scala 41:52:@27818.4]
  wire  output_28_1; // @[Switch.scala 41:38:@27819.4]
  wire  _T_66662; // @[Switch.scala 41:52:@27821.4]
  wire  output_28_2; // @[Switch.scala 41:38:@27822.4]
  wire  _T_66665; // @[Switch.scala 41:52:@27824.4]
  wire  output_28_3; // @[Switch.scala 41:38:@27825.4]
  wire  _T_66668; // @[Switch.scala 41:52:@27827.4]
  wire  output_28_4; // @[Switch.scala 41:38:@27828.4]
  wire  _T_66671; // @[Switch.scala 41:52:@27830.4]
  wire  output_28_5; // @[Switch.scala 41:38:@27831.4]
  wire  _T_66674; // @[Switch.scala 41:52:@27833.4]
  wire  output_28_6; // @[Switch.scala 41:38:@27834.4]
  wire  _T_66677; // @[Switch.scala 41:52:@27836.4]
  wire  output_28_7; // @[Switch.scala 41:38:@27837.4]
  wire  _T_66680; // @[Switch.scala 41:52:@27839.4]
  wire  output_28_8; // @[Switch.scala 41:38:@27840.4]
  wire  _T_66683; // @[Switch.scala 41:52:@27842.4]
  wire  output_28_9; // @[Switch.scala 41:38:@27843.4]
  wire  _T_66686; // @[Switch.scala 41:52:@27845.4]
  wire  output_28_10; // @[Switch.scala 41:38:@27846.4]
  wire  _T_66689; // @[Switch.scala 41:52:@27848.4]
  wire  output_28_11; // @[Switch.scala 41:38:@27849.4]
  wire  _T_66692; // @[Switch.scala 41:52:@27851.4]
  wire  output_28_12; // @[Switch.scala 41:38:@27852.4]
  wire  _T_66695; // @[Switch.scala 41:52:@27854.4]
  wire  output_28_13; // @[Switch.scala 41:38:@27855.4]
  wire  _T_66698; // @[Switch.scala 41:52:@27857.4]
  wire  output_28_14; // @[Switch.scala 41:38:@27858.4]
  wire  _T_66701; // @[Switch.scala 41:52:@27860.4]
  wire  output_28_15; // @[Switch.scala 41:38:@27861.4]
  wire  _T_66704; // @[Switch.scala 41:52:@27863.4]
  wire  output_28_16; // @[Switch.scala 41:38:@27864.4]
  wire  _T_66707; // @[Switch.scala 41:52:@27866.4]
  wire  output_28_17; // @[Switch.scala 41:38:@27867.4]
  wire  _T_66710; // @[Switch.scala 41:52:@27869.4]
  wire  output_28_18; // @[Switch.scala 41:38:@27870.4]
  wire  _T_66713; // @[Switch.scala 41:52:@27872.4]
  wire  output_28_19; // @[Switch.scala 41:38:@27873.4]
  wire  _T_66716; // @[Switch.scala 41:52:@27875.4]
  wire  output_28_20; // @[Switch.scala 41:38:@27876.4]
  wire  _T_66719; // @[Switch.scala 41:52:@27878.4]
  wire  output_28_21; // @[Switch.scala 41:38:@27879.4]
  wire  _T_66722; // @[Switch.scala 41:52:@27881.4]
  wire  output_28_22; // @[Switch.scala 41:38:@27882.4]
  wire  _T_66725; // @[Switch.scala 41:52:@27884.4]
  wire  output_28_23; // @[Switch.scala 41:38:@27885.4]
  wire  _T_66728; // @[Switch.scala 41:52:@27887.4]
  wire  output_28_24; // @[Switch.scala 41:38:@27888.4]
  wire  _T_66731; // @[Switch.scala 41:52:@27890.4]
  wire  output_28_25; // @[Switch.scala 41:38:@27891.4]
  wire  _T_66734; // @[Switch.scala 41:52:@27893.4]
  wire  output_28_26; // @[Switch.scala 41:38:@27894.4]
  wire  _T_66737; // @[Switch.scala 41:52:@27896.4]
  wire  output_28_27; // @[Switch.scala 41:38:@27897.4]
  wire  _T_66740; // @[Switch.scala 41:52:@27899.4]
  wire  output_28_28; // @[Switch.scala 41:38:@27900.4]
  wire  _T_66743; // @[Switch.scala 41:52:@27902.4]
  wire  output_28_29; // @[Switch.scala 41:38:@27903.4]
  wire  _T_66746; // @[Switch.scala 41:52:@27905.4]
  wire  output_28_30; // @[Switch.scala 41:38:@27906.4]
  wire  _T_66749; // @[Switch.scala 41:52:@27908.4]
  wire  output_28_31; // @[Switch.scala 41:38:@27909.4]
  wire  _T_66752; // @[Switch.scala 41:52:@27911.4]
  wire  output_28_32; // @[Switch.scala 41:38:@27912.4]
  wire  _T_66755; // @[Switch.scala 41:52:@27914.4]
  wire  output_28_33; // @[Switch.scala 41:38:@27915.4]
  wire  _T_66758; // @[Switch.scala 41:52:@27917.4]
  wire  output_28_34; // @[Switch.scala 41:38:@27918.4]
  wire  _T_66761; // @[Switch.scala 41:52:@27920.4]
  wire  output_28_35; // @[Switch.scala 41:38:@27921.4]
  wire  _T_66764; // @[Switch.scala 41:52:@27923.4]
  wire  output_28_36; // @[Switch.scala 41:38:@27924.4]
  wire  _T_66767; // @[Switch.scala 41:52:@27926.4]
  wire  output_28_37; // @[Switch.scala 41:38:@27927.4]
  wire  _T_66770; // @[Switch.scala 41:52:@27929.4]
  wire  output_28_38; // @[Switch.scala 41:38:@27930.4]
  wire  _T_66773; // @[Switch.scala 41:52:@27932.4]
  wire  output_28_39; // @[Switch.scala 41:38:@27933.4]
  wire  _T_66776; // @[Switch.scala 41:52:@27935.4]
  wire  output_28_40; // @[Switch.scala 41:38:@27936.4]
  wire  _T_66779; // @[Switch.scala 41:52:@27938.4]
  wire  output_28_41; // @[Switch.scala 41:38:@27939.4]
  wire  _T_66782; // @[Switch.scala 41:52:@27941.4]
  wire  output_28_42; // @[Switch.scala 41:38:@27942.4]
  wire  _T_66785; // @[Switch.scala 41:52:@27944.4]
  wire  output_28_43; // @[Switch.scala 41:38:@27945.4]
  wire  _T_66788; // @[Switch.scala 41:52:@27947.4]
  wire  output_28_44; // @[Switch.scala 41:38:@27948.4]
  wire  _T_66791; // @[Switch.scala 41:52:@27950.4]
  wire  output_28_45; // @[Switch.scala 41:38:@27951.4]
  wire  _T_66794; // @[Switch.scala 41:52:@27953.4]
  wire  output_28_46; // @[Switch.scala 41:38:@27954.4]
  wire  _T_66797; // @[Switch.scala 41:52:@27956.4]
  wire  output_28_47; // @[Switch.scala 41:38:@27957.4]
  wire  _T_66800; // @[Switch.scala 41:52:@27959.4]
  wire  output_28_48; // @[Switch.scala 41:38:@27960.4]
  wire  _T_66803; // @[Switch.scala 41:52:@27962.4]
  wire  output_28_49; // @[Switch.scala 41:38:@27963.4]
  wire  _T_66806; // @[Switch.scala 41:52:@27965.4]
  wire  output_28_50; // @[Switch.scala 41:38:@27966.4]
  wire  _T_66809; // @[Switch.scala 41:52:@27968.4]
  wire  output_28_51; // @[Switch.scala 41:38:@27969.4]
  wire  _T_66812; // @[Switch.scala 41:52:@27971.4]
  wire  output_28_52; // @[Switch.scala 41:38:@27972.4]
  wire  _T_66815; // @[Switch.scala 41:52:@27974.4]
  wire  output_28_53; // @[Switch.scala 41:38:@27975.4]
  wire  _T_66818; // @[Switch.scala 41:52:@27977.4]
  wire  output_28_54; // @[Switch.scala 41:38:@27978.4]
  wire  _T_66821; // @[Switch.scala 41:52:@27980.4]
  wire  output_28_55; // @[Switch.scala 41:38:@27981.4]
  wire  _T_66824; // @[Switch.scala 41:52:@27983.4]
  wire  output_28_56; // @[Switch.scala 41:38:@27984.4]
  wire  _T_66827; // @[Switch.scala 41:52:@27986.4]
  wire  output_28_57; // @[Switch.scala 41:38:@27987.4]
  wire  _T_66830; // @[Switch.scala 41:52:@27989.4]
  wire  output_28_58; // @[Switch.scala 41:38:@27990.4]
  wire  _T_66833; // @[Switch.scala 41:52:@27992.4]
  wire  output_28_59; // @[Switch.scala 41:38:@27993.4]
  wire  _T_66836; // @[Switch.scala 41:52:@27995.4]
  wire  output_28_60; // @[Switch.scala 41:38:@27996.4]
  wire  _T_66839; // @[Switch.scala 41:52:@27998.4]
  wire  output_28_61; // @[Switch.scala 41:38:@27999.4]
  wire  _T_66842; // @[Switch.scala 41:52:@28001.4]
  wire  output_28_62; // @[Switch.scala 41:38:@28002.4]
  wire  _T_66845; // @[Switch.scala 41:52:@28004.4]
  wire  output_28_63; // @[Switch.scala 41:38:@28005.4]
  wire [7:0] _T_66853; // @[Switch.scala 43:31:@28013.4]
  wire [15:0] _T_66861; // @[Switch.scala 43:31:@28021.4]
  wire [7:0] _T_66868; // @[Switch.scala 43:31:@28028.4]
  wire [31:0] _T_66877; // @[Switch.scala 43:31:@28037.4]
  wire [7:0] _T_66884; // @[Switch.scala 43:31:@28044.4]
  wire [15:0] _T_66892; // @[Switch.scala 43:31:@28052.4]
  wire [7:0] _T_66899; // @[Switch.scala 43:31:@28059.4]
  wire [31:0] _T_66908; // @[Switch.scala 43:31:@28068.4]
  wire [63:0] _T_66909; // @[Switch.scala 43:31:@28069.4]
  wire  _T_66913; // @[Switch.scala 41:52:@28072.4]
  wire  output_29_0; // @[Switch.scala 41:38:@28073.4]
  wire  _T_66916; // @[Switch.scala 41:52:@28075.4]
  wire  output_29_1; // @[Switch.scala 41:38:@28076.4]
  wire  _T_66919; // @[Switch.scala 41:52:@28078.4]
  wire  output_29_2; // @[Switch.scala 41:38:@28079.4]
  wire  _T_66922; // @[Switch.scala 41:52:@28081.4]
  wire  output_29_3; // @[Switch.scala 41:38:@28082.4]
  wire  _T_66925; // @[Switch.scala 41:52:@28084.4]
  wire  output_29_4; // @[Switch.scala 41:38:@28085.4]
  wire  _T_66928; // @[Switch.scala 41:52:@28087.4]
  wire  output_29_5; // @[Switch.scala 41:38:@28088.4]
  wire  _T_66931; // @[Switch.scala 41:52:@28090.4]
  wire  output_29_6; // @[Switch.scala 41:38:@28091.4]
  wire  _T_66934; // @[Switch.scala 41:52:@28093.4]
  wire  output_29_7; // @[Switch.scala 41:38:@28094.4]
  wire  _T_66937; // @[Switch.scala 41:52:@28096.4]
  wire  output_29_8; // @[Switch.scala 41:38:@28097.4]
  wire  _T_66940; // @[Switch.scala 41:52:@28099.4]
  wire  output_29_9; // @[Switch.scala 41:38:@28100.4]
  wire  _T_66943; // @[Switch.scala 41:52:@28102.4]
  wire  output_29_10; // @[Switch.scala 41:38:@28103.4]
  wire  _T_66946; // @[Switch.scala 41:52:@28105.4]
  wire  output_29_11; // @[Switch.scala 41:38:@28106.4]
  wire  _T_66949; // @[Switch.scala 41:52:@28108.4]
  wire  output_29_12; // @[Switch.scala 41:38:@28109.4]
  wire  _T_66952; // @[Switch.scala 41:52:@28111.4]
  wire  output_29_13; // @[Switch.scala 41:38:@28112.4]
  wire  _T_66955; // @[Switch.scala 41:52:@28114.4]
  wire  output_29_14; // @[Switch.scala 41:38:@28115.4]
  wire  _T_66958; // @[Switch.scala 41:52:@28117.4]
  wire  output_29_15; // @[Switch.scala 41:38:@28118.4]
  wire  _T_66961; // @[Switch.scala 41:52:@28120.4]
  wire  output_29_16; // @[Switch.scala 41:38:@28121.4]
  wire  _T_66964; // @[Switch.scala 41:52:@28123.4]
  wire  output_29_17; // @[Switch.scala 41:38:@28124.4]
  wire  _T_66967; // @[Switch.scala 41:52:@28126.4]
  wire  output_29_18; // @[Switch.scala 41:38:@28127.4]
  wire  _T_66970; // @[Switch.scala 41:52:@28129.4]
  wire  output_29_19; // @[Switch.scala 41:38:@28130.4]
  wire  _T_66973; // @[Switch.scala 41:52:@28132.4]
  wire  output_29_20; // @[Switch.scala 41:38:@28133.4]
  wire  _T_66976; // @[Switch.scala 41:52:@28135.4]
  wire  output_29_21; // @[Switch.scala 41:38:@28136.4]
  wire  _T_66979; // @[Switch.scala 41:52:@28138.4]
  wire  output_29_22; // @[Switch.scala 41:38:@28139.4]
  wire  _T_66982; // @[Switch.scala 41:52:@28141.4]
  wire  output_29_23; // @[Switch.scala 41:38:@28142.4]
  wire  _T_66985; // @[Switch.scala 41:52:@28144.4]
  wire  output_29_24; // @[Switch.scala 41:38:@28145.4]
  wire  _T_66988; // @[Switch.scala 41:52:@28147.4]
  wire  output_29_25; // @[Switch.scala 41:38:@28148.4]
  wire  _T_66991; // @[Switch.scala 41:52:@28150.4]
  wire  output_29_26; // @[Switch.scala 41:38:@28151.4]
  wire  _T_66994; // @[Switch.scala 41:52:@28153.4]
  wire  output_29_27; // @[Switch.scala 41:38:@28154.4]
  wire  _T_66997; // @[Switch.scala 41:52:@28156.4]
  wire  output_29_28; // @[Switch.scala 41:38:@28157.4]
  wire  _T_67000; // @[Switch.scala 41:52:@28159.4]
  wire  output_29_29; // @[Switch.scala 41:38:@28160.4]
  wire  _T_67003; // @[Switch.scala 41:52:@28162.4]
  wire  output_29_30; // @[Switch.scala 41:38:@28163.4]
  wire  _T_67006; // @[Switch.scala 41:52:@28165.4]
  wire  output_29_31; // @[Switch.scala 41:38:@28166.4]
  wire  _T_67009; // @[Switch.scala 41:52:@28168.4]
  wire  output_29_32; // @[Switch.scala 41:38:@28169.4]
  wire  _T_67012; // @[Switch.scala 41:52:@28171.4]
  wire  output_29_33; // @[Switch.scala 41:38:@28172.4]
  wire  _T_67015; // @[Switch.scala 41:52:@28174.4]
  wire  output_29_34; // @[Switch.scala 41:38:@28175.4]
  wire  _T_67018; // @[Switch.scala 41:52:@28177.4]
  wire  output_29_35; // @[Switch.scala 41:38:@28178.4]
  wire  _T_67021; // @[Switch.scala 41:52:@28180.4]
  wire  output_29_36; // @[Switch.scala 41:38:@28181.4]
  wire  _T_67024; // @[Switch.scala 41:52:@28183.4]
  wire  output_29_37; // @[Switch.scala 41:38:@28184.4]
  wire  _T_67027; // @[Switch.scala 41:52:@28186.4]
  wire  output_29_38; // @[Switch.scala 41:38:@28187.4]
  wire  _T_67030; // @[Switch.scala 41:52:@28189.4]
  wire  output_29_39; // @[Switch.scala 41:38:@28190.4]
  wire  _T_67033; // @[Switch.scala 41:52:@28192.4]
  wire  output_29_40; // @[Switch.scala 41:38:@28193.4]
  wire  _T_67036; // @[Switch.scala 41:52:@28195.4]
  wire  output_29_41; // @[Switch.scala 41:38:@28196.4]
  wire  _T_67039; // @[Switch.scala 41:52:@28198.4]
  wire  output_29_42; // @[Switch.scala 41:38:@28199.4]
  wire  _T_67042; // @[Switch.scala 41:52:@28201.4]
  wire  output_29_43; // @[Switch.scala 41:38:@28202.4]
  wire  _T_67045; // @[Switch.scala 41:52:@28204.4]
  wire  output_29_44; // @[Switch.scala 41:38:@28205.4]
  wire  _T_67048; // @[Switch.scala 41:52:@28207.4]
  wire  output_29_45; // @[Switch.scala 41:38:@28208.4]
  wire  _T_67051; // @[Switch.scala 41:52:@28210.4]
  wire  output_29_46; // @[Switch.scala 41:38:@28211.4]
  wire  _T_67054; // @[Switch.scala 41:52:@28213.4]
  wire  output_29_47; // @[Switch.scala 41:38:@28214.4]
  wire  _T_67057; // @[Switch.scala 41:52:@28216.4]
  wire  output_29_48; // @[Switch.scala 41:38:@28217.4]
  wire  _T_67060; // @[Switch.scala 41:52:@28219.4]
  wire  output_29_49; // @[Switch.scala 41:38:@28220.4]
  wire  _T_67063; // @[Switch.scala 41:52:@28222.4]
  wire  output_29_50; // @[Switch.scala 41:38:@28223.4]
  wire  _T_67066; // @[Switch.scala 41:52:@28225.4]
  wire  output_29_51; // @[Switch.scala 41:38:@28226.4]
  wire  _T_67069; // @[Switch.scala 41:52:@28228.4]
  wire  output_29_52; // @[Switch.scala 41:38:@28229.4]
  wire  _T_67072; // @[Switch.scala 41:52:@28231.4]
  wire  output_29_53; // @[Switch.scala 41:38:@28232.4]
  wire  _T_67075; // @[Switch.scala 41:52:@28234.4]
  wire  output_29_54; // @[Switch.scala 41:38:@28235.4]
  wire  _T_67078; // @[Switch.scala 41:52:@28237.4]
  wire  output_29_55; // @[Switch.scala 41:38:@28238.4]
  wire  _T_67081; // @[Switch.scala 41:52:@28240.4]
  wire  output_29_56; // @[Switch.scala 41:38:@28241.4]
  wire  _T_67084; // @[Switch.scala 41:52:@28243.4]
  wire  output_29_57; // @[Switch.scala 41:38:@28244.4]
  wire  _T_67087; // @[Switch.scala 41:52:@28246.4]
  wire  output_29_58; // @[Switch.scala 41:38:@28247.4]
  wire  _T_67090; // @[Switch.scala 41:52:@28249.4]
  wire  output_29_59; // @[Switch.scala 41:38:@28250.4]
  wire  _T_67093; // @[Switch.scala 41:52:@28252.4]
  wire  output_29_60; // @[Switch.scala 41:38:@28253.4]
  wire  _T_67096; // @[Switch.scala 41:52:@28255.4]
  wire  output_29_61; // @[Switch.scala 41:38:@28256.4]
  wire  _T_67099; // @[Switch.scala 41:52:@28258.4]
  wire  output_29_62; // @[Switch.scala 41:38:@28259.4]
  wire  _T_67102; // @[Switch.scala 41:52:@28261.4]
  wire  output_29_63; // @[Switch.scala 41:38:@28262.4]
  wire [7:0] _T_67110; // @[Switch.scala 43:31:@28270.4]
  wire [15:0] _T_67118; // @[Switch.scala 43:31:@28278.4]
  wire [7:0] _T_67125; // @[Switch.scala 43:31:@28285.4]
  wire [31:0] _T_67134; // @[Switch.scala 43:31:@28294.4]
  wire [7:0] _T_67141; // @[Switch.scala 43:31:@28301.4]
  wire [15:0] _T_67149; // @[Switch.scala 43:31:@28309.4]
  wire [7:0] _T_67156; // @[Switch.scala 43:31:@28316.4]
  wire [31:0] _T_67165; // @[Switch.scala 43:31:@28325.4]
  wire [63:0] _T_67166; // @[Switch.scala 43:31:@28326.4]
  wire  _T_67170; // @[Switch.scala 41:52:@28329.4]
  wire  output_30_0; // @[Switch.scala 41:38:@28330.4]
  wire  _T_67173; // @[Switch.scala 41:52:@28332.4]
  wire  output_30_1; // @[Switch.scala 41:38:@28333.4]
  wire  _T_67176; // @[Switch.scala 41:52:@28335.4]
  wire  output_30_2; // @[Switch.scala 41:38:@28336.4]
  wire  _T_67179; // @[Switch.scala 41:52:@28338.4]
  wire  output_30_3; // @[Switch.scala 41:38:@28339.4]
  wire  _T_67182; // @[Switch.scala 41:52:@28341.4]
  wire  output_30_4; // @[Switch.scala 41:38:@28342.4]
  wire  _T_67185; // @[Switch.scala 41:52:@28344.4]
  wire  output_30_5; // @[Switch.scala 41:38:@28345.4]
  wire  _T_67188; // @[Switch.scala 41:52:@28347.4]
  wire  output_30_6; // @[Switch.scala 41:38:@28348.4]
  wire  _T_67191; // @[Switch.scala 41:52:@28350.4]
  wire  output_30_7; // @[Switch.scala 41:38:@28351.4]
  wire  _T_67194; // @[Switch.scala 41:52:@28353.4]
  wire  output_30_8; // @[Switch.scala 41:38:@28354.4]
  wire  _T_67197; // @[Switch.scala 41:52:@28356.4]
  wire  output_30_9; // @[Switch.scala 41:38:@28357.4]
  wire  _T_67200; // @[Switch.scala 41:52:@28359.4]
  wire  output_30_10; // @[Switch.scala 41:38:@28360.4]
  wire  _T_67203; // @[Switch.scala 41:52:@28362.4]
  wire  output_30_11; // @[Switch.scala 41:38:@28363.4]
  wire  _T_67206; // @[Switch.scala 41:52:@28365.4]
  wire  output_30_12; // @[Switch.scala 41:38:@28366.4]
  wire  _T_67209; // @[Switch.scala 41:52:@28368.4]
  wire  output_30_13; // @[Switch.scala 41:38:@28369.4]
  wire  _T_67212; // @[Switch.scala 41:52:@28371.4]
  wire  output_30_14; // @[Switch.scala 41:38:@28372.4]
  wire  _T_67215; // @[Switch.scala 41:52:@28374.4]
  wire  output_30_15; // @[Switch.scala 41:38:@28375.4]
  wire  _T_67218; // @[Switch.scala 41:52:@28377.4]
  wire  output_30_16; // @[Switch.scala 41:38:@28378.4]
  wire  _T_67221; // @[Switch.scala 41:52:@28380.4]
  wire  output_30_17; // @[Switch.scala 41:38:@28381.4]
  wire  _T_67224; // @[Switch.scala 41:52:@28383.4]
  wire  output_30_18; // @[Switch.scala 41:38:@28384.4]
  wire  _T_67227; // @[Switch.scala 41:52:@28386.4]
  wire  output_30_19; // @[Switch.scala 41:38:@28387.4]
  wire  _T_67230; // @[Switch.scala 41:52:@28389.4]
  wire  output_30_20; // @[Switch.scala 41:38:@28390.4]
  wire  _T_67233; // @[Switch.scala 41:52:@28392.4]
  wire  output_30_21; // @[Switch.scala 41:38:@28393.4]
  wire  _T_67236; // @[Switch.scala 41:52:@28395.4]
  wire  output_30_22; // @[Switch.scala 41:38:@28396.4]
  wire  _T_67239; // @[Switch.scala 41:52:@28398.4]
  wire  output_30_23; // @[Switch.scala 41:38:@28399.4]
  wire  _T_67242; // @[Switch.scala 41:52:@28401.4]
  wire  output_30_24; // @[Switch.scala 41:38:@28402.4]
  wire  _T_67245; // @[Switch.scala 41:52:@28404.4]
  wire  output_30_25; // @[Switch.scala 41:38:@28405.4]
  wire  _T_67248; // @[Switch.scala 41:52:@28407.4]
  wire  output_30_26; // @[Switch.scala 41:38:@28408.4]
  wire  _T_67251; // @[Switch.scala 41:52:@28410.4]
  wire  output_30_27; // @[Switch.scala 41:38:@28411.4]
  wire  _T_67254; // @[Switch.scala 41:52:@28413.4]
  wire  output_30_28; // @[Switch.scala 41:38:@28414.4]
  wire  _T_67257; // @[Switch.scala 41:52:@28416.4]
  wire  output_30_29; // @[Switch.scala 41:38:@28417.4]
  wire  _T_67260; // @[Switch.scala 41:52:@28419.4]
  wire  output_30_30; // @[Switch.scala 41:38:@28420.4]
  wire  _T_67263; // @[Switch.scala 41:52:@28422.4]
  wire  output_30_31; // @[Switch.scala 41:38:@28423.4]
  wire  _T_67266; // @[Switch.scala 41:52:@28425.4]
  wire  output_30_32; // @[Switch.scala 41:38:@28426.4]
  wire  _T_67269; // @[Switch.scala 41:52:@28428.4]
  wire  output_30_33; // @[Switch.scala 41:38:@28429.4]
  wire  _T_67272; // @[Switch.scala 41:52:@28431.4]
  wire  output_30_34; // @[Switch.scala 41:38:@28432.4]
  wire  _T_67275; // @[Switch.scala 41:52:@28434.4]
  wire  output_30_35; // @[Switch.scala 41:38:@28435.4]
  wire  _T_67278; // @[Switch.scala 41:52:@28437.4]
  wire  output_30_36; // @[Switch.scala 41:38:@28438.4]
  wire  _T_67281; // @[Switch.scala 41:52:@28440.4]
  wire  output_30_37; // @[Switch.scala 41:38:@28441.4]
  wire  _T_67284; // @[Switch.scala 41:52:@28443.4]
  wire  output_30_38; // @[Switch.scala 41:38:@28444.4]
  wire  _T_67287; // @[Switch.scala 41:52:@28446.4]
  wire  output_30_39; // @[Switch.scala 41:38:@28447.4]
  wire  _T_67290; // @[Switch.scala 41:52:@28449.4]
  wire  output_30_40; // @[Switch.scala 41:38:@28450.4]
  wire  _T_67293; // @[Switch.scala 41:52:@28452.4]
  wire  output_30_41; // @[Switch.scala 41:38:@28453.4]
  wire  _T_67296; // @[Switch.scala 41:52:@28455.4]
  wire  output_30_42; // @[Switch.scala 41:38:@28456.4]
  wire  _T_67299; // @[Switch.scala 41:52:@28458.4]
  wire  output_30_43; // @[Switch.scala 41:38:@28459.4]
  wire  _T_67302; // @[Switch.scala 41:52:@28461.4]
  wire  output_30_44; // @[Switch.scala 41:38:@28462.4]
  wire  _T_67305; // @[Switch.scala 41:52:@28464.4]
  wire  output_30_45; // @[Switch.scala 41:38:@28465.4]
  wire  _T_67308; // @[Switch.scala 41:52:@28467.4]
  wire  output_30_46; // @[Switch.scala 41:38:@28468.4]
  wire  _T_67311; // @[Switch.scala 41:52:@28470.4]
  wire  output_30_47; // @[Switch.scala 41:38:@28471.4]
  wire  _T_67314; // @[Switch.scala 41:52:@28473.4]
  wire  output_30_48; // @[Switch.scala 41:38:@28474.4]
  wire  _T_67317; // @[Switch.scala 41:52:@28476.4]
  wire  output_30_49; // @[Switch.scala 41:38:@28477.4]
  wire  _T_67320; // @[Switch.scala 41:52:@28479.4]
  wire  output_30_50; // @[Switch.scala 41:38:@28480.4]
  wire  _T_67323; // @[Switch.scala 41:52:@28482.4]
  wire  output_30_51; // @[Switch.scala 41:38:@28483.4]
  wire  _T_67326; // @[Switch.scala 41:52:@28485.4]
  wire  output_30_52; // @[Switch.scala 41:38:@28486.4]
  wire  _T_67329; // @[Switch.scala 41:52:@28488.4]
  wire  output_30_53; // @[Switch.scala 41:38:@28489.4]
  wire  _T_67332; // @[Switch.scala 41:52:@28491.4]
  wire  output_30_54; // @[Switch.scala 41:38:@28492.4]
  wire  _T_67335; // @[Switch.scala 41:52:@28494.4]
  wire  output_30_55; // @[Switch.scala 41:38:@28495.4]
  wire  _T_67338; // @[Switch.scala 41:52:@28497.4]
  wire  output_30_56; // @[Switch.scala 41:38:@28498.4]
  wire  _T_67341; // @[Switch.scala 41:52:@28500.4]
  wire  output_30_57; // @[Switch.scala 41:38:@28501.4]
  wire  _T_67344; // @[Switch.scala 41:52:@28503.4]
  wire  output_30_58; // @[Switch.scala 41:38:@28504.4]
  wire  _T_67347; // @[Switch.scala 41:52:@28506.4]
  wire  output_30_59; // @[Switch.scala 41:38:@28507.4]
  wire  _T_67350; // @[Switch.scala 41:52:@28509.4]
  wire  output_30_60; // @[Switch.scala 41:38:@28510.4]
  wire  _T_67353; // @[Switch.scala 41:52:@28512.4]
  wire  output_30_61; // @[Switch.scala 41:38:@28513.4]
  wire  _T_67356; // @[Switch.scala 41:52:@28515.4]
  wire  output_30_62; // @[Switch.scala 41:38:@28516.4]
  wire  _T_67359; // @[Switch.scala 41:52:@28518.4]
  wire  output_30_63; // @[Switch.scala 41:38:@28519.4]
  wire [7:0] _T_67367; // @[Switch.scala 43:31:@28527.4]
  wire [15:0] _T_67375; // @[Switch.scala 43:31:@28535.4]
  wire [7:0] _T_67382; // @[Switch.scala 43:31:@28542.4]
  wire [31:0] _T_67391; // @[Switch.scala 43:31:@28551.4]
  wire [7:0] _T_67398; // @[Switch.scala 43:31:@28558.4]
  wire [15:0] _T_67406; // @[Switch.scala 43:31:@28566.4]
  wire [7:0] _T_67413; // @[Switch.scala 43:31:@28573.4]
  wire [31:0] _T_67422; // @[Switch.scala 43:31:@28582.4]
  wire [63:0] _T_67423; // @[Switch.scala 43:31:@28583.4]
  wire  _T_67427; // @[Switch.scala 41:52:@28586.4]
  wire  output_31_0; // @[Switch.scala 41:38:@28587.4]
  wire  _T_67430; // @[Switch.scala 41:52:@28589.4]
  wire  output_31_1; // @[Switch.scala 41:38:@28590.4]
  wire  _T_67433; // @[Switch.scala 41:52:@28592.4]
  wire  output_31_2; // @[Switch.scala 41:38:@28593.4]
  wire  _T_67436; // @[Switch.scala 41:52:@28595.4]
  wire  output_31_3; // @[Switch.scala 41:38:@28596.4]
  wire  _T_67439; // @[Switch.scala 41:52:@28598.4]
  wire  output_31_4; // @[Switch.scala 41:38:@28599.4]
  wire  _T_67442; // @[Switch.scala 41:52:@28601.4]
  wire  output_31_5; // @[Switch.scala 41:38:@28602.4]
  wire  _T_67445; // @[Switch.scala 41:52:@28604.4]
  wire  output_31_6; // @[Switch.scala 41:38:@28605.4]
  wire  _T_67448; // @[Switch.scala 41:52:@28607.4]
  wire  output_31_7; // @[Switch.scala 41:38:@28608.4]
  wire  _T_67451; // @[Switch.scala 41:52:@28610.4]
  wire  output_31_8; // @[Switch.scala 41:38:@28611.4]
  wire  _T_67454; // @[Switch.scala 41:52:@28613.4]
  wire  output_31_9; // @[Switch.scala 41:38:@28614.4]
  wire  _T_67457; // @[Switch.scala 41:52:@28616.4]
  wire  output_31_10; // @[Switch.scala 41:38:@28617.4]
  wire  _T_67460; // @[Switch.scala 41:52:@28619.4]
  wire  output_31_11; // @[Switch.scala 41:38:@28620.4]
  wire  _T_67463; // @[Switch.scala 41:52:@28622.4]
  wire  output_31_12; // @[Switch.scala 41:38:@28623.4]
  wire  _T_67466; // @[Switch.scala 41:52:@28625.4]
  wire  output_31_13; // @[Switch.scala 41:38:@28626.4]
  wire  _T_67469; // @[Switch.scala 41:52:@28628.4]
  wire  output_31_14; // @[Switch.scala 41:38:@28629.4]
  wire  _T_67472; // @[Switch.scala 41:52:@28631.4]
  wire  output_31_15; // @[Switch.scala 41:38:@28632.4]
  wire  _T_67475; // @[Switch.scala 41:52:@28634.4]
  wire  output_31_16; // @[Switch.scala 41:38:@28635.4]
  wire  _T_67478; // @[Switch.scala 41:52:@28637.4]
  wire  output_31_17; // @[Switch.scala 41:38:@28638.4]
  wire  _T_67481; // @[Switch.scala 41:52:@28640.4]
  wire  output_31_18; // @[Switch.scala 41:38:@28641.4]
  wire  _T_67484; // @[Switch.scala 41:52:@28643.4]
  wire  output_31_19; // @[Switch.scala 41:38:@28644.4]
  wire  _T_67487; // @[Switch.scala 41:52:@28646.4]
  wire  output_31_20; // @[Switch.scala 41:38:@28647.4]
  wire  _T_67490; // @[Switch.scala 41:52:@28649.4]
  wire  output_31_21; // @[Switch.scala 41:38:@28650.4]
  wire  _T_67493; // @[Switch.scala 41:52:@28652.4]
  wire  output_31_22; // @[Switch.scala 41:38:@28653.4]
  wire  _T_67496; // @[Switch.scala 41:52:@28655.4]
  wire  output_31_23; // @[Switch.scala 41:38:@28656.4]
  wire  _T_67499; // @[Switch.scala 41:52:@28658.4]
  wire  output_31_24; // @[Switch.scala 41:38:@28659.4]
  wire  _T_67502; // @[Switch.scala 41:52:@28661.4]
  wire  output_31_25; // @[Switch.scala 41:38:@28662.4]
  wire  _T_67505; // @[Switch.scala 41:52:@28664.4]
  wire  output_31_26; // @[Switch.scala 41:38:@28665.4]
  wire  _T_67508; // @[Switch.scala 41:52:@28667.4]
  wire  output_31_27; // @[Switch.scala 41:38:@28668.4]
  wire  _T_67511; // @[Switch.scala 41:52:@28670.4]
  wire  output_31_28; // @[Switch.scala 41:38:@28671.4]
  wire  _T_67514; // @[Switch.scala 41:52:@28673.4]
  wire  output_31_29; // @[Switch.scala 41:38:@28674.4]
  wire  _T_67517; // @[Switch.scala 41:52:@28676.4]
  wire  output_31_30; // @[Switch.scala 41:38:@28677.4]
  wire  _T_67520; // @[Switch.scala 41:52:@28679.4]
  wire  output_31_31; // @[Switch.scala 41:38:@28680.4]
  wire  _T_67523; // @[Switch.scala 41:52:@28682.4]
  wire  output_31_32; // @[Switch.scala 41:38:@28683.4]
  wire  _T_67526; // @[Switch.scala 41:52:@28685.4]
  wire  output_31_33; // @[Switch.scala 41:38:@28686.4]
  wire  _T_67529; // @[Switch.scala 41:52:@28688.4]
  wire  output_31_34; // @[Switch.scala 41:38:@28689.4]
  wire  _T_67532; // @[Switch.scala 41:52:@28691.4]
  wire  output_31_35; // @[Switch.scala 41:38:@28692.4]
  wire  _T_67535; // @[Switch.scala 41:52:@28694.4]
  wire  output_31_36; // @[Switch.scala 41:38:@28695.4]
  wire  _T_67538; // @[Switch.scala 41:52:@28697.4]
  wire  output_31_37; // @[Switch.scala 41:38:@28698.4]
  wire  _T_67541; // @[Switch.scala 41:52:@28700.4]
  wire  output_31_38; // @[Switch.scala 41:38:@28701.4]
  wire  _T_67544; // @[Switch.scala 41:52:@28703.4]
  wire  output_31_39; // @[Switch.scala 41:38:@28704.4]
  wire  _T_67547; // @[Switch.scala 41:52:@28706.4]
  wire  output_31_40; // @[Switch.scala 41:38:@28707.4]
  wire  _T_67550; // @[Switch.scala 41:52:@28709.4]
  wire  output_31_41; // @[Switch.scala 41:38:@28710.4]
  wire  _T_67553; // @[Switch.scala 41:52:@28712.4]
  wire  output_31_42; // @[Switch.scala 41:38:@28713.4]
  wire  _T_67556; // @[Switch.scala 41:52:@28715.4]
  wire  output_31_43; // @[Switch.scala 41:38:@28716.4]
  wire  _T_67559; // @[Switch.scala 41:52:@28718.4]
  wire  output_31_44; // @[Switch.scala 41:38:@28719.4]
  wire  _T_67562; // @[Switch.scala 41:52:@28721.4]
  wire  output_31_45; // @[Switch.scala 41:38:@28722.4]
  wire  _T_67565; // @[Switch.scala 41:52:@28724.4]
  wire  output_31_46; // @[Switch.scala 41:38:@28725.4]
  wire  _T_67568; // @[Switch.scala 41:52:@28727.4]
  wire  output_31_47; // @[Switch.scala 41:38:@28728.4]
  wire  _T_67571; // @[Switch.scala 41:52:@28730.4]
  wire  output_31_48; // @[Switch.scala 41:38:@28731.4]
  wire  _T_67574; // @[Switch.scala 41:52:@28733.4]
  wire  output_31_49; // @[Switch.scala 41:38:@28734.4]
  wire  _T_67577; // @[Switch.scala 41:52:@28736.4]
  wire  output_31_50; // @[Switch.scala 41:38:@28737.4]
  wire  _T_67580; // @[Switch.scala 41:52:@28739.4]
  wire  output_31_51; // @[Switch.scala 41:38:@28740.4]
  wire  _T_67583; // @[Switch.scala 41:52:@28742.4]
  wire  output_31_52; // @[Switch.scala 41:38:@28743.4]
  wire  _T_67586; // @[Switch.scala 41:52:@28745.4]
  wire  output_31_53; // @[Switch.scala 41:38:@28746.4]
  wire  _T_67589; // @[Switch.scala 41:52:@28748.4]
  wire  output_31_54; // @[Switch.scala 41:38:@28749.4]
  wire  _T_67592; // @[Switch.scala 41:52:@28751.4]
  wire  output_31_55; // @[Switch.scala 41:38:@28752.4]
  wire  _T_67595; // @[Switch.scala 41:52:@28754.4]
  wire  output_31_56; // @[Switch.scala 41:38:@28755.4]
  wire  _T_67598; // @[Switch.scala 41:52:@28757.4]
  wire  output_31_57; // @[Switch.scala 41:38:@28758.4]
  wire  _T_67601; // @[Switch.scala 41:52:@28760.4]
  wire  output_31_58; // @[Switch.scala 41:38:@28761.4]
  wire  _T_67604; // @[Switch.scala 41:52:@28763.4]
  wire  output_31_59; // @[Switch.scala 41:38:@28764.4]
  wire  _T_67607; // @[Switch.scala 41:52:@28766.4]
  wire  output_31_60; // @[Switch.scala 41:38:@28767.4]
  wire  _T_67610; // @[Switch.scala 41:52:@28769.4]
  wire  output_31_61; // @[Switch.scala 41:38:@28770.4]
  wire  _T_67613; // @[Switch.scala 41:52:@28772.4]
  wire  output_31_62; // @[Switch.scala 41:38:@28773.4]
  wire  _T_67616; // @[Switch.scala 41:52:@28775.4]
  wire  output_31_63; // @[Switch.scala 41:38:@28776.4]
  wire [7:0] _T_67624; // @[Switch.scala 43:31:@28784.4]
  wire [15:0] _T_67632; // @[Switch.scala 43:31:@28792.4]
  wire [7:0] _T_67639; // @[Switch.scala 43:31:@28799.4]
  wire [31:0] _T_67648; // @[Switch.scala 43:31:@28808.4]
  wire [7:0] _T_67655; // @[Switch.scala 43:31:@28815.4]
  wire [15:0] _T_67663; // @[Switch.scala 43:31:@28823.4]
  wire [7:0] _T_67670; // @[Switch.scala 43:31:@28830.4]
  wire [31:0] _T_67679; // @[Switch.scala 43:31:@28839.4]
  wire [63:0] _T_67680; // @[Switch.scala 43:31:@28840.4]
  wire  _T_67684; // @[Switch.scala 41:52:@28843.4]
  wire  output_32_0; // @[Switch.scala 41:38:@28844.4]
  wire  _T_67687; // @[Switch.scala 41:52:@28846.4]
  wire  output_32_1; // @[Switch.scala 41:38:@28847.4]
  wire  _T_67690; // @[Switch.scala 41:52:@28849.4]
  wire  output_32_2; // @[Switch.scala 41:38:@28850.4]
  wire  _T_67693; // @[Switch.scala 41:52:@28852.4]
  wire  output_32_3; // @[Switch.scala 41:38:@28853.4]
  wire  _T_67696; // @[Switch.scala 41:52:@28855.4]
  wire  output_32_4; // @[Switch.scala 41:38:@28856.4]
  wire  _T_67699; // @[Switch.scala 41:52:@28858.4]
  wire  output_32_5; // @[Switch.scala 41:38:@28859.4]
  wire  _T_67702; // @[Switch.scala 41:52:@28861.4]
  wire  output_32_6; // @[Switch.scala 41:38:@28862.4]
  wire  _T_67705; // @[Switch.scala 41:52:@28864.4]
  wire  output_32_7; // @[Switch.scala 41:38:@28865.4]
  wire  _T_67708; // @[Switch.scala 41:52:@28867.4]
  wire  output_32_8; // @[Switch.scala 41:38:@28868.4]
  wire  _T_67711; // @[Switch.scala 41:52:@28870.4]
  wire  output_32_9; // @[Switch.scala 41:38:@28871.4]
  wire  _T_67714; // @[Switch.scala 41:52:@28873.4]
  wire  output_32_10; // @[Switch.scala 41:38:@28874.4]
  wire  _T_67717; // @[Switch.scala 41:52:@28876.4]
  wire  output_32_11; // @[Switch.scala 41:38:@28877.4]
  wire  _T_67720; // @[Switch.scala 41:52:@28879.4]
  wire  output_32_12; // @[Switch.scala 41:38:@28880.4]
  wire  _T_67723; // @[Switch.scala 41:52:@28882.4]
  wire  output_32_13; // @[Switch.scala 41:38:@28883.4]
  wire  _T_67726; // @[Switch.scala 41:52:@28885.4]
  wire  output_32_14; // @[Switch.scala 41:38:@28886.4]
  wire  _T_67729; // @[Switch.scala 41:52:@28888.4]
  wire  output_32_15; // @[Switch.scala 41:38:@28889.4]
  wire  _T_67732; // @[Switch.scala 41:52:@28891.4]
  wire  output_32_16; // @[Switch.scala 41:38:@28892.4]
  wire  _T_67735; // @[Switch.scala 41:52:@28894.4]
  wire  output_32_17; // @[Switch.scala 41:38:@28895.4]
  wire  _T_67738; // @[Switch.scala 41:52:@28897.4]
  wire  output_32_18; // @[Switch.scala 41:38:@28898.4]
  wire  _T_67741; // @[Switch.scala 41:52:@28900.4]
  wire  output_32_19; // @[Switch.scala 41:38:@28901.4]
  wire  _T_67744; // @[Switch.scala 41:52:@28903.4]
  wire  output_32_20; // @[Switch.scala 41:38:@28904.4]
  wire  _T_67747; // @[Switch.scala 41:52:@28906.4]
  wire  output_32_21; // @[Switch.scala 41:38:@28907.4]
  wire  _T_67750; // @[Switch.scala 41:52:@28909.4]
  wire  output_32_22; // @[Switch.scala 41:38:@28910.4]
  wire  _T_67753; // @[Switch.scala 41:52:@28912.4]
  wire  output_32_23; // @[Switch.scala 41:38:@28913.4]
  wire  _T_67756; // @[Switch.scala 41:52:@28915.4]
  wire  output_32_24; // @[Switch.scala 41:38:@28916.4]
  wire  _T_67759; // @[Switch.scala 41:52:@28918.4]
  wire  output_32_25; // @[Switch.scala 41:38:@28919.4]
  wire  _T_67762; // @[Switch.scala 41:52:@28921.4]
  wire  output_32_26; // @[Switch.scala 41:38:@28922.4]
  wire  _T_67765; // @[Switch.scala 41:52:@28924.4]
  wire  output_32_27; // @[Switch.scala 41:38:@28925.4]
  wire  _T_67768; // @[Switch.scala 41:52:@28927.4]
  wire  output_32_28; // @[Switch.scala 41:38:@28928.4]
  wire  _T_67771; // @[Switch.scala 41:52:@28930.4]
  wire  output_32_29; // @[Switch.scala 41:38:@28931.4]
  wire  _T_67774; // @[Switch.scala 41:52:@28933.4]
  wire  output_32_30; // @[Switch.scala 41:38:@28934.4]
  wire  _T_67777; // @[Switch.scala 41:52:@28936.4]
  wire  output_32_31; // @[Switch.scala 41:38:@28937.4]
  wire  _T_67780; // @[Switch.scala 41:52:@28939.4]
  wire  output_32_32; // @[Switch.scala 41:38:@28940.4]
  wire  _T_67783; // @[Switch.scala 41:52:@28942.4]
  wire  output_32_33; // @[Switch.scala 41:38:@28943.4]
  wire  _T_67786; // @[Switch.scala 41:52:@28945.4]
  wire  output_32_34; // @[Switch.scala 41:38:@28946.4]
  wire  _T_67789; // @[Switch.scala 41:52:@28948.4]
  wire  output_32_35; // @[Switch.scala 41:38:@28949.4]
  wire  _T_67792; // @[Switch.scala 41:52:@28951.4]
  wire  output_32_36; // @[Switch.scala 41:38:@28952.4]
  wire  _T_67795; // @[Switch.scala 41:52:@28954.4]
  wire  output_32_37; // @[Switch.scala 41:38:@28955.4]
  wire  _T_67798; // @[Switch.scala 41:52:@28957.4]
  wire  output_32_38; // @[Switch.scala 41:38:@28958.4]
  wire  _T_67801; // @[Switch.scala 41:52:@28960.4]
  wire  output_32_39; // @[Switch.scala 41:38:@28961.4]
  wire  _T_67804; // @[Switch.scala 41:52:@28963.4]
  wire  output_32_40; // @[Switch.scala 41:38:@28964.4]
  wire  _T_67807; // @[Switch.scala 41:52:@28966.4]
  wire  output_32_41; // @[Switch.scala 41:38:@28967.4]
  wire  _T_67810; // @[Switch.scala 41:52:@28969.4]
  wire  output_32_42; // @[Switch.scala 41:38:@28970.4]
  wire  _T_67813; // @[Switch.scala 41:52:@28972.4]
  wire  output_32_43; // @[Switch.scala 41:38:@28973.4]
  wire  _T_67816; // @[Switch.scala 41:52:@28975.4]
  wire  output_32_44; // @[Switch.scala 41:38:@28976.4]
  wire  _T_67819; // @[Switch.scala 41:52:@28978.4]
  wire  output_32_45; // @[Switch.scala 41:38:@28979.4]
  wire  _T_67822; // @[Switch.scala 41:52:@28981.4]
  wire  output_32_46; // @[Switch.scala 41:38:@28982.4]
  wire  _T_67825; // @[Switch.scala 41:52:@28984.4]
  wire  output_32_47; // @[Switch.scala 41:38:@28985.4]
  wire  _T_67828; // @[Switch.scala 41:52:@28987.4]
  wire  output_32_48; // @[Switch.scala 41:38:@28988.4]
  wire  _T_67831; // @[Switch.scala 41:52:@28990.4]
  wire  output_32_49; // @[Switch.scala 41:38:@28991.4]
  wire  _T_67834; // @[Switch.scala 41:52:@28993.4]
  wire  output_32_50; // @[Switch.scala 41:38:@28994.4]
  wire  _T_67837; // @[Switch.scala 41:52:@28996.4]
  wire  output_32_51; // @[Switch.scala 41:38:@28997.4]
  wire  _T_67840; // @[Switch.scala 41:52:@28999.4]
  wire  output_32_52; // @[Switch.scala 41:38:@29000.4]
  wire  _T_67843; // @[Switch.scala 41:52:@29002.4]
  wire  output_32_53; // @[Switch.scala 41:38:@29003.4]
  wire  _T_67846; // @[Switch.scala 41:52:@29005.4]
  wire  output_32_54; // @[Switch.scala 41:38:@29006.4]
  wire  _T_67849; // @[Switch.scala 41:52:@29008.4]
  wire  output_32_55; // @[Switch.scala 41:38:@29009.4]
  wire  _T_67852; // @[Switch.scala 41:52:@29011.4]
  wire  output_32_56; // @[Switch.scala 41:38:@29012.4]
  wire  _T_67855; // @[Switch.scala 41:52:@29014.4]
  wire  output_32_57; // @[Switch.scala 41:38:@29015.4]
  wire  _T_67858; // @[Switch.scala 41:52:@29017.4]
  wire  output_32_58; // @[Switch.scala 41:38:@29018.4]
  wire  _T_67861; // @[Switch.scala 41:52:@29020.4]
  wire  output_32_59; // @[Switch.scala 41:38:@29021.4]
  wire  _T_67864; // @[Switch.scala 41:52:@29023.4]
  wire  output_32_60; // @[Switch.scala 41:38:@29024.4]
  wire  _T_67867; // @[Switch.scala 41:52:@29026.4]
  wire  output_32_61; // @[Switch.scala 41:38:@29027.4]
  wire  _T_67870; // @[Switch.scala 41:52:@29029.4]
  wire  output_32_62; // @[Switch.scala 41:38:@29030.4]
  wire  _T_67873; // @[Switch.scala 41:52:@29032.4]
  wire  output_32_63; // @[Switch.scala 41:38:@29033.4]
  wire [7:0] _T_67881; // @[Switch.scala 43:31:@29041.4]
  wire [15:0] _T_67889; // @[Switch.scala 43:31:@29049.4]
  wire [7:0] _T_67896; // @[Switch.scala 43:31:@29056.4]
  wire [31:0] _T_67905; // @[Switch.scala 43:31:@29065.4]
  wire [7:0] _T_67912; // @[Switch.scala 43:31:@29072.4]
  wire [15:0] _T_67920; // @[Switch.scala 43:31:@29080.4]
  wire [7:0] _T_67927; // @[Switch.scala 43:31:@29087.4]
  wire [31:0] _T_67936; // @[Switch.scala 43:31:@29096.4]
  wire [63:0] _T_67937; // @[Switch.scala 43:31:@29097.4]
  wire  _T_67941; // @[Switch.scala 41:52:@29100.4]
  wire  output_33_0; // @[Switch.scala 41:38:@29101.4]
  wire  _T_67944; // @[Switch.scala 41:52:@29103.4]
  wire  output_33_1; // @[Switch.scala 41:38:@29104.4]
  wire  _T_67947; // @[Switch.scala 41:52:@29106.4]
  wire  output_33_2; // @[Switch.scala 41:38:@29107.4]
  wire  _T_67950; // @[Switch.scala 41:52:@29109.4]
  wire  output_33_3; // @[Switch.scala 41:38:@29110.4]
  wire  _T_67953; // @[Switch.scala 41:52:@29112.4]
  wire  output_33_4; // @[Switch.scala 41:38:@29113.4]
  wire  _T_67956; // @[Switch.scala 41:52:@29115.4]
  wire  output_33_5; // @[Switch.scala 41:38:@29116.4]
  wire  _T_67959; // @[Switch.scala 41:52:@29118.4]
  wire  output_33_6; // @[Switch.scala 41:38:@29119.4]
  wire  _T_67962; // @[Switch.scala 41:52:@29121.4]
  wire  output_33_7; // @[Switch.scala 41:38:@29122.4]
  wire  _T_67965; // @[Switch.scala 41:52:@29124.4]
  wire  output_33_8; // @[Switch.scala 41:38:@29125.4]
  wire  _T_67968; // @[Switch.scala 41:52:@29127.4]
  wire  output_33_9; // @[Switch.scala 41:38:@29128.4]
  wire  _T_67971; // @[Switch.scala 41:52:@29130.4]
  wire  output_33_10; // @[Switch.scala 41:38:@29131.4]
  wire  _T_67974; // @[Switch.scala 41:52:@29133.4]
  wire  output_33_11; // @[Switch.scala 41:38:@29134.4]
  wire  _T_67977; // @[Switch.scala 41:52:@29136.4]
  wire  output_33_12; // @[Switch.scala 41:38:@29137.4]
  wire  _T_67980; // @[Switch.scala 41:52:@29139.4]
  wire  output_33_13; // @[Switch.scala 41:38:@29140.4]
  wire  _T_67983; // @[Switch.scala 41:52:@29142.4]
  wire  output_33_14; // @[Switch.scala 41:38:@29143.4]
  wire  _T_67986; // @[Switch.scala 41:52:@29145.4]
  wire  output_33_15; // @[Switch.scala 41:38:@29146.4]
  wire  _T_67989; // @[Switch.scala 41:52:@29148.4]
  wire  output_33_16; // @[Switch.scala 41:38:@29149.4]
  wire  _T_67992; // @[Switch.scala 41:52:@29151.4]
  wire  output_33_17; // @[Switch.scala 41:38:@29152.4]
  wire  _T_67995; // @[Switch.scala 41:52:@29154.4]
  wire  output_33_18; // @[Switch.scala 41:38:@29155.4]
  wire  _T_67998; // @[Switch.scala 41:52:@29157.4]
  wire  output_33_19; // @[Switch.scala 41:38:@29158.4]
  wire  _T_68001; // @[Switch.scala 41:52:@29160.4]
  wire  output_33_20; // @[Switch.scala 41:38:@29161.4]
  wire  _T_68004; // @[Switch.scala 41:52:@29163.4]
  wire  output_33_21; // @[Switch.scala 41:38:@29164.4]
  wire  _T_68007; // @[Switch.scala 41:52:@29166.4]
  wire  output_33_22; // @[Switch.scala 41:38:@29167.4]
  wire  _T_68010; // @[Switch.scala 41:52:@29169.4]
  wire  output_33_23; // @[Switch.scala 41:38:@29170.4]
  wire  _T_68013; // @[Switch.scala 41:52:@29172.4]
  wire  output_33_24; // @[Switch.scala 41:38:@29173.4]
  wire  _T_68016; // @[Switch.scala 41:52:@29175.4]
  wire  output_33_25; // @[Switch.scala 41:38:@29176.4]
  wire  _T_68019; // @[Switch.scala 41:52:@29178.4]
  wire  output_33_26; // @[Switch.scala 41:38:@29179.4]
  wire  _T_68022; // @[Switch.scala 41:52:@29181.4]
  wire  output_33_27; // @[Switch.scala 41:38:@29182.4]
  wire  _T_68025; // @[Switch.scala 41:52:@29184.4]
  wire  output_33_28; // @[Switch.scala 41:38:@29185.4]
  wire  _T_68028; // @[Switch.scala 41:52:@29187.4]
  wire  output_33_29; // @[Switch.scala 41:38:@29188.4]
  wire  _T_68031; // @[Switch.scala 41:52:@29190.4]
  wire  output_33_30; // @[Switch.scala 41:38:@29191.4]
  wire  _T_68034; // @[Switch.scala 41:52:@29193.4]
  wire  output_33_31; // @[Switch.scala 41:38:@29194.4]
  wire  _T_68037; // @[Switch.scala 41:52:@29196.4]
  wire  output_33_32; // @[Switch.scala 41:38:@29197.4]
  wire  _T_68040; // @[Switch.scala 41:52:@29199.4]
  wire  output_33_33; // @[Switch.scala 41:38:@29200.4]
  wire  _T_68043; // @[Switch.scala 41:52:@29202.4]
  wire  output_33_34; // @[Switch.scala 41:38:@29203.4]
  wire  _T_68046; // @[Switch.scala 41:52:@29205.4]
  wire  output_33_35; // @[Switch.scala 41:38:@29206.4]
  wire  _T_68049; // @[Switch.scala 41:52:@29208.4]
  wire  output_33_36; // @[Switch.scala 41:38:@29209.4]
  wire  _T_68052; // @[Switch.scala 41:52:@29211.4]
  wire  output_33_37; // @[Switch.scala 41:38:@29212.4]
  wire  _T_68055; // @[Switch.scala 41:52:@29214.4]
  wire  output_33_38; // @[Switch.scala 41:38:@29215.4]
  wire  _T_68058; // @[Switch.scala 41:52:@29217.4]
  wire  output_33_39; // @[Switch.scala 41:38:@29218.4]
  wire  _T_68061; // @[Switch.scala 41:52:@29220.4]
  wire  output_33_40; // @[Switch.scala 41:38:@29221.4]
  wire  _T_68064; // @[Switch.scala 41:52:@29223.4]
  wire  output_33_41; // @[Switch.scala 41:38:@29224.4]
  wire  _T_68067; // @[Switch.scala 41:52:@29226.4]
  wire  output_33_42; // @[Switch.scala 41:38:@29227.4]
  wire  _T_68070; // @[Switch.scala 41:52:@29229.4]
  wire  output_33_43; // @[Switch.scala 41:38:@29230.4]
  wire  _T_68073; // @[Switch.scala 41:52:@29232.4]
  wire  output_33_44; // @[Switch.scala 41:38:@29233.4]
  wire  _T_68076; // @[Switch.scala 41:52:@29235.4]
  wire  output_33_45; // @[Switch.scala 41:38:@29236.4]
  wire  _T_68079; // @[Switch.scala 41:52:@29238.4]
  wire  output_33_46; // @[Switch.scala 41:38:@29239.4]
  wire  _T_68082; // @[Switch.scala 41:52:@29241.4]
  wire  output_33_47; // @[Switch.scala 41:38:@29242.4]
  wire  _T_68085; // @[Switch.scala 41:52:@29244.4]
  wire  output_33_48; // @[Switch.scala 41:38:@29245.4]
  wire  _T_68088; // @[Switch.scala 41:52:@29247.4]
  wire  output_33_49; // @[Switch.scala 41:38:@29248.4]
  wire  _T_68091; // @[Switch.scala 41:52:@29250.4]
  wire  output_33_50; // @[Switch.scala 41:38:@29251.4]
  wire  _T_68094; // @[Switch.scala 41:52:@29253.4]
  wire  output_33_51; // @[Switch.scala 41:38:@29254.4]
  wire  _T_68097; // @[Switch.scala 41:52:@29256.4]
  wire  output_33_52; // @[Switch.scala 41:38:@29257.4]
  wire  _T_68100; // @[Switch.scala 41:52:@29259.4]
  wire  output_33_53; // @[Switch.scala 41:38:@29260.4]
  wire  _T_68103; // @[Switch.scala 41:52:@29262.4]
  wire  output_33_54; // @[Switch.scala 41:38:@29263.4]
  wire  _T_68106; // @[Switch.scala 41:52:@29265.4]
  wire  output_33_55; // @[Switch.scala 41:38:@29266.4]
  wire  _T_68109; // @[Switch.scala 41:52:@29268.4]
  wire  output_33_56; // @[Switch.scala 41:38:@29269.4]
  wire  _T_68112; // @[Switch.scala 41:52:@29271.4]
  wire  output_33_57; // @[Switch.scala 41:38:@29272.4]
  wire  _T_68115; // @[Switch.scala 41:52:@29274.4]
  wire  output_33_58; // @[Switch.scala 41:38:@29275.4]
  wire  _T_68118; // @[Switch.scala 41:52:@29277.4]
  wire  output_33_59; // @[Switch.scala 41:38:@29278.4]
  wire  _T_68121; // @[Switch.scala 41:52:@29280.4]
  wire  output_33_60; // @[Switch.scala 41:38:@29281.4]
  wire  _T_68124; // @[Switch.scala 41:52:@29283.4]
  wire  output_33_61; // @[Switch.scala 41:38:@29284.4]
  wire  _T_68127; // @[Switch.scala 41:52:@29286.4]
  wire  output_33_62; // @[Switch.scala 41:38:@29287.4]
  wire  _T_68130; // @[Switch.scala 41:52:@29289.4]
  wire  output_33_63; // @[Switch.scala 41:38:@29290.4]
  wire [7:0] _T_68138; // @[Switch.scala 43:31:@29298.4]
  wire [15:0] _T_68146; // @[Switch.scala 43:31:@29306.4]
  wire [7:0] _T_68153; // @[Switch.scala 43:31:@29313.4]
  wire [31:0] _T_68162; // @[Switch.scala 43:31:@29322.4]
  wire [7:0] _T_68169; // @[Switch.scala 43:31:@29329.4]
  wire [15:0] _T_68177; // @[Switch.scala 43:31:@29337.4]
  wire [7:0] _T_68184; // @[Switch.scala 43:31:@29344.4]
  wire [31:0] _T_68193; // @[Switch.scala 43:31:@29353.4]
  wire [63:0] _T_68194; // @[Switch.scala 43:31:@29354.4]
  wire  _T_68198; // @[Switch.scala 41:52:@29357.4]
  wire  output_34_0; // @[Switch.scala 41:38:@29358.4]
  wire  _T_68201; // @[Switch.scala 41:52:@29360.4]
  wire  output_34_1; // @[Switch.scala 41:38:@29361.4]
  wire  _T_68204; // @[Switch.scala 41:52:@29363.4]
  wire  output_34_2; // @[Switch.scala 41:38:@29364.4]
  wire  _T_68207; // @[Switch.scala 41:52:@29366.4]
  wire  output_34_3; // @[Switch.scala 41:38:@29367.4]
  wire  _T_68210; // @[Switch.scala 41:52:@29369.4]
  wire  output_34_4; // @[Switch.scala 41:38:@29370.4]
  wire  _T_68213; // @[Switch.scala 41:52:@29372.4]
  wire  output_34_5; // @[Switch.scala 41:38:@29373.4]
  wire  _T_68216; // @[Switch.scala 41:52:@29375.4]
  wire  output_34_6; // @[Switch.scala 41:38:@29376.4]
  wire  _T_68219; // @[Switch.scala 41:52:@29378.4]
  wire  output_34_7; // @[Switch.scala 41:38:@29379.4]
  wire  _T_68222; // @[Switch.scala 41:52:@29381.4]
  wire  output_34_8; // @[Switch.scala 41:38:@29382.4]
  wire  _T_68225; // @[Switch.scala 41:52:@29384.4]
  wire  output_34_9; // @[Switch.scala 41:38:@29385.4]
  wire  _T_68228; // @[Switch.scala 41:52:@29387.4]
  wire  output_34_10; // @[Switch.scala 41:38:@29388.4]
  wire  _T_68231; // @[Switch.scala 41:52:@29390.4]
  wire  output_34_11; // @[Switch.scala 41:38:@29391.4]
  wire  _T_68234; // @[Switch.scala 41:52:@29393.4]
  wire  output_34_12; // @[Switch.scala 41:38:@29394.4]
  wire  _T_68237; // @[Switch.scala 41:52:@29396.4]
  wire  output_34_13; // @[Switch.scala 41:38:@29397.4]
  wire  _T_68240; // @[Switch.scala 41:52:@29399.4]
  wire  output_34_14; // @[Switch.scala 41:38:@29400.4]
  wire  _T_68243; // @[Switch.scala 41:52:@29402.4]
  wire  output_34_15; // @[Switch.scala 41:38:@29403.4]
  wire  _T_68246; // @[Switch.scala 41:52:@29405.4]
  wire  output_34_16; // @[Switch.scala 41:38:@29406.4]
  wire  _T_68249; // @[Switch.scala 41:52:@29408.4]
  wire  output_34_17; // @[Switch.scala 41:38:@29409.4]
  wire  _T_68252; // @[Switch.scala 41:52:@29411.4]
  wire  output_34_18; // @[Switch.scala 41:38:@29412.4]
  wire  _T_68255; // @[Switch.scala 41:52:@29414.4]
  wire  output_34_19; // @[Switch.scala 41:38:@29415.4]
  wire  _T_68258; // @[Switch.scala 41:52:@29417.4]
  wire  output_34_20; // @[Switch.scala 41:38:@29418.4]
  wire  _T_68261; // @[Switch.scala 41:52:@29420.4]
  wire  output_34_21; // @[Switch.scala 41:38:@29421.4]
  wire  _T_68264; // @[Switch.scala 41:52:@29423.4]
  wire  output_34_22; // @[Switch.scala 41:38:@29424.4]
  wire  _T_68267; // @[Switch.scala 41:52:@29426.4]
  wire  output_34_23; // @[Switch.scala 41:38:@29427.4]
  wire  _T_68270; // @[Switch.scala 41:52:@29429.4]
  wire  output_34_24; // @[Switch.scala 41:38:@29430.4]
  wire  _T_68273; // @[Switch.scala 41:52:@29432.4]
  wire  output_34_25; // @[Switch.scala 41:38:@29433.4]
  wire  _T_68276; // @[Switch.scala 41:52:@29435.4]
  wire  output_34_26; // @[Switch.scala 41:38:@29436.4]
  wire  _T_68279; // @[Switch.scala 41:52:@29438.4]
  wire  output_34_27; // @[Switch.scala 41:38:@29439.4]
  wire  _T_68282; // @[Switch.scala 41:52:@29441.4]
  wire  output_34_28; // @[Switch.scala 41:38:@29442.4]
  wire  _T_68285; // @[Switch.scala 41:52:@29444.4]
  wire  output_34_29; // @[Switch.scala 41:38:@29445.4]
  wire  _T_68288; // @[Switch.scala 41:52:@29447.4]
  wire  output_34_30; // @[Switch.scala 41:38:@29448.4]
  wire  _T_68291; // @[Switch.scala 41:52:@29450.4]
  wire  output_34_31; // @[Switch.scala 41:38:@29451.4]
  wire  _T_68294; // @[Switch.scala 41:52:@29453.4]
  wire  output_34_32; // @[Switch.scala 41:38:@29454.4]
  wire  _T_68297; // @[Switch.scala 41:52:@29456.4]
  wire  output_34_33; // @[Switch.scala 41:38:@29457.4]
  wire  _T_68300; // @[Switch.scala 41:52:@29459.4]
  wire  output_34_34; // @[Switch.scala 41:38:@29460.4]
  wire  _T_68303; // @[Switch.scala 41:52:@29462.4]
  wire  output_34_35; // @[Switch.scala 41:38:@29463.4]
  wire  _T_68306; // @[Switch.scala 41:52:@29465.4]
  wire  output_34_36; // @[Switch.scala 41:38:@29466.4]
  wire  _T_68309; // @[Switch.scala 41:52:@29468.4]
  wire  output_34_37; // @[Switch.scala 41:38:@29469.4]
  wire  _T_68312; // @[Switch.scala 41:52:@29471.4]
  wire  output_34_38; // @[Switch.scala 41:38:@29472.4]
  wire  _T_68315; // @[Switch.scala 41:52:@29474.4]
  wire  output_34_39; // @[Switch.scala 41:38:@29475.4]
  wire  _T_68318; // @[Switch.scala 41:52:@29477.4]
  wire  output_34_40; // @[Switch.scala 41:38:@29478.4]
  wire  _T_68321; // @[Switch.scala 41:52:@29480.4]
  wire  output_34_41; // @[Switch.scala 41:38:@29481.4]
  wire  _T_68324; // @[Switch.scala 41:52:@29483.4]
  wire  output_34_42; // @[Switch.scala 41:38:@29484.4]
  wire  _T_68327; // @[Switch.scala 41:52:@29486.4]
  wire  output_34_43; // @[Switch.scala 41:38:@29487.4]
  wire  _T_68330; // @[Switch.scala 41:52:@29489.4]
  wire  output_34_44; // @[Switch.scala 41:38:@29490.4]
  wire  _T_68333; // @[Switch.scala 41:52:@29492.4]
  wire  output_34_45; // @[Switch.scala 41:38:@29493.4]
  wire  _T_68336; // @[Switch.scala 41:52:@29495.4]
  wire  output_34_46; // @[Switch.scala 41:38:@29496.4]
  wire  _T_68339; // @[Switch.scala 41:52:@29498.4]
  wire  output_34_47; // @[Switch.scala 41:38:@29499.4]
  wire  _T_68342; // @[Switch.scala 41:52:@29501.4]
  wire  output_34_48; // @[Switch.scala 41:38:@29502.4]
  wire  _T_68345; // @[Switch.scala 41:52:@29504.4]
  wire  output_34_49; // @[Switch.scala 41:38:@29505.4]
  wire  _T_68348; // @[Switch.scala 41:52:@29507.4]
  wire  output_34_50; // @[Switch.scala 41:38:@29508.4]
  wire  _T_68351; // @[Switch.scala 41:52:@29510.4]
  wire  output_34_51; // @[Switch.scala 41:38:@29511.4]
  wire  _T_68354; // @[Switch.scala 41:52:@29513.4]
  wire  output_34_52; // @[Switch.scala 41:38:@29514.4]
  wire  _T_68357; // @[Switch.scala 41:52:@29516.4]
  wire  output_34_53; // @[Switch.scala 41:38:@29517.4]
  wire  _T_68360; // @[Switch.scala 41:52:@29519.4]
  wire  output_34_54; // @[Switch.scala 41:38:@29520.4]
  wire  _T_68363; // @[Switch.scala 41:52:@29522.4]
  wire  output_34_55; // @[Switch.scala 41:38:@29523.4]
  wire  _T_68366; // @[Switch.scala 41:52:@29525.4]
  wire  output_34_56; // @[Switch.scala 41:38:@29526.4]
  wire  _T_68369; // @[Switch.scala 41:52:@29528.4]
  wire  output_34_57; // @[Switch.scala 41:38:@29529.4]
  wire  _T_68372; // @[Switch.scala 41:52:@29531.4]
  wire  output_34_58; // @[Switch.scala 41:38:@29532.4]
  wire  _T_68375; // @[Switch.scala 41:52:@29534.4]
  wire  output_34_59; // @[Switch.scala 41:38:@29535.4]
  wire  _T_68378; // @[Switch.scala 41:52:@29537.4]
  wire  output_34_60; // @[Switch.scala 41:38:@29538.4]
  wire  _T_68381; // @[Switch.scala 41:52:@29540.4]
  wire  output_34_61; // @[Switch.scala 41:38:@29541.4]
  wire  _T_68384; // @[Switch.scala 41:52:@29543.4]
  wire  output_34_62; // @[Switch.scala 41:38:@29544.4]
  wire  _T_68387; // @[Switch.scala 41:52:@29546.4]
  wire  output_34_63; // @[Switch.scala 41:38:@29547.4]
  wire [7:0] _T_68395; // @[Switch.scala 43:31:@29555.4]
  wire [15:0] _T_68403; // @[Switch.scala 43:31:@29563.4]
  wire [7:0] _T_68410; // @[Switch.scala 43:31:@29570.4]
  wire [31:0] _T_68419; // @[Switch.scala 43:31:@29579.4]
  wire [7:0] _T_68426; // @[Switch.scala 43:31:@29586.4]
  wire [15:0] _T_68434; // @[Switch.scala 43:31:@29594.4]
  wire [7:0] _T_68441; // @[Switch.scala 43:31:@29601.4]
  wire [31:0] _T_68450; // @[Switch.scala 43:31:@29610.4]
  wire [63:0] _T_68451; // @[Switch.scala 43:31:@29611.4]
  wire  _T_68455; // @[Switch.scala 41:52:@29614.4]
  wire  output_35_0; // @[Switch.scala 41:38:@29615.4]
  wire  _T_68458; // @[Switch.scala 41:52:@29617.4]
  wire  output_35_1; // @[Switch.scala 41:38:@29618.4]
  wire  _T_68461; // @[Switch.scala 41:52:@29620.4]
  wire  output_35_2; // @[Switch.scala 41:38:@29621.4]
  wire  _T_68464; // @[Switch.scala 41:52:@29623.4]
  wire  output_35_3; // @[Switch.scala 41:38:@29624.4]
  wire  _T_68467; // @[Switch.scala 41:52:@29626.4]
  wire  output_35_4; // @[Switch.scala 41:38:@29627.4]
  wire  _T_68470; // @[Switch.scala 41:52:@29629.4]
  wire  output_35_5; // @[Switch.scala 41:38:@29630.4]
  wire  _T_68473; // @[Switch.scala 41:52:@29632.4]
  wire  output_35_6; // @[Switch.scala 41:38:@29633.4]
  wire  _T_68476; // @[Switch.scala 41:52:@29635.4]
  wire  output_35_7; // @[Switch.scala 41:38:@29636.4]
  wire  _T_68479; // @[Switch.scala 41:52:@29638.4]
  wire  output_35_8; // @[Switch.scala 41:38:@29639.4]
  wire  _T_68482; // @[Switch.scala 41:52:@29641.4]
  wire  output_35_9; // @[Switch.scala 41:38:@29642.4]
  wire  _T_68485; // @[Switch.scala 41:52:@29644.4]
  wire  output_35_10; // @[Switch.scala 41:38:@29645.4]
  wire  _T_68488; // @[Switch.scala 41:52:@29647.4]
  wire  output_35_11; // @[Switch.scala 41:38:@29648.4]
  wire  _T_68491; // @[Switch.scala 41:52:@29650.4]
  wire  output_35_12; // @[Switch.scala 41:38:@29651.4]
  wire  _T_68494; // @[Switch.scala 41:52:@29653.4]
  wire  output_35_13; // @[Switch.scala 41:38:@29654.4]
  wire  _T_68497; // @[Switch.scala 41:52:@29656.4]
  wire  output_35_14; // @[Switch.scala 41:38:@29657.4]
  wire  _T_68500; // @[Switch.scala 41:52:@29659.4]
  wire  output_35_15; // @[Switch.scala 41:38:@29660.4]
  wire  _T_68503; // @[Switch.scala 41:52:@29662.4]
  wire  output_35_16; // @[Switch.scala 41:38:@29663.4]
  wire  _T_68506; // @[Switch.scala 41:52:@29665.4]
  wire  output_35_17; // @[Switch.scala 41:38:@29666.4]
  wire  _T_68509; // @[Switch.scala 41:52:@29668.4]
  wire  output_35_18; // @[Switch.scala 41:38:@29669.4]
  wire  _T_68512; // @[Switch.scala 41:52:@29671.4]
  wire  output_35_19; // @[Switch.scala 41:38:@29672.4]
  wire  _T_68515; // @[Switch.scala 41:52:@29674.4]
  wire  output_35_20; // @[Switch.scala 41:38:@29675.4]
  wire  _T_68518; // @[Switch.scala 41:52:@29677.4]
  wire  output_35_21; // @[Switch.scala 41:38:@29678.4]
  wire  _T_68521; // @[Switch.scala 41:52:@29680.4]
  wire  output_35_22; // @[Switch.scala 41:38:@29681.4]
  wire  _T_68524; // @[Switch.scala 41:52:@29683.4]
  wire  output_35_23; // @[Switch.scala 41:38:@29684.4]
  wire  _T_68527; // @[Switch.scala 41:52:@29686.4]
  wire  output_35_24; // @[Switch.scala 41:38:@29687.4]
  wire  _T_68530; // @[Switch.scala 41:52:@29689.4]
  wire  output_35_25; // @[Switch.scala 41:38:@29690.4]
  wire  _T_68533; // @[Switch.scala 41:52:@29692.4]
  wire  output_35_26; // @[Switch.scala 41:38:@29693.4]
  wire  _T_68536; // @[Switch.scala 41:52:@29695.4]
  wire  output_35_27; // @[Switch.scala 41:38:@29696.4]
  wire  _T_68539; // @[Switch.scala 41:52:@29698.4]
  wire  output_35_28; // @[Switch.scala 41:38:@29699.4]
  wire  _T_68542; // @[Switch.scala 41:52:@29701.4]
  wire  output_35_29; // @[Switch.scala 41:38:@29702.4]
  wire  _T_68545; // @[Switch.scala 41:52:@29704.4]
  wire  output_35_30; // @[Switch.scala 41:38:@29705.4]
  wire  _T_68548; // @[Switch.scala 41:52:@29707.4]
  wire  output_35_31; // @[Switch.scala 41:38:@29708.4]
  wire  _T_68551; // @[Switch.scala 41:52:@29710.4]
  wire  output_35_32; // @[Switch.scala 41:38:@29711.4]
  wire  _T_68554; // @[Switch.scala 41:52:@29713.4]
  wire  output_35_33; // @[Switch.scala 41:38:@29714.4]
  wire  _T_68557; // @[Switch.scala 41:52:@29716.4]
  wire  output_35_34; // @[Switch.scala 41:38:@29717.4]
  wire  _T_68560; // @[Switch.scala 41:52:@29719.4]
  wire  output_35_35; // @[Switch.scala 41:38:@29720.4]
  wire  _T_68563; // @[Switch.scala 41:52:@29722.4]
  wire  output_35_36; // @[Switch.scala 41:38:@29723.4]
  wire  _T_68566; // @[Switch.scala 41:52:@29725.4]
  wire  output_35_37; // @[Switch.scala 41:38:@29726.4]
  wire  _T_68569; // @[Switch.scala 41:52:@29728.4]
  wire  output_35_38; // @[Switch.scala 41:38:@29729.4]
  wire  _T_68572; // @[Switch.scala 41:52:@29731.4]
  wire  output_35_39; // @[Switch.scala 41:38:@29732.4]
  wire  _T_68575; // @[Switch.scala 41:52:@29734.4]
  wire  output_35_40; // @[Switch.scala 41:38:@29735.4]
  wire  _T_68578; // @[Switch.scala 41:52:@29737.4]
  wire  output_35_41; // @[Switch.scala 41:38:@29738.4]
  wire  _T_68581; // @[Switch.scala 41:52:@29740.4]
  wire  output_35_42; // @[Switch.scala 41:38:@29741.4]
  wire  _T_68584; // @[Switch.scala 41:52:@29743.4]
  wire  output_35_43; // @[Switch.scala 41:38:@29744.4]
  wire  _T_68587; // @[Switch.scala 41:52:@29746.4]
  wire  output_35_44; // @[Switch.scala 41:38:@29747.4]
  wire  _T_68590; // @[Switch.scala 41:52:@29749.4]
  wire  output_35_45; // @[Switch.scala 41:38:@29750.4]
  wire  _T_68593; // @[Switch.scala 41:52:@29752.4]
  wire  output_35_46; // @[Switch.scala 41:38:@29753.4]
  wire  _T_68596; // @[Switch.scala 41:52:@29755.4]
  wire  output_35_47; // @[Switch.scala 41:38:@29756.4]
  wire  _T_68599; // @[Switch.scala 41:52:@29758.4]
  wire  output_35_48; // @[Switch.scala 41:38:@29759.4]
  wire  _T_68602; // @[Switch.scala 41:52:@29761.4]
  wire  output_35_49; // @[Switch.scala 41:38:@29762.4]
  wire  _T_68605; // @[Switch.scala 41:52:@29764.4]
  wire  output_35_50; // @[Switch.scala 41:38:@29765.4]
  wire  _T_68608; // @[Switch.scala 41:52:@29767.4]
  wire  output_35_51; // @[Switch.scala 41:38:@29768.4]
  wire  _T_68611; // @[Switch.scala 41:52:@29770.4]
  wire  output_35_52; // @[Switch.scala 41:38:@29771.4]
  wire  _T_68614; // @[Switch.scala 41:52:@29773.4]
  wire  output_35_53; // @[Switch.scala 41:38:@29774.4]
  wire  _T_68617; // @[Switch.scala 41:52:@29776.4]
  wire  output_35_54; // @[Switch.scala 41:38:@29777.4]
  wire  _T_68620; // @[Switch.scala 41:52:@29779.4]
  wire  output_35_55; // @[Switch.scala 41:38:@29780.4]
  wire  _T_68623; // @[Switch.scala 41:52:@29782.4]
  wire  output_35_56; // @[Switch.scala 41:38:@29783.4]
  wire  _T_68626; // @[Switch.scala 41:52:@29785.4]
  wire  output_35_57; // @[Switch.scala 41:38:@29786.4]
  wire  _T_68629; // @[Switch.scala 41:52:@29788.4]
  wire  output_35_58; // @[Switch.scala 41:38:@29789.4]
  wire  _T_68632; // @[Switch.scala 41:52:@29791.4]
  wire  output_35_59; // @[Switch.scala 41:38:@29792.4]
  wire  _T_68635; // @[Switch.scala 41:52:@29794.4]
  wire  output_35_60; // @[Switch.scala 41:38:@29795.4]
  wire  _T_68638; // @[Switch.scala 41:52:@29797.4]
  wire  output_35_61; // @[Switch.scala 41:38:@29798.4]
  wire  _T_68641; // @[Switch.scala 41:52:@29800.4]
  wire  output_35_62; // @[Switch.scala 41:38:@29801.4]
  wire  _T_68644; // @[Switch.scala 41:52:@29803.4]
  wire  output_35_63; // @[Switch.scala 41:38:@29804.4]
  wire [7:0] _T_68652; // @[Switch.scala 43:31:@29812.4]
  wire [15:0] _T_68660; // @[Switch.scala 43:31:@29820.4]
  wire [7:0] _T_68667; // @[Switch.scala 43:31:@29827.4]
  wire [31:0] _T_68676; // @[Switch.scala 43:31:@29836.4]
  wire [7:0] _T_68683; // @[Switch.scala 43:31:@29843.4]
  wire [15:0] _T_68691; // @[Switch.scala 43:31:@29851.4]
  wire [7:0] _T_68698; // @[Switch.scala 43:31:@29858.4]
  wire [31:0] _T_68707; // @[Switch.scala 43:31:@29867.4]
  wire [63:0] _T_68708; // @[Switch.scala 43:31:@29868.4]
  wire  _T_68712; // @[Switch.scala 41:52:@29871.4]
  wire  output_36_0; // @[Switch.scala 41:38:@29872.4]
  wire  _T_68715; // @[Switch.scala 41:52:@29874.4]
  wire  output_36_1; // @[Switch.scala 41:38:@29875.4]
  wire  _T_68718; // @[Switch.scala 41:52:@29877.4]
  wire  output_36_2; // @[Switch.scala 41:38:@29878.4]
  wire  _T_68721; // @[Switch.scala 41:52:@29880.4]
  wire  output_36_3; // @[Switch.scala 41:38:@29881.4]
  wire  _T_68724; // @[Switch.scala 41:52:@29883.4]
  wire  output_36_4; // @[Switch.scala 41:38:@29884.4]
  wire  _T_68727; // @[Switch.scala 41:52:@29886.4]
  wire  output_36_5; // @[Switch.scala 41:38:@29887.4]
  wire  _T_68730; // @[Switch.scala 41:52:@29889.4]
  wire  output_36_6; // @[Switch.scala 41:38:@29890.4]
  wire  _T_68733; // @[Switch.scala 41:52:@29892.4]
  wire  output_36_7; // @[Switch.scala 41:38:@29893.4]
  wire  _T_68736; // @[Switch.scala 41:52:@29895.4]
  wire  output_36_8; // @[Switch.scala 41:38:@29896.4]
  wire  _T_68739; // @[Switch.scala 41:52:@29898.4]
  wire  output_36_9; // @[Switch.scala 41:38:@29899.4]
  wire  _T_68742; // @[Switch.scala 41:52:@29901.4]
  wire  output_36_10; // @[Switch.scala 41:38:@29902.4]
  wire  _T_68745; // @[Switch.scala 41:52:@29904.4]
  wire  output_36_11; // @[Switch.scala 41:38:@29905.4]
  wire  _T_68748; // @[Switch.scala 41:52:@29907.4]
  wire  output_36_12; // @[Switch.scala 41:38:@29908.4]
  wire  _T_68751; // @[Switch.scala 41:52:@29910.4]
  wire  output_36_13; // @[Switch.scala 41:38:@29911.4]
  wire  _T_68754; // @[Switch.scala 41:52:@29913.4]
  wire  output_36_14; // @[Switch.scala 41:38:@29914.4]
  wire  _T_68757; // @[Switch.scala 41:52:@29916.4]
  wire  output_36_15; // @[Switch.scala 41:38:@29917.4]
  wire  _T_68760; // @[Switch.scala 41:52:@29919.4]
  wire  output_36_16; // @[Switch.scala 41:38:@29920.4]
  wire  _T_68763; // @[Switch.scala 41:52:@29922.4]
  wire  output_36_17; // @[Switch.scala 41:38:@29923.4]
  wire  _T_68766; // @[Switch.scala 41:52:@29925.4]
  wire  output_36_18; // @[Switch.scala 41:38:@29926.4]
  wire  _T_68769; // @[Switch.scala 41:52:@29928.4]
  wire  output_36_19; // @[Switch.scala 41:38:@29929.4]
  wire  _T_68772; // @[Switch.scala 41:52:@29931.4]
  wire  output_36_20; // @[Switch.scala 41:38:@29932.4]
  wire  _T_68775; // @[Switch.scala 41:52:@29934.4]
  wire  output_36_21; // @[Switch.scala 41:38:@29935.4]
  wire  _T_68778; // @[Switch.scala 41:52:@29937.4]
  wire  output_36_22; // @[Switch.scala 41:38:@29938.4]
  wire  _T_68781; // @[Switch.scala 41:52:@29940.4]
  wire  output_36_23; // @[Switch.scala 41:38:@29941.4]
  wire  _T_68784; // @[Switch.scala 41:52:@29943.4]
  wire  output_36_24; // @[Switch.scala 41:38:@29944.4]
  wire  _T_68787; // @[Switch.scala 41:52:@29946.4]
  wire  output_36_25; // @[Switch.scala 41:38:@29947.4]
  wire  _T_68790; // @[Switch.scala 41:52:@29949.4]
  wire  output_36_26; // @[Switch.scala 41:38:@29950.4]
  wire  _T_68793; // @[Switch.scala 41:52:@29952.4]
  wire  output_36_27; // @[Switch.scala 41:38:@29953.4]
  wire  _T_68796; // @[Switch.scala 41:52:@29955.4]
  wire  output_36_28; // @[Switch.scala 41:38:@29956.4]
  wire  _T_68799; // @[Switch.scala 41:52:@29958.4]
  wire  output_36_29; // @[Switch.scala 41:38:@29959.4]
  wire  _T_68802; // @[Switch.scala 41:52:@29961.4]
  wire  output_36_30; // @[Switch.scala 41:38:@29962.4]
  wire  _T_68805; // @[Switch.scala 41:52:@29964.4]
  wire  output_36_31; // @[Switch.scala 41:38:@29965.4]
  wire  _T_68808; // @[Switch.scala 41:52:@29967.4]
  wire  output_36_32; // @[Switch.scala 41:38:@29968.4]
  wire  _T_68811; // @[Switch.scala 41:52:@29970.4]
  wire  output_36_33; // @[Switch.scala 41:38:@29971.4]
  wire  _T_68814; // @[Switch.scala 41:52:@29973.4]
  wire  output_36_34; // @[Switch.scala 41:38:@29974.4]
  wire  _T_68817; // @[Switch.scala 41:52:@29976.4]
  wire  output_36_35; // @[Switch.scala 41:38:@29977.4]
  wire  _T_68820; // @[Switch.scala 41:52:@29979.4]
  wire  output_36_36; // @[Switch.scala 41:38:@29980.4]
  wire  _T_68823; // @[Switch.scala 41:52:@29982.4]
  wire  output_36_37; // @[Switch.scala 41:38:@29983.4]
  wire  _T_68826; // @[Switch.scala 41:52:@29985.4]
  wire  output_36_38; // @[Switch.scala 41:38:@29986.4]
  wire  _T_68829; // @[Switch.scala 41:52:@29988.4]
  wire  output_36_39; // @[Switch.scala 41:38:@29989.4]
  wire  _T_68832; // @[Switch.scala 41:52:@29991.4]
  wire  output_36_40; // @[Switch.scala 41:38:@29992.4]
  wire  _T_68835; // @[Switch.scala 41:52:@29994.4]
  wire  output_36_41; // @[Switch.scala 41:38:@29995.4]
  wire  _T_68838; // @[Switch.scala 41:52:@29997.4]
  wire  output_36_42; // @[Switch.scala 41:38:@29998.4]
  wire  _T_68841; // @[Switch.scala 41:52:@30000.4]
  wire  output_36_43; // @[Switch.scala 41:38:@30001.4]
  wire  _T_68844; // @[Switch.scala 41:52:@30003.4]
  wire  output_36_44; // @[Switch.scala 41:38:@30004.4]
  wire  _T_68847; // @[Switch.scala 41:52:@30006.4]
  wire  output_36_45; // @[Switch.scala 41:38:@30007.4]
  wire  _T_68850; // @[Switch.scala 41:52:@30009.4]
  wire  output_36_46; // @[Switch.scala 41:38:@30010.4]
  wire  _T_68853; // @[Switch.scala 41:52:@30012.4]
  wire  output_36_47; // @[Switch.scala 41:38:@30013.4]
  wire  _T_68856; // @[Switch.scala 41:52:@30015.4]
  wire  output_36_48; // @[Switch.scala 41:38:@30016.4]
  wire  _T_68859; // @[Switch.scala 41:52:@30018.4]
  wire  output_36_49; // @[Switch.scala 41:38:@30019.4]
  wire  _T_68862; // @[Switch.scala 41:52:@30021.4]
  wire  output_36_50; // @[Switch.scala 41:38:@30022.4]
  wire  _T_68865; // @[Switch.scala 41:52:@30024.4]
  wire  output_36_51; // @[Switch.scala 41:38:@30025.4]
  wire  _T_68868; // @[Switch.scala 41:52:@30027.4]
  wire  output_36_52; // @[Switch.scala 41:38:@30028.4]
  wire  _T_68871; // @[Switch.scala 41:52:@30030.4]
  wire  output_36_53; // @[Switch.scala 41:38:@30031.4]
  wire  _T_68874; // @[Switch.scala 41:52:@30033.4]
  wire  output_36_54; // @[Switch.scala 41:38:@30034.4]
  wire  _T_68877; // @[Switch.scala 41:52:@30036.4]
  wire  output_36_55; // @[Switch.scala 41:38:@30037.4]
  wire  _T_68880; // @[Switch.scala 41:52:@30039.4]
  wire  output_36_56; // @[Switch.scala 41:38:@30040.4]
  wire  _T_68883; // @[Switch.scala 41:52:@30042.4]
  wire  output_36_57; // @[Switch.scala 41:38:@30043.4]
  wire  _T_68886; // @[Switch.scala 41:52:@30045.4]
  wire  output_36_58; // @[Switch.scala 41:38:@30046.4]
  wire  _T_68889; // @[Switch.scala 41:52:@30048.4]
  wire  output_36_59; // @[Switch.scala 41:38:@30049.4]
  wire  _T_68892; // @[Switch.scala 41:52:@30051.4]
  wire  output_36_60; // @[Switch.scala 41:38:@30052.4]
  wire  _T_68895; // @[Switch.scala 41:52:@30054.4]
  wire  output_36_61; // @[Switch.scala 41:38:@30055.4]
  wire  _T_68898; // @[Switch.scala 41:52:@30057.4]
  wire  output_36_62; // @[Switch.scala 41:38:@30058.4]
  wire  _T_68901; // @[Switch.scala 41:52:@30060.4]
  wire  output_36_63; // @[Switch.scala 41:38:@30061.4]
  wire [7:0] _T_68909; // @[Switch.scala 43:31:@30069.4]
  wire [15:0] _T_68917; // @[Switch.scala 43:31:@30077.4]
  wire [7:0] _T_68924; // @[Switch.scala 43:31:@30084.4]
  wire [31:0] _T_68933; // @[Switch.scala 43:31:@30093.4]
  wire [7:0] _T_68940; // @[Switch.scala 43:31:@30100.4]
  wire [15:0] _T_68948; // @[Switch.scala 43:31:@30108.4]
  wire [7:0] _T_68955; // @[Switch.scala 43:31:@30115.4]
  wire [31:0] _T_68964; // @[Switch.scala 43:31:@30124.4]
  wire [63:0] _T_68965; // @[Switch.scala 43:31:@30125.4]
  wire  _T_68969; // @[Switch.scala 41:52:@30128.4]
  wire  output_37_0; // @[Switch.scala 41:38:@30129.4]
  wire  _T_68972; // @[Switch.scala 41:52:@30131.4]
  wire  output_37_1; // @[Switch.scala 41:38:@30132.4]
  wire  _T_68975; // @[Switch.scala 41:52:@30134.4]
  wire  output_37_2; // @[Switch.scala 41:38:@30135.4]
  wire  _T_68978; // @[Switch.scala 41:52:@30137.4]
  wire  output_37_3; // @[Switch.scala 41:38:@30138.4]
  wire  _T_68981; // @[Switch.scala 41:52:@30140.4]
  wire  output_37_4; // @[Switch.scala 41:38:@30141.4]
  wire  _T_68984; // @[Switch.scala 41:52:@30143.4]
  wire  output_37_5; // @[Switch.scala 41:38:@30144.4]
  wire  _T_68987; // @[Switch.scala 41:52:@30146.4]
  wire  output_37_6; // @[Switch.scala 41:38:@30147.4]
  wire  _T_68990; // @[Switch.scala 41:52:@30149.4]
  wire  output_37_7; // @[Switch.scala 41:38:@30150.4]
  wire  _T_68993; // @[Switch.scala 41:52:@30152.4]
  wire  output_37_8; // @[Switch.scala 41:38:@30153.4]
  wire  _T_68996; // @[Switch.scala 41:52:@30155.4]
  wire  output_37_9; // @[Switch.scala 41:38:@30156.4]
  wire  _T_68999; // @[Switch.scala 41:52:@30158.4]
  wire  output_37_10; // @[Switch.scala 41:38:@30159.4]
  wire  _T_69002; // @[Switch.scala 41:52:@30161.4]
  wire  output_37_11; // @[Switch.scala 41:38:@30162.4]
  wire  _T_69005; // @[Switch.scala 41:52:@30164.4]
  wire  output_37_12; // @[Switch.scala 41:38:@30165.4]
  wire  _T_69008; // @[Switch.scala 41:52:@30167.4]
  wire  output_37_13; // @[Switch.scala 41:38:@30168.4]
  wire  _T_69011; // @[Switch.scala 41:52:@30170.4]
  wire  output_37_14; // @[Switch.scala 41:38:@30171.4]
  wire  _T_69014; // @[Switch.scala 41:52:@30173.4]
  wire  output_37_15; // @[Switch.scala 41:38:@30174.4]
  wire  _T_69017; // @[Switch.scala 41:52:@30176.4]
  wire  output_37_16; // @[Switch.scala 41:38:@30177.4]
  wire  _T_69020; // @[Switch.scala 41:52:@30179.4]
  wire  output_37_17; // @[Switch.scala 41:38:@30180.4]
  wire  _T_69023; // @[Switch.scala 41:52:@30182.4]
  wire  output_37_18; // @[Switch.scala 41:38:@30183.4]
  wire  _T_69026; // @[Switch.scala 41:52:@30185.4]
  wire  output_37_19; // @[Switch.scala 41:38:@30186.4]
  wire  _T_69029; // @[Switch.scala 41:52:@30188.4]
  wire  output_37_20; // @[Switch.scala 41:38:@30189.4]
  wire  _T_69032; // @[Switch.scala 41:52:@30191.4]
  wire  output_37_21; // @[Switch.scala 41:38:@30192.4]
  wire  _T_69035; // @[Switch.scala 41:52:@30194.4]
  wire  output_37_22; // @[Switch.scala 41:38:@30195.4]
  wire  _T_69038; // @[Switch.scala 41:52:@30197.4]
  wire  output_37_23; // @[Switch.scala 41:38:@30198.4]
  wire  _T_69041; // @[Switch.scala 41:52:@30200.4]
  wire  output_37_24; // @[Switch.scala 41:38:@30201.4]
  wire  _T_69044; // @[Switch.scala 41:52:@30203.4]
  wire  output_37_25; // @[Switch.scala 41:38:@30204.4]
  wire  _T_69047; // @[Switch.scala 41:52:@30206.4]
  wire  output_37_26; // @[Switch.scala 41:38:@30207.4]
  wire  _T_69050; // @[Switch.scala 41:52:@30209.4]
  wire  output_37_27; // @[Switch.scala 41:38:@30210.4]
  wire  _T_69053; // @[Switch.scala 41:52:@30212.4]
  wire  output_37_28; // @[Switch.scala 41:38:@30213.4]
  wire  _T_69056; // @[Switch.scala 41:52:@30215.4]
  wire  output_37_29; // @[Switch.scala 41:38:@30216.4]
  wire  _T_69059; // @[Switch.scala 41:52:@30218.4]
  wire  output_37_30; // @[Switch.scala 41:38:@30219.4]
  wire  _T_69062; // @[Switch.scala 41:52:@30221.4]
  wire  output_37_31; // @[Switch.scala 41:38:@30222.4]
  wire  _T_69065; // @[Switch.scala 41:52:@30224.4]
  wire  output_37_32; // @[Switch.scala 41:38:@30225.4]
  wire  _T_69068; // @[Switch.scala 41:52:@30227.4]
  wire  output_37_33; // @[Switch.scala 41:38:@30228.4]
  wire  _T_69071; // @[Switch.scala 41:52:@30230.4]
  wire  output_37_34; // @[Switch.scala 41:38:@30231.4]
  wire  _T_69074; // @[Switch.scala 41:52:@30233.4]
  wire  output_37_35; // @[Switch.scala 41:38:@30234.4]
  wire  _T_69077; // @[Switch.scala 41:52:@30236.4]
  wire  output_37_36; // @[Switch.scala 41:38:@30237.4]
  wire  _T_69080; // @[Switch.scala 41:52:@30239.4]
  wire  output_37_37; // @[Switch.scala 41:38:@30240.4]
  wire  _T_69083; // @[Switch.scala 41:52:@30242.4]
  wire  output_37_38; // @[Switch.scala 41:38:@30243.4]
  wire  _T_69086; // @[Switch.scala 41:52:@30245.4]
  wire  output_37_39; // @[Switch.scala 41:38:@30246.4]
  wire  _T_69089; // @[Switch.scala 41:52:@30248.4]
  wire  output_37_40; // @[Switch.scala 41:38:@30249.4]
  wire  _T_69092; // @[Switch.scala 41:52:@30251.4]
  wire  output_37_41; // @[Switch.scala 41:38:@30252.4]
  wire  _T_69095; // @[Switch.scala 41:52:@30254.4]
  wire  output_37_42; // @[Switch.scala 41:38:@30255.4]
  wire  _T_69098; // @[Switch.scala 41:52:@30257.4]
  wire  output_37_43; // @[Switch.scala 41:38:@30258.4]
  wire  _T_69101; // @[Switch.scala 41:52:@30260.4]
  wire  output_37_44; // @[Switch.scala 41:38:@30261.4]
  wire  _T_69104; // @[Switch.scala 41:52:@30263.4]
  wire  output_37_45; // @[Switch.scala 41:38:@30264.4]
  wire  _T_69107; // @[Switch.scala 41:52:@30266.4]
  wire  output_37_46; // @[Switch.scala 41:38:@30267.4]
  wire  _T_69110; // @[Switch.scala 41:52:@30269.4]
  wire  output_37_47; // @[Switch.scala 41:38:@30270.4]
  wire  _T_69113; // @[Switch.scala 41:52:@30272.4]
  wire  output_37_48; // @[Switch.scala 41:38:@30273.4]
  wire  _T_69116; // @[Switch.scala 41:52:@30275.4]
  wire  output_37_49; // @[Switch.scala 41:38:@30276.4]
  wire  _T_69119; // @[Switch.scala 41:52:@30278.4]
  wire  output_37_50; // @[Switch.scala 41:38:@30279.4]
  wire  _T_69122; // @[Switch.scala 41:52:@30281.4]
  wire  output_37_51; // @[Switch.scala 41:38:@30282.4]
  wire  _T_69125; // @[Switch.scala 41:52:@30284.4]
  wire  output_37_52; // @[Switch.scala 41:38:@30285.4]
  wire  _T_69128; // @[Switch.scala 41:52:@30287.4]
  wire  output_37_53; // @[Switch.scala 41:38:@30288.4]
  wire  _T_69131; // @[Switch.scala 41:52:@30290.4]
  wire  output_37_54; // @[Switch.scala 41:38:@30291.4]
  wire  _T_69134; // @[Switch.scala 41:52:@30293.4]
  wire  output_37_55; // @[Switch.scala 41:38:@30294.4]
  wire  _T_69137; // @[Switch.scala 41:52:@30296.4]
  wire  output_37_56; // @[Switch.scala 41:38:@30297.4]
  wire  _T_69140; // @[Switch.scala 41:52:@30299.4]
  wire  output_37_57; // @[Switch.scala 41:38:@30300.4]
  wire  _T_69143; // @[Switch.scala 41:52:@30302.4]
  wire  output_37_58; // @[Switch.scala 41:38:@30303.4]
  wire  _T_69146; // @[Switch.scala 41:52:@30305.4]
  wire  output_37_59; // @[Switch.scala 41:38:@30306.4]
  wire  _T_69149; // @[Switch.scala 41:52:@30308.4]
  wire  output_37_60; // @[Switch.scala 41:38:@30309.4]
  wire  _T_69152; // @[Switch.scala 41:52:@30311.4]
  wire  output_37_61; // @[Switch.scala 41:38:@30312.4]
  wire  _T_69155; // @[Switch.scala 41:52:@30314.4]
  wire  output_37_62; // @[Switch.scala 41:38:@30315.4]
  wire  _T_69158; // @[Switch.scala 41:52:@30317.4]
  wire  output_37_63; // @[Switch.scala 41:38:@30318.4]
  wire [7:0] _T_69166; // @[Switch.scala 43:31:@30326.4]
  wire [15:0] _T_69174; // @[Switch.scala 43:31:@30334.4]
  wire [7:0] _T_69181; // @[Switch.scala 43:31:@30341.4]
  wire [31:0] _T_69190; // @[Switch.scala 43:31:@30350.4]
  wire [7:0] _T_69197; // @[Switch.scala 43:31:@30357.4]
  wire [15:0] _T_69205; // @[Switch.scala 43:31:@30365.4]
  wire [7:0] _T_69212; // @[Switch.scala 43:31:@30372.4]
  wire [31:0] _T_69221; // @[Switch.scala 43:31:@30381.4]
  wire [63:0] _T_69222; // @[Switch.scala 43:31:@30382.4]
  wire  _T_69226; // @[Switch.scala 41:52:@30385.4]
  wire  output_38_0; // @[Switch.scala 41:38:@30386.4]
  wire  _T_69229; // @[Switch.scala 41:52:@30388.4]
  wire  output_38_1; // @[Switch.scala 41:38:@30389.4]
  wire  _T_69232; // @[Switch.scala 41:52:@30391.4]
  wire  output_38_2; // @[Switch.scala 41:38:@30392.4]
  wire  _T_69235; // @[Switch.scala 41:52:@30394.4]
  wire  output_38_3; // @[Switch.scala 41:38:@30395.4]
  wire  _T_69238; // @[Switch.scala 41:52:@30397.4]
  wire  output_38_4; // @[Switch.scala 41:38:@30398.4]
  wire  _T_69241; // @[Switch.scala 41:52:@30400.4]
  wire  output_38_5; // @[Switch.scala 41:38:@30401.4]
  wire  _T_69244; // @[Switch.scala 41:52:@30403.4]
  wire  output_38_6; // @[Switch.scala 41:38:@30404.4]
  wire  _T_69247; // @[Switch.scala 41:52:@30406.4]
  wire  output_38_7; // @[Switch.scala 41:38:@30407.4]
  wire  _T_69250; // @[Switch.scala 41:52:@30409.4]
  wire  output_38_8; // @[Switch.scala 41:38:@30410.4]
  wire  _T_69253; // @[Switch.scala 41:52:@30412.4]
  wire  output_38_9; // @[Switch.scala 41:38:@30413.4]
  wire  _T_69256; // @[Switch.scala 41:52:@30415.4]
  wire  output_38_10; // @[Switch.scala 41:38:@30416.4]
  wire  _T_69259; // @[Switch.scala 41:52:@30418.4]
  wire  output_38_11; // @[Switch.scala 41:38:@30419.4]
  wire  _T_69262; // @[Switch.scala 41:52:@30421.4]
  wire  output_38_12; // @[Switch.scala 41:38:@30422.4]
  wire  _T_69265; // @[Switch.scala 41:52:@30424.4]
  wire  output_38_13; // @[Switch.scala 41:38:@30425.4]
  wire  _T_69268; // @[Switch.scala 41:52:@30427.4]
  wire  output_38_14; // @[Switch.scala 41:38:@30428.4]
  wire  _T_69271; // @[Switch.scala 41:52:@30430.4]
  wire  output_38_15; // @[Switch.scala 41:38:@30431.4]
  wire  _T_69274; // @[Switch.scala 41:52:@30433.4]
  wire  output_38_16; // @[Switch.scala 41:38:@30434.4]
  wire  _T_69277; // @[Switch.scala 41:52:@30436.4]
  wire  output_38_17; // @[Switch.scala 41:38:@30437.4]
  wire  _T_69280; // @[Switch.scala 41:52:@30439.4]
  wire  output_38_18; // @[Switch.scala 41:38:@30440.4]
  wire  _T_69283; // @[Switch.scala 41:52:@30442.4]
  wire  output_38_19; // @[Switch.scala 41:38:@30443.4]
  wire  _T_69286; // @[Switch.scala 41:52:@30445.4]
  wire  output_38_20; // @[Switch.scala 41:38:@30446.4]
  wire  _T_69289; // @[Switch.scala 41:52:@30448.4]
  wire  output_38_21; // @[Switch.scala 41:38:@30449.4]
  wire  _T_69292; // @[Switch.scala 41:52:@30451.4]
  wire  output_38_22; // @[Switch.scala 41:38:@30452.4]
  wire  _T_69295; // @[Switch.scala 41:52:@30454.4]
  wire  output_38_23; // @[Switch.scala 41:38:@30455.4]
  wire  _T_69298; // @[Switch.scala 41:52:@30457.4]
  wire  output_38_24; // @[Switch.scala 41:38:@30458.4]
  wire  _T_69301; // @[Switch.scala 41:52:@30460.4]
  wire  output_38_25; // @[Switch.scala 41:38:@30461.4]
  wire  _T_69304; // @[Switch.scala 41:52:@30463.4]
  wire  output_38_26; // @[Switch.scala 41:38:@30464.4]
  wire  _T_69307; // @[Switch.scala 41:52:@30466.4]
  wire  output_38_27; // @[Switch.scala 41:38:@30467.4]
  wire  _T_69310; // @[Switch.scala 41:52:@30469.4]
  wire  output_38_28; // @[Switch.scala 41:38:@30470.4]
  wire  _T_69313; // @[Switch.scala 41:52:@30472.4]
  wire  output_38_29; // @[Switch.scala 41:38:@30473.4]
  wire  _T_69316; // @[Switch.scala 41:52:@30475.4]
  wire  output_38_30; // @[Switch.scala 41:38:@30476.4]
  wire  _T_69319; // @[Switch.scala 41:52:@30478.4]
  wire  output_38_31; // @[Switch.scala 41:38:@30479.4]
  wire  _T_69322; // @[Switch.scala 41:52:@30481.4]
  wire  output_38_32; // @[Switch.scala 41:38:@30482.4]
  wire  _T_69325; // @[Switch.scala 41:52:@30484.4]
  wire  output_38_33; // @[Switch.scala 41:38:@30485.4]
  wire  _T_69328; // @[Switch.scala 41:52:@30487.4]
  wire  output_38_34; // @[Switch.scala 41:38:@30488.4]
  wire  _T_69331; // @[Switch.scala 41:52:@30490.4]
  wire  output_38_35; // @[Switch.scala 41:38:@30491.4]
  wire  _T_69334; // @[Switch.scala 41:52:@30493.4]
  wire  output_38_36; // @[Switch.scala 41:38:@30494.4]
  wire  _T_69337; // @[Switch.scala 41:52:@30496.4]
  wire  output_38_37; // @[Switch.scala 41:38:@30497.4]
  wire  _T_69340; // @[Switch.scala 41:52:@30499.4]
  wire  output_38_38; // @[Switch.scala 41:38:@30500.4]
  wire  _T_69343; // @[Switch.scala 41:52:@30502.4]
  wire  output_38_39; // @[Switch.scala 41:38:@30503.4]
  wire  _T_69346; // @[Switch.scala 41:52:@30505.4]
  wire  output_38_40; // @[Switch.scala 41:38:@30506.4]
  wire  _T_69349; // @[Switch.scala 41:52:@30508.4]
  wire  output_38_41; // @[Switch.scala 41:38:@30509.4]
  wire  _T_69352; // @[Switch.scala 41:52:@30511.4]
  wire  output_38_42; // @[Switch.scala 41:38:@30512.4]
  wire  _T_69355; // @[Switch.scala 41:52:@30514.4]
  wire  output_38_43; // @[Switch.scala 41:38:@30515.4]
  wire  _T_69358; // @[Switch.scala 41:52:@30517.4]
  wire  output_38_44; // @[Switch.scala 41:38:@30518.4]
  wire  _T_69361; // @[Switch.scala 41:52:@30520.4]
  wire  output_38_45; // @[Switch.scala 41:38:@30521.4]
  wire  _T_69364; // @[Switch.scala 41:52:@30523.4]
  wire  output_38_46; // @[Switch.scala 41:38:@30524.4]
  wire  _T_69367; // @[Switch.scala 41:52:@30526.4]
  wire  output_38_47; // @[Switch.scala 41:38:@30527.4]
  wire  _T_69370; // @[Switch.scala 41:52:@30529.4]
  wire  output_38_48; // @[Switch.scala 41:38:@30530.4]
  wire  _T_69373; // @[Switch.scala 41:52:@30532.4]
  wire  output_38_49; // @[Switch.scala 41:38:@30533.4]
  wire  _T_69376; // @[Switch.scala 41:52:@30535.4]
  wire  output_38_50; // @[Switch.scala 41:38:@30536.4]
  wire  _T_69379; // @[Switch.scala 41:52:@30538.4]
  wire  output_38_51; // @[Switch.scala 41:38:@30539.4]
  wire  _T_69382; // @[Switch.scala 41:52:@30541.4]
  wire  output_38_52; // @[Switch.scala 41:38:@30542.4]
  wire  _T_69385; // @[Switch.scala 41:52:@30544.4]
  wire  output_38_53; // @[Switch.scala 41:38:@30545.4]
  wire  _T_69388; // @[Switch.scala 41:52:@30547.4]
  wire  output_38_54; // @[Switch.scala 41:38:@30548.4]
  wire  _T_69391; // @[Switch.scala 41:52:@30550.4]
  wire  output_38_55; // @[Switch.scala 41:38:@30551.4]
  wire  _T_69394; // @[Switch.scala 41:52:@30553.4]
  wire  output_38_56; // @[Switch.scala 41:38:@30554.4]
  wire  _T_69397; // @[Switch.scala 41:52:@30556.4]
  wire  output_38_57; // @[Switch.scala 41:38:@30557.4]
  wire  _T_69400; // @[Switch.scala 41:52:@30559.4]
  wire  output_38_58; // @[Switch.scala 41:38:@30560.4]
  wire  _T_69403; // @[Switch.scala 41:52:@30562.4]
  wire  output_38_59; // @[Switch.scala 41:38:@30563.4]
  wire  _T_69406; // @[Switch.scala 41:52:@30565.4]
  wire  output_38_60; // @[Switch.scala 41:38:@30566.4]
  wire  _T_69409; // @[Switch.scala 41:52:@30568.4]
  wire  output_38_61; // @[Switch.scala 41:38:@30569.4]
  wire  _T_69412; // @[Switch.scala 41:52:@30571.4]
  wire  output_38_62; // @[Switch.scala 41:38:@30572.4]
  wire  _T_69415; // @[Switch.scala 41:52:@30574.4]
  wire  output_38_63; // @[Switch.scala 41:38:@30575.4]
  wire [7:0] _T_69423; // @[Switch.scala 43:31:@30583.4]
  wire [15:0] _T_69431; // @[Switch.scala 43:31:@30591.4]
  wire [7:0] _T_69438; // @[Switch.scala 43:31:@30598.4]
  wire [31:0] _T_69447; // @[Switch.scala 43:31:@30607.4]
  wire [7:0] _T_69454; // @[Switch.scala 43:31:@30614.4]
  wire [15:0] _T_69462; // @[Switch.scala 43:31:@30622.4]
  wire [7:0] _T_69469; // @[Switch.scala 43:31:@30629.4]
  wire [31:0] _T_69478; // @[Switch.scala 43:31:@30638.4]
  wire [63:0] _T_69479; // @[Switch.scala 43:31:@30639.4]
  wire  _T_69483; // @[Switch.scala 41:52:@30642.4]
  wire  output_39_0; // @[Switch.scala 41:38:@30643.4]
  wire  _T_69486; // @[Switch.scala 41:52:@30645.4]
  wire  output_39_1; // @[Switch.scala 41:38:@30646.4]
  wire  _T_69489; // @[Switch.scala 41:52:@30648.4]
  wire  output_39_2; // @[Switch.scala 41:38:@30649.4]
  wire  _T_69492; // @[Switch.scala 41:52:@30651.4]
  wire  output_39_3; // @[Switch.scala 41:38:@30652.4]
  wire  _T_69495; // @[Switch.scala 41:52:@30654.4]
  wire  output_39_4; // @[Switch.scala 41:38:@30655.4]
  wire  _T_69498; // @[Switch.scala 41:52:@30657.4]
  wire  output_39_5; // @[Switch.scala 41:38:@30658.4]
  wire  _T_69501; // @[Switch.scala 41:52:@30660.4]
  wire  output_39_6; // @[Switch.scala 41:38:@30661.4]
  wire  _T_69504; // @[Switch.scala 41:52:@30663.4]
  wire  output_39_7; // @[Switch.scala 41:38:@30664.4]
  wire  _T_69507; // @[Switch.scala 41:52:@30666.4]
  wire  output_39_8; // @[Switch.scala 41:38:@30667.4]
  wire  _T_69510; // @[Switch.scala 41:52:@30669.4]
  wire  output_39_9; // @[Switch.scala 41:38:@30670.4]
  wire  _T_69513; // @[Switch.scala 41:52:@30672.4]
  wire  output_39_10; // @[Switch.scala 41:38:@30673.4]
  wire  _T_69516; // @[Switch.scala 41:52:@30675.4]
  wire  output_39_11; // @[Switch.scala 41:38:@30676.4]
  wire  _T_69519; // @[Switch.scala 41:52:@30678.4]
  wire  output_39_12; // @[Switch.scala 41:38:@30679.4]
  wire  _T_69522; // @[Switch.scala 41:52:@30681.4]
  wire  output_39_13; // @[Switch.scala 41:38:@30682.4]
  wire  _T_69525; // @[Switch.scala 41:52:@30684.4]
  wire  output_39_14; // @[Switch.scala 41:38:@30685.4]
  wire  _T_69528; // @[Switch.scala 41:52:@30687.4]
  wire  output_39_15; // @[Switch.scala 41:38:@30688.4]
  wire  _T_69531; // @[Switch.scala 41:52:@30690.4]
  wire  output_39_16; // @[Switch.scala 41:38:@30691.4]
  wire  _T_69534; // @[Switch.scala 41:52:@30693.4]
  wire  output_39_17; // @[Switch.scala 41:38:@30694.4]
  wire  _T_69537; // @[Switch.scala 41:52:@30696.4]
  wire  output_39_18; // @[Switch.scala 41:38:@30697.4]
  wire  _T_69540; // @[Switch.scala 41:52:@30699.4]
  wire  output_39_19; // @[Switch.scala 41:38:@30700.4]
  wire  _T_69543; // @[Switch.scala 41:52:@30702.4]
  wire  output_39_20; // @[Switch.scala 41:38:@30703.4]
  wire  _T_69546; // @[Switch.scala 41:52:@30705.4]
  wire  output_39_21; // @[Switch.scala 41:38:@30706.4]
  wire  _T_69549; // @[Switch.scala 41:52:@30708.4]
  wire  output_39_22; // @[Switch.scala 41:38:@30709.4]
  wire  _T_69552; // @[Switch.scala 41:52:@30711.4]
  wire  output_39_23; // @[Switch.scala 41:38:@30712.4]
  wire  _T_69555; // @[Switch.scala 41:52:@30714.4]
  wire  output_39_24; // @[Switch.scala 41:38:@30715.4]
  wire  _T_69558; // @[Switch.scala 41:52:@30717.4]
  wire  output_39_25; // @[Switch.scala 41:38:@30718.4]
  wire  _T_69561; // @[Switch.scala 41:52:@30720.4]
  wire  output_39_26; // @[Switch.scala 41:38:@30721.4]
  wire  _T_69564; // @[Switch.scala 41:52:@30723.4]
  wire  output_39_27; // @[Switch.scala 41:38:@30724.4]
  wire  _T_69567; // @[Switch.scala 41:52:@30726.4]
  wire  output_39_28; // @[Switch.scala 41:38:@30727.4]
  wire  _T_69570; // @[Switch.scala 41:52:@30729.4]
  wire  output_39_29; // @[Switch.scala 41:38:@30730.4]
  wire  _T_69573; // @[Switch.scala 41:52:@30732.4]
  wire  output_39_30; // @[Switch.scala 41:38:@30733.4]
  wire  _T_69576; // @[Switch.scala 41:52:@30735.4]
  wire  output_39_31; // @[Switch.scala 41:38:@30736.4]
  wire  _T_69579; // @[Switch.scala 41:52:@30738.4]
  wire  output_39_32; // @[Switch.scala 41:38:@30739.4]
  wire  _T_69582; // @[Switch.scala 41:52:@30741.4]
  wire  output_39_33; // @[Switch.scala 41:38:@30742.4]
  wire  _T_69585; // @[Switch.scala 41:52:@30744.4]
  wire  output_39_34; // @[Switch.scala 41:38:@30745.4]
  wire  _T_69588; // @[Switch.scala 41:52:@30747.4]
  wire  output_39_35; // @[Switch.scala 41:38:@30748.4]
  wire  _T_69591; // @[Switch.scala 41:52:@30750.4]
  wire  output_39_36; // @[Switch.scala 41:38:@30751.4]
  wire  _T_69594; // @[Switch.scala 41:52:@30753.4]
  wire  output_39_37; // @[Switch.scala 41:38:@30754.4]
  wire  _T_69597; // @[Switch.scala 41:52:@30756.4]
  wire  output_39_38; // @[Switch.scala 41:38:@30757.4]
  wire  _T_69600; // @[Switch.scala 41:52:@30759.4]
  wire  output_39_39; // @[Switch.scala 41:38:@30760.4]
  wire  _T_69603; // @[Switch.scala 41:52:@30762.4]
  wire  output_39_40; // @[Switch.scala 41:38:@30763.4]
  wire  _T_69606; // @[Switch.scala 41:52:@30765.4]
  wire  output_39_41; // @[Switch.scala 41:38:@30766.4]
  wire  _T_69609; // @[Switch.scala 41:52:@30768.4]
  wire  output_39_42; // @[Switch.scala 41:38:@30769.4]
  wire  _T_69612; // @[Switch.scala 41:52:@30771.4]
  wire  output_39_43; // @[Switch.scala 41:38:@30772.4]
  wire  _T_69615; // @[Switch.scala 41:52:@30774.4]
  wire  output_39_44; // @[Switch.scala 41:38:@30775.4]
  wire  _T_69618; // @[Switch.scala 41:52:@30777.4]
  wire  output_39_45; // @[Switch.scala 41:38:@30778.4]
  wire  _T_69621; // @[Switch.scala 41:52:@30780.4]
  wire  output_39_46; // @[Switch.scala 41:38:@30781.4]
  wire  _T_69624; // @[Switch.scala 41:52:@30783.4]
  wire  output_39_47; // @[Switch.scala 41:38:@30784.4]
  wire  _T_69627; // @[Switch.scala 41:52:@30786.4]
  wire  output_39_48; // @[Switch.scala 41:38:@30787.4]
  wire  _T_69630; // @[Switch.scala 41:52:@30789.4]
  wire  output_39_49; // @[Switch.scala 41:38:@30790.4]
  wire  _T_69633; // @[Switch.scala 41:52:@30792.4]
  wire  output_39_50; // @[Switch.scala 41:38:@30793.4]
  wire  _T_69636; // @[Switch.scala 41:52:@30795.4]
  wire  output_39_51; // @[Switch.scala 41:38:@30796.4]
  wire  _T_69639; // @[Switch.scala 41:52:@30798.4]
  wire  output_39_52; // @[Switch.scala 41:38:@30799.4]
  wire  _T_69642; // @[Switch.scala 41:52:@30801.4]
  wire  output_39_53; // @[Switch.scala 41:38:@30802.4]
  wire  _T_69645; // @[Switch.scala 41:52:@30804.4]
  wire  output_39_54; // @[Switch.scala 41:38:@30805.4]
  wire  _T_69648; // @[Switch.scala 41:52:@30807.4]
  wire  output_39_55; // @[Switch.scala 41:38:@30808.4]
  wire  _T_69651; // @[Switch.scala 41:52:@30810.4]
  wire  output_39_56; // @[Switch.scala 41:38:@30811.4]
  wire  _T_69654; // @[Switch.scala 41:52:@30813.4]
  wire  output_39_57; // @[Switch.scala 41:38:@30814.4]
  wire  _T_69657; // @[Switch.scala 41:52:@30816.4]
  wire  output_39_58; // @[Switch.scala 41:38:@30817.4]
  wire  _T_69660; // @[Switch.scala 41:52:@30819.4]
  wire  output_39_59; // @[Switch.scala 41:38:@30820.4]
  wire  _T_69663; // @[Switch.scala 41:52:@30822.4]
  wire  output_39_60; // @[Switch.scala 41:38:@30823.4]
  wire  _T_69666; // @[Switch.scala 41:52:@30825.4]
  wire  output_39_61; // @[Switch.scala 41:38:@30826.4]
  wire  _T_69669; // @[Switch.scala 41:52:@30828.4]
  wire  output_39_62; // @[Switch.scala 41:38:@30829.4]
  wire  _T_69672; // @[Switch.scala 41:52:@30831.4]
  wire  output_39_63; // @[Switch.scala 41:38:@30832.4]
  wire [7:0] _T_69680; // @[Switch.scala 43:31:@30840.4]
  wire [15:0] _T_69688; // @[Switch.scala 43:31:@30848.4]
  wire [7:0] _T_69695; // @[Switch.scala 43:31:@30855.4]
  wire [31:0] _T_69704; // @[Switch.scala 43:31:@30864.4]
  wire [7:0] _T_69711; // @[Switch.scala 43:31:@30871.4]
  wire [15:0] _T_69719; // @[Switch.scala 43:31:@30879.4]
  wire [7:0] _T_69726; // @[Switch.scala 43:31:@30886.4]
  wire [31:0] _T_69735; // @[Switch.scala 43:31:@30895.4]
  wire [63:0] _T_69736; // @[Switch.scala 43:31:@30896.4]
  wire  _T_69740; // @[Switch.scala 41:52:@30899.4]
  wire  output_40_0; // @[Switch.scala 41:38:@30900.4]
  wire  _T_69743; // @[Switch.scala 41:52:@30902.4]
  wire  output_40_1; // @[Switch.scala 41:38:@30903.4]
  wire  _T_69746; // @[Switch.scala 41:52:@30905.4]
  wire  output_40_2; // @[Switch.scala 41:38:@30906.4]
  wire  _T_69749; // @[Switch.scala 41:52:@30908.4]
  wire  output_40_3; // @[Switch.scala 41:38:@30909.4]
  wire  _T_69752; // @[Switch.scala 41:52:@30911.4]
  wire  output_40_4; // @[Switch.scala 41:38:@30912.4]
  wire  _T_69755; // @[Switch.scala 41:52:@30914.4]
  wire  output_40_5; // @[Switch.scala 41:38:@30915.4]
  wire  _T_69758; // @[Switch.scala 41:52:@30917.4]
  wire  output_40_6; // @[Switch.scala 41:38:@30918.4]
  wire  _T_69761; // @[Switch.scala 41:52:@30920.4]
  wire  output_40_7; // @[Switch.scala 41:38:@30921.4]
  wire  _T_69764; // @[Switch.scala 41:52:@30923.4]
  wire  output_40_8; // @[Switch.scala 41:38:@30924.4]
  wire  _T_69767; // @[Switch.scala 41:52:@30926.4]
  wire  output_40_9; // @[Switch.scala 41:38:@30927.4]
  wire  _T_69770; // @[Switch.scala 41:52:@30929.4]
  wire  output_40_10; // @[Switch.scala 41:38:@30930.4]
  wire  _T_69773; // @[Switch.scala 41:52:@30932.4]
  wire  output_40_11; // @[Switch.scala 41:38:@30933.4]
  wire  _T_69776; // @[Switch.scala 41:52:@30935.4]
  wire  output_40_12; // @[Switch.scala 41:38:@30936.4]
  wire  _T_69779; // @[Switch.scala 41:52:@30938.4]
  wire  output_40_13; // @[Switch.scala 41:38:@30939.4]
  wire  _T_69782; // @[Switch.scala 41:52:@30941.4]
  wire  output_40_14; // @[Switch.scala 41:38:@30942.4]
  wire  _T_69785; // @[Switch.scala 41:52:@30944.4]
  wire  output_40_15; // @[Switch.scala 41:38:@30945.4]
  wire  _T_69788; // @[Switch.scala 41:52:@30947.4]
  wire  output_40_16; // @[Switch.scala 41:38:@30948.4]
  wire  _T_69791; // @[Switch.scala 41:52:@30950.4]
  wire  output_40_17; // @[Switch.scala 41:38:@30951.4]
  wire  _T_69794; // @[Switch.scala 41:52:@30953.4]
  wire  output_40_18; // @[Switch.scala 41:38:@30954.4]
  wire  _T_69797; // @[Switch.scala 41:52:@30956.4]
  wire  output_40_19; // @[Switch.scala 41:38:@30957.4]
  wire  _T_69800; // @[Switch.scala 41:52:@30959.4]
  wire  output_40_20; // @[Switch.scala 41:38:@30960.4]
  wire  _T_69803; // @[Switch.scala 41:52:@30962.4]
  wire  output_40_21; // @[Switch.scala 41:38:@30963.4]
  wire  _T_69806; // @[Switch.scala 41:52:@30965.4]
  wire  output_40_22; // @[Switch.scala 41:38:@30966.4]
  wire  _T_69809; // @[Switch.scala 41:52:@30968.4]
  wire  output_40_23; // @[Switch.scala 41:38:@30969.4]
  wire  _T_69812; // @[Switch.scala 41:52:@30971.4]
  wire  output_40_24; // @[Switch.scala 41:38:@30972.4]
  wire  _T_69815; // @[Switch.scala 41:52:@30974.4]
  wire  output_40_25; // @[Switch.scala 41:38:@30975.4]
  wire  _T_69818; // @[Switch.scala 41:52:@30977.4]
  wire  output_40_26; // @[Switch.scala 41:38:@30978.4]
  wire  _T_69821; // @[Switch.scala 41:52:@30980.4]
  wire  output_40_27; // @[Switch.scala 41:38:@30981.4]
  wire  _T_69824; // @[Switch.scala 41:52:@30983.4]
  wire  output_40_28; // @[Switch.scala 41:38:@30984.4]
  wire  _T_69827; // @[Switch.scala 41:52:@30986.4]
  wire  output_40_29; // @[Switch.scala 41:38:@30987.4]
  wire  _T_69830; // @[Switch.scala 41:52:@30989.4]
  wire  output_40_30; // @[Switch.scala 41:38:@30990.4]
  wire  _T_69833; // @[Switch.scala 41:52:@30992.4]
  wire  output_40_31; // @[Switch.scala 41:38:@30993.4]
  wire  _T_69836; // @[Switch.scala 41:52:@30995.4]
  wire  output_40_32; // @[Switch.scala 41:38:@30996.4]
  wire  _T_69839; // @[Switch.scala 41:52:@30998.4]
  wire  output_40_33; // @[Switch.scala 41:38:@30999.4]
  wire  _T_69842; // @[Switch.scala 41:52:@31001.4]
  wire  output_40_34; // @[Switch.scala 41:38:@31002.4]
  wire  _T_69845; // @[Switch.scala 41:52:@31004.4]
  wire  output_40_35; // @[Switch.scala 41:38:@31005.4]
  wire  _T_69848; // @[Switch.scala 41:52:@31007.4]
  wire  output_40_36; // @[Switch.scala 41:38:@31008.4]
  wire  _T_69851; // @[Switch.scala 41:52:@31010.4]
  wire  output_40_37; // @[Switch.scala 41:38:@31011.4]
  wire  _T_69854; // @[Switch.scala 41:52:@31013.4]
  wire  output_40_38; // @[Switch.scala 41:38:@31014.4]
  wire  _T_69857; // @[Switch.scala 41:52:@31016.4]
  wire  output_40_39; // @[Switch.scala 41:38:@31017.4]
  wire  _T_69860; // @[Switch.scala 41:52:@31019.4]
  wire  output_40_40; // @[Switch.scala 41:38:@31020.4]
  wire  _T_69863; // @[Switch.scala 41:52:@31022.4]
  wire  output_40_41; // @[Switch.scala 41:38:@31023.4]
  wire  _T_69866; // @[Switch.scala 41:52:@31025.4]
  wire  output_40_42; // @[Switch.scala 41:38:@31026.4]
  wire  _T_69869; // @[Switch.scala 41:52:@31028.4]
  wire  output_40_43; // @[Switch.scala 41:38:@31029.4]
  wire  _T_69872; // @[Switch.scala 41:52:@31031.4]
  wire  output_40_44; // @[Switch.scala 41:38:@31032.4]
  wire  _T_69875; // @[Switch.scala 41:52:@31034.4]
  wire  output_40_45; // @[Switch.scala 41:38:@31035.4]
  wire  _T_69878; // @[Switch.scala 41:52:@31037.4]
  wire  output_40_46; // @[Switch.scala 41:38:@31038.4]
  wire  _T_69881; // @[Switch.scala 41:52:@31040.4]
  wire  output_40_47; // @[Switch.scala 41:38:@31041.4]
  wire  _T_69884; // @[Switch.scala 41:52:@31043.4]
  wire  output_40_48; // @[Switch.scala 41:38:@31044.4]
  wire  _T_69887; // @[Switch.scala 41:52:@31046.4]
  wire  output_40_49; // @[Switch.scala 41:38:@31047.4]
  wire  _T_69890; // @[Switch.scala 41:52:@31049.4]
  wire  output_40_50; // @[Switch.scala 41:38:@31050.4]
  wire  _T_69893; // @[Switch.scala 41:52:@31052.4]
  wire  output_40_51; // @[Switch.scala 41:38:@31053.4]
  wire  _T_69896; // @[Switch.scala 41:52:@31055.4]
  wire  output_40_52; // @[Switch.scala 41:38:@31056.4]
  wire  _T_69899; // @[Switch.scala 41:52:@31058.4]
  wire  output_40_53; // @[Switch.scala 41:38:@31059.4]
  wire  _T_69902; // @[Switch.scala 41:52:@31061.4]
  wire  output_40_54; // @[Switch.scala 41:38:@31062.4]
  wire  _T_69905; // @[Switch.scala 41:52:@31064.4]
  wire  output_40_55; // @[Switch.scala 41:38:@31065.4]
  wire  _T_69908; // @[Switch.scala 41:52:@31067.4]
  wire  output_40_56; // @[Switch.scala 41:38:@31068.4]
  wire  _T_69911; // @[Switch.scala 41:52:@31070.4]
  wire  output_40_57; // @[Switch.scala 41:38:@31071.4]
  wire  _T_69914; // @[Switch.scala 41:52:@31073.4]
  wire  output_40_58; // @[Switch.scala 41:38:@31074.4]
  wire  _T_69917; // @[Switch.scala 41:52:@31076.4]
  wire  output_40_59; // @[Switch.scala 41:38:@31077.4]
  wire  _T_69920; // @[Switch.scala 41:52:@31079.4]
  wire  output_40_60; // @[Switch.scala 41:38:@31080.4]
  wire  _T_69923; // @[Switch.scala 41:52:@31082.4]
  wire  output_40_61; // @[Switch.scala 41:38:@31083.4]
  wire  _T_69926; // @[Switch.scala 41:52:@31085.4]
  wire  output_40_62; // @[Switch.scala 41:38:@31086.4]
  wire  _T_69929; // @[Switch.scala 41:52:@31088.4]
  wire  output_40_63; // @[Switch.scala 41:38:@31089.4]
  wire [7:0] _T_69937; // @[Switch.scala 43:31:@31097.4]
  wire [15:0] _T_69945; // @[Switch.scala 43:31:@31105.4]
  wire [7:0] _T_69952; // @[Switch.scala 43:31:@31112.4]
  wire [31:0] _T_69961; // @[Switch.scala 43:31:@31121.4]
  wire [7:0] _T_69968; // @[Switch.scala 43:31:@31128.4]
  wire [15:0] _T_69976; // @[Switch.scala 43:31:@31136.4]
  wire [7:0] _T_69983; // @[Switch.scala 43:31:@31143.4]
  wire [31:0] _T_69992; // @[Switch.scala 43:31:@31152.4]
  wire [63:0] _T_69993; // @[Switch.scala 43:31:@31153.4]
  wire  _T_69997; // @[Switch.scala 41:52:@31156.4]
  wire  output_41_0; // @[Switch.scala 41:38:@31157.4]
  wire  _T_70000; // @[Switch.scala 41:52:@31159.4]
  wire  output_41_1; // @[Switch.scala 41:38:@31160.4]
  wire  _T_70003; // @[Switch.scala 41:52:@31162.4]
  wire  output_41_2; // @[Switch.scala 41:38:@31163.4]
  wire  _T_70006; // @[Switch.scala 41:52:@31165.4]
  wire  output_41_3; // @[Switch.scala 41:38:@31166.4]
  wire  _T_70009; // @[Switch.scala 41:52:@31168.4]
  wire  output_41_4; // @[Switch.scala 41:38:@31169.4]
  wire  _T_70012; // @[Switch.scala 41:52:@31171.4]
  wire  output_41_5; // @[Switch.scala 41:38:@31172.4]
  wire  _T_70015; // @[Switch.scala 41:52:@31174.4]
  wire  output_41_6; // @[Switch.scala 41:38:@31175.4]
  wire  _T_70018; // @[Switch.scala 41:52:@31177.4]
  wire  output_41_7; // @[Switch.scala 41:38:@31178.4]
  wire  _T_70021; // @[Switch.scala 41:52:@31180.4]
  wire  output_41_8; // @[Switch.scala 41:38:@31181.4]
  wire  _T_70024; // @[Switch.scala 41:52:@31183.4]
  wire  output_41_9; // @[Switch.scala 41:38:@31184.4]
  wire  _T_70027; // @[Switch.scala 41:52:@31186.4]
  wire  output_41_10; // @[Switch.scala 41:38:@31187.4]
  wire  _T_70030; // @[Switch.scala 41:52:@31189.4]
  wire  output_41_11; // @[Switch.scala 41:38:@31190.4]
  wire  _T_70033; // @[Switch.scala 41:52:@31192.4]
  wire  output_41_12; // @[Switch.scala 41:38:@31193.4]
  wire  _T_70036; // @[Switch.scala 41:52:@31195.4]
  wire  output_41_13; // @[Switch.scala 41:38:@31196.4]
  wire  _T_70039; // @[Switch.scala 41:52:@31198.4]
  wire  output_41_14; // @[Switch.scala 41:38:@31199.4]
  wire  _T_70042; // @[Switch.scala 41:52:@31201.4]
  wire  output_41_15; // @[Switch.scala 41:38:@31202.4]
  wire  _T_70045; // @[Switch.scala 41:52:@31204.4]
  wire  output_41_16; // @[Switch.scala 41:38:@31205.4]
  wire  _T_70048; // @[Switch.scala 41:52:@31207.4]
  wire  output_41_17; // @[Switch.scala 41:38:@31208.4]
  wire  _T_70051; // @[Switch.scala 41:52:@31210.4]
  wire  output_41_18; // @[Switch.scala 41:38:@31211.4]
  wire  _T_70054; // @[Switch.scala 41:52:@31213.4]
  wire  output_41_19; // @[Switch.scala 41:38:@31214.4]
  wire  _T_70057; // @[Switch.scala 41:52:@31216.4]
  wire  output_41_20; // @[Switch.scala 41:38:@31217.4]
  wire  _T_70060; // @[Switch.scala 41:52:@31219.4]
  wire  output_41_21; // @[Switch.scala 41:38:@31220.4]
  wire  _T_70063; // @[Switch.scala 41:52:@31222.4]
  wire  output_41_22; // @[Switch.scala 41:38:@31223.4]
  wire  _T_70066; // @[Switch.scala 41:52:@31225.4]
  wire  output_41_23; // @[Switch.scala 41:38:@31226.4]
  wire  _T_70069; // @[Switch.scala 41:52:@31228.4]
  wire  output_41_24; // @[Switch.scala 41:38:@31229.4]
  wire  _T_70072; // @[Switch.scala 41:52:@31231.4]
  wire  output_41_25; // @[Switch.scala 41:38:@31232.4]
  wire  _T_70075; // @[Switch.scala 41:52:@31234.4]
  wire  output_41_26; // @[Switch.scala 41:38:@31235.4]
  wire  _T_70078; // @[Switch.scala 41:52:@31237.4]
  wire  output_41_27; // @[Switch.scala 41:38:@31238.4]
  wire  _T_70081; // @[Switch.scala 41:52:@31240.4]
  wire  output_41_28; // @[Switch.scala 41:38:@31241.4]
  wire  _T_70084; // @[Switch.scala 41:52:@31243.4]
  wire  output_41_29; // @[Switch.scala 41:38:@31244.4]
  wire  _T_70087; // @[Switch.scala 41:52:@31246.4]
  wire  output_41_30; // @[Switch.scala 41:38:@31247.4]
  wire  _T_70090; // @[Switch.scala 41:52:@31249.4]
  wire  output_41_31; // @[Switch.scala 41:38:@31250.4]
  wire  _T_70093; // @[Switch.scala 41:52:@31252.4]
  wire  output_41_32; // @[Switch.scala 41:38:@31253.4]
  wire  _T_70096; // @[Switch.scala 41:52:@31255.4]
  wire  output_41_33; // @[Switch.scala 41:38:@31256.4]
  wire  _T_70099; // @[Switch.scala 41:52:@31258.4]
  wire  output_41_34; // @[Switch.scala 41:38:@31259.4]
  wire  _T_70102; // @[Switch.scala 41:52:@31261.4]
  wire  output_41_35; // @[Switch.scala 41:38:@31262.4]
  wire  _T_70105; // @[Switch.scala 41:52:@31264.4]
  wire  output_41_36; // @[Switch.scala 41:38:@31265.4]
  wire  _T_70108; // @[Switch.scala 41:52:@31267.4]
  wire  output_41_37; // @[Switch.scala 41:38:@31268.4]
  wire  _T_70111; // @[Switch.scala 41:52:@31270.4]
  wire  output_41_38; // @[Switch.scala 41:38:@31271.4]
  wire  _T_70114; // @[Switch.scala 41:52:@31273.4]
  wire  output_41_39; // @[Switch.scala 41:38:@31274.4]
  wire  _T_70117; // @[Switch.scala 41:52:@31276.4]
  wire  output_41_40; // @[Switch.scala 41:38:@31277.4]
  wire  _T_70120; // @[Switch.scala 41:52:@31279.4]
  wire  output_41_41; // @[Switch.scala 41:38:@31280.4]
  wire  _T_70123; // @[Switch.scala 41:52:@31282.4]
  wire  output_41_42; // @[Switch.scala 41:38:@31283.4]
  wire  _T_70126; // @[Switch.scala 41:52:@31285.4]
  wire  output_41_43; // @[Switch.scala 41:38:@31286.4]
  wire  _T_70129; // @[Switch.scala 41:52:@31288.4]
  wire  output_41_44; // @[Switch.scala 41:38:@31289.4]
  wire  _T_70132; // @[Switch.scala 41:52:@31291.4]
  wire  output_41_45; // @[Switch.scala 41:38:@31292.4]
  wire  _T_70135; // @[Switch.scala 41:52:@31294.4]
  wire  output_41_46; // @[Switch.scala 41:38:@31295.4]
  wire  _T_70138; // @[Switch.scala 41:52:@31297.4]
  wire  output_41_47; // @[Switch.scala 41:38:@31298.4]
  wire  _T_70141; // @[Switch.scala 41:52:@31300.4]
  wire  output_41_48; // @[Switch.scala 41:38:@31301.4]
  wire  _T_70144; // @[Switch.scala 41:52:@31303.4]
  wire  output_41_49; // @[Switch.scala 41:38:@31304.4]
  wire  _T_70147; // @[Switch.scala 41:52:@31306.4]
  wire  output_41_50; // @[Switch.scala 41:38:@31307.4]
  wire  _T_70150; // @[Switch.scala 41:52:@31309.4]
  wire  output_41_51; // @[Switch.scala 41:38:@31310.4]
  wire  _T_70153; // @[Switch.scala 41:52:@31312.4]
  wire  output_41_52; // @[Switch.scala 41:38:@31313.4]
  wire  _T_70156; // @[Switch.scala 41:52:@31315.4]
  wire  output_41_53; // @[Switch.scala 41:38:@31316.4]
  wire  _T_70159; // @[Switch.scala 41:52:@31318.4]
  wire  output_41_54; // @[Switch.scala 41:38:@31319.4]
  wire  _T_70162; // @[Switch.scala 41:52:@31321.4]
  wire  output_41_55; // @[Switch.scala 41:38:@31322.4]
  wire  _T_70165; // @[Switch.scala 41:52:@31324.4]
  wire  output_41_56; // @[Switch.scala 41:38:@31325.4]
  wire  _T_70168; // @[Switch.scala 41:52:@31327.4]
  wire  output_41_57; // @[Switch.scala 41:38:@31328.4]
  wire  _T_70171; // @[Switch.scala 41:52:@31330.4]
  wire  output_41_58; // @[Switch.scala 41:38:@31331.4]
  wire  _T_70174; // @[Switch.scala 41:52:@31333.4]
  wire  output_41_59; // @[Switch.scala 41:38:@31334.4]
  wire  _T_70177; // @[Switch.scala 41:52:@31336.4]
  wire  output_41_60; // @[Switch.scala 41:38:@31337.4]
  wire  _T_70180; // @[Switch.scala 41:52:@31339.4]
  wire  output_41_61; // @[Switch.scala 41:38:@31340.4]
  wire  _T_70183; // @[Switch.scala 41:52:@31342.4]
  wire  output_41_62; // @[Switch.scala 41:38:@31343.4]
  wire  _T_70186; // @[Switch.scala 41:52:@31345.4]
  wire  output_41_63; // @[Switch.scala 41:38:@31346.4]
  wire [7:0] _T_70194; // @[Switch.scala 43:31:@31354.4]
  wire [15:0] _T_70202; // @[Switch.scala 43:31:@31362.4]
  wire [7:0] _T_70209; // @[Switch.scala 43:31:@31369.4]
  wire [31:0] _T_70218; // @[Switch.scala 43:31:@31378.4]
  wire [7:0] _T_70225; // @[Switch.scala 43:31:@31385.4]
  wire [15:0] _T_70233; // @[Switch.scala 43:31:@31393.4]
  wire [7:0] _T_70240; // @[Switch.scala 43:31:@31400.4]
  wire [31:0] _T_70249; // @[Switch.scala 43:31:@31409.4]
  wire [63:0] _T_70250; // @[Switch.scala 43:31:@31410.4]
  wire  _T_70254; // @[Switch.scala 41:52:@31413.4]
  wire  output_42_0; // @[Switch.scala 41:38:@31414.4]
  wire  _T_70257; // @[Switch.scala 41:52:@31416.4]
  wire  output_42_1; // @[Switch.scala 41:38:@31417.4]
  wire  _T_70260; // @[Switch.scala 41:52:@31419.4]
  wire  output_42_2; // @[Switch.scala 41:38:@31420.4]
  wire  _T_70263; // @[Switch.scala 41:52:@31422.4]
  wire  output_42_3; // @[Switch.scala 41:38:@31423.4]
  wire  _T_70266; // @[Switch.scala 41:52:@31425.4]
  wire  output_42_4; // @[Switch.scala 41:38:@31426.4]
  wire  _T_70269; // @[Switch.scala 41:52:@31428.4]
  wire  output_42_5; // @[Switch.scala 41:38:@31429.4]
  wire  _T_70272; // @[Switch.scala 41:52:@31431.4]
  wire  output_42_6; // @[Switch.scala 41:38:@31432.4]
  wire  _T_70275; // @[Switch.scala 41:52:@31434.4]
  wire  output_42_7; // @[Switch.scala 41:38:@31435.4]
  wire  _T_70278; // @[Switch.scala 41:52:@31437.4]
  wire  output_42_8; // @[Switch.scala 41:38:@31438.4]
  wire  _T_70281; // @[Switch.scala 41:52:@31440.4]
  wire  output_42_9; // @[Switch.scala 41:38:@31441.4]
  wire  _T_70284; // @[Switch.scala 41:52:@31443.4]
  wire  output_42_10; // @[Switch.scala 41:38:@31444.4]
  wire  _T_70287; // @[Switch.scala 41:52:@31446.4]
  wire  output_42_11; // @[Switch.scala 41:38:@31447.4]
  wire  _T_70290; // @[Switch.scala 41:52:@31449.4]
  wire  output_42_12; // @[Switch.scala 41:38:@31450.4]
  wire  _T_70293; // @[Switch.scala 41:52:@31452.4]
  wire  output_42_13; // @[Switch.scala 41:38:@31453.4]
  wire  _T_70296; // @[Switch.scala 41:52:@31455.4]
  wire  output_42_14; // @[Switch.scala 41:38:@31456.4]
  wire  _T_70299; // @[Switch.scala 41:52:@31458.4]
  wire  output_42_15; // @[Switch.scala 41:38:@31459.4]
  wire  _T_70302; // @[Switch.scala 41:52:@31461.4]
  wire  output_42_16; // @[Switch.scala 41:38:@31462.4]
  wire  _T_70305; // @[Switch.scala 41:52:@31464.4]
  wire  output_42_17; // @[Switch.scala 41:38:@31465.4]
  wire  _T_70308; // @[Switch.scala 41:52:@31467.4]
  wire  output_42_18; // @[Switch.scala 41:38:@31468.4]
  wire  _T_70311; // @[Switch.scala 41:52:@31470.4]
  wire  output_42_19; // @[Switch.scala 41:38:@31471.4]
  wire  _T_70314; // @[Switch.scala 41:52:@31473.4]
  wire  output_42_20; // @[Switch.scala 41:38:@31474.4]
  wire  _T_70317; // @[Switch.scala 41:52:@31476.4]
  wire  output_42_21; // @[Switch.scala 41:38:@31477.4]
  wire  _T_70320; // @[Switch.scala 41:52:@31479.4]
  wire  output_42_22; // @[Switch.scala 41:38:@31480.4]
  wire  _T_70323; // @[Switch.scala 41:52:@31482.4]
  wire  output_42_23; // @[Switch.scala 41:38:@31483.4]
  wire  _T_70326; // @[Switch.scala 41:52:@31485.4]
  wire  output_42_24; // @[Switch.scala 41:38:@31486.4]
  wire  _T_70329; // @[Switch.scala 41:52:@31488.4]
  wire  output_42_25; // @[Switch.scala 41:38:@31489.4]
  wire  _T_70332; // @[Switch.scala 41:52:@31491.4]
  wire  output_42_26; // @[Switch.scala 41:38:@31492.4]
  wire  _T_70335; // @[Switch.scala 41:52:@31494.4]
  wire  output_42_27; // @[Switch.scala 41:38:@31495.4]
  wire  _T_70338; // @[Switch.scala 41:52:@31497.4]
  wire  output_42_28; // @[Switch.scala 41:38:@31498.4]
  wire  _T_70341; // @[Switch.scala 41:52:@31500.4]
  wire  output_42_29; // @[Switch.scala 41:38:@31501.4]
  wire  _T_70344; // @[Switch.scala 41:52:@31503.4]
  wire  output_42_30; // @[Switch.scala 41:38:@31504.4]
  wire  _T_70347; // @[Switch.scala 41:52:@31506.4]
  wire  output_42_31; // @[Switch.scala 41:38:@31507.4]
  wire  _T_70350; // @[Switch.scala 41:52:@31509.4]
  wire  output_42_32; // @[Switch.scala 41:38:@31510.4]
  wire  _T_70353; // @[Switch.scala 41:52:@31512.4]
  wire  output_42_33; // @[Switch.scala 41:38:@31513.4]
  wire  _T_70356; // @[Switch.scala 41:52:@31515.4]
  wire  output_42_34; // @[Switch.scala 41:38:@31516.4]
  wire  _T_70359; // @[Switch.scala 41:52:@31518.4]
  wire  output_42_35; // @[Switch.scala 41:38:@31519.4]
  wire  _T_70362; // @[Switch.scala 41:52:@31521.4]
  wire  output_42_36; // @[Switch.scala 41:38:@31522.4]
  wire  _T_70365; // @[Switch.scala 41:52:@31524.4]
  wire  output_42_37; // @[Switch.scala 41:38:@31525.4]
  wire  _T_70368; // @[Switch.scala 41:52:@31527.4]
  wire  output_42_38; // @[Switch.scala 41:38:@31528.4]
  wire  _T_70371; // @[Switch.scala 41:52:@31530.4]
  wire  output_42_39; // @[Switch.scala 41:38:@31531.4]
  wire  _T_70374; // @[Switch.scala 41:52:@31533.4]
  wire  output_42_40; // @[Switch.scala 41:38:@31534.4]
  wire  _T_70377; // @[Switch.scala 41:52:@31536.4]
  wire  output_42_41; // @[Switch.scala 41:38:@31537.4]
  wire  _T_70380; // @[Switch.scala 41:52:@31539.4]
  wire  output_42_42; // @[Switch.scala 41:38:@31540.4]
  wire  _T_70383; // @[Switch.scala 41:52:@31542.4]
  wire  output_42_43; // @[Switch.scala 41:38:@31543.4]
  wire  _T_70386; // @[Switch.scala 41:52:@31545.4]
  wire  output_42_44; // @[Switch.scala 41:38:@31546.4]
  wire  _T_70389; // @[Switch.scala 41:52:@31548.4]
  wire  output_42_45; // @[Switch.scala 41:38:@31549.4]
  wire  _T_70392; // @[Switch.scala 41:52:@31551.4]
  wire  output_42_46; // @[Switch.scala 41:38:@31552.4]
  wire  _T_70395; // @[Switch.scala 41:52:@31554.4]
  wire  output_42_47; // @[Switch.scala 41:38:@31555.4]
  wire  _T_70398; // @[Switch.scala 41:52:@31557.4]
  wire  output_42_48; // @[Switch.scala 41:38:@31558.4]
  wire  _T_70401; // @[Switch.scala 41:52:@31560.4]
  wire  output_42_49; // @[Switch.scala 41:38:@31561.4]
  wire  _T_70404; // @[Switch.scala 41:52:@31563.4]
  wire  output_42_50; // @[Switch.scala 41:38:@31564.4]
  wire  _T_70407; // @[Switch.scala 41:52:@31566.4]
  wire  output_42_51; // @[Switch.scala 41:38:@31567.4]
  wire  _T_70410; // @[Switch.scala 41:52:@31569.4]
  wire  output_42_52; // @[Switch.scala 41:38:@31570.4]
  wire  _T_70413; // @[Switch.scala 41:52:@31572.4]
  wire  output_42_53; // @[Switch.scala 41:38:@31573.4]
  wire  _T_70416; // @[Switch.scala 41:52:@31575.4]
  wire  output_42_54; // @[Switch.scala 41:38:@31576.4]
  wire  _T_70419; // @[Switch.scala 41:52:@31578.4]
  wire  output_42_55; // @[Switch.scala 41:38:@31579.4]
  wire  _T_70422; // @[Switch.scala 41:52:@31581.4]
  wire  output_42_56; // @[Switch.scala 41:38:@31582.4]
  wire  _T_70425; // @[Switch.scala 41:52:@31584.4]
  wire  output_42_57; // @[Switch.scala 41:38:@31585.4]
  wire  _T_70428; // @[Switch.scala 41:52:@31587.4]
  wire  output_42_58; // @[Switch.scala 41:38:@31588.4]
  wire  _T_70431; // @[Switch.scala 41:52:@31590.4]
  wire  output_42_59; // @[Switch.scala 41:38:@31591.4]
  wire  _T_70434; // @[Switch.scala 41:52:@31593.4]
  wire  output_42_60; // @[Switch.scala 41:38:@31594.4]
  wire  _T_70437; // @[Switch.scala 41:52:@31596.4]
  wire  output_42_61; // @[Switch.scala 41:38:@31597.4]
  wire  _T_70440; // @[Switch.scala 41:52:@31599.4]
  wire  output_42_62; // @[Switch.scala 41:38:@31600.4]
  wire  _T_70443; // @[Switch.scala 41:52:@31602.4]
  wire  output_42_63; // @[Switch.scala 41:38:@31603.4]
  wire [7:0] _T_70451; // @[Switch.scala 43:31:@31611.4]
  wire [15:0] _T_70459; // @[Switch.scala 43:31:@31619.4]
  wire [7:0] _T_70466; // @[Switch.scala 43:31:@31626.4]
  wire [31:0] _T_70475; // @[Switch.scala 43:31:@31635.4]
  wire [7:0] _T_70482; // @[Switch.scala 43:31:@31642.4]
  wire [15:0] _T_70490; // @[Switch.scala 43:31:@31650.4]
  wire [7:0] _T_70497; // @[Switch.scala 43:31:@31657.4]
  wire [31:0] _T_70506; // @[Switch.scala 43:31:@31666.4]
  wire [63:0] _T_70507; // @[Switch.scala 43:31:@31667.4]
  wire  _T_70511; // @[Switch.scala 41:52:@31670.4]
  wire  output_43_0; // @[Switch.scala 41:38:@31671.4]
  wire  _T_70514; // @[Switch.scala 41:52:@31673.4]
  wire  output_43_1; // @[Switch.scala 41:38:@31674.4]
  wire  _T_70517; // @[Switch.scala 41:52:@31676.4]
  wire  output_43_2; // @[Switch.scala 41:38:@31677.4]
  wire  _T_70520; // @[Switch.scala 41:52:@31679.4]
  wire  output_43_3; // @[Switch.scala 41:38:@31680.4]
  wire  _T_70523; // @[Switch.scala 41:52:@31682.4]
  wire  output_43_4; // @[Switch.scala 41:38:@31683.4]
  wire  _T_70526; // @[Switch.scala 41:52:@31685.4]
  wire  output_43_5; // @[Switch.scala 41:38:@31686.4]
  wire  _T_70529; // @[Switch.scala 41:52:@31688.4]
  wire  output_43_6; // @[Switch.scala 41:38:@31689.4]
  wire  _T_70532; // @[Switch.scala 41:52:@31691.4]
  wire  output_43_7; // @[Switch.scala 41:38:@31692.4]
  wire  _T_70535; // @[Switch.scala 41:52:@31694.4]
  wire  output_43_8; // @[Switch.scala 41:38:@31695.4]
  wire  _T_70538; // @[Switch.scala 41:52:@31697.4]
  wire  output_43_9; // @[Switch.scala 41:38:@31698.4]
  wire  _T_70541; // @[Switch.scala 41:52:@31700.4]
  wire  output_43_10; // @[Switch.scala 41:38:@31701.4]
  wire  _T_70544; // @[Switch.scala 41:52:@31703.4]
  wire  output_43_11; // @[Switch.scala 41:38:@31704.4]
  wire  _T_70547; // @[Switch.scala 41:52:@31706.4]
  wire  output_43_12; // @[Switch.scala 41:38:@31707.4]
  wire  _T_70550; // @[Switch.scala 41:52:@31709.4]
  wire  output_43_13; // @[Switch.scala 41:38:@31710.4]
  wire  _T_70553; // @[Switch.scala 41:52:@31712.4]
  wire  output_43_14; // @[Switch.scala 41:38:@31713.4]
  wire  _T_70556; // @[Switch.scala 41:52:@31715.4]
  wire  output_43_15; // @[Switch.scala 41:38:@31716.4]
  wire  _T_70559; // @[Switch.scala 41:52:@31718.4]
  wire  output_43_16; // @[Switch.scala 41:38:@31719.4]
  wire  _T_70562; // @[Switch.scala 41:52:@31721.4]
  wire  output_43_17; // @[Switch.scala 41:38:@31722.4]
  wire  _T_70565; // @[Switch.scala 41:52:@31724.4]
  wire  output_43_18; // @[Switch.scala 41:38:@31725.4]
  wire  _T_70568; // @[Switch.scala 41:52:@31727.4]
  wire  output_43_19; // @[Switch.scala 41:38:@31728.4]
  wire  _T_70571; // @[Switch.scala 41:52:@31730.4]
  wire  output_43_20; // @[Switch.scala 41:38:@31731.4]
  wire  _T_70574; // @[Switch.scala 41:52:@31733.4]
  wire  output_43_21; // @[Switch.scala 41:38:@31734.4]
  wire  _T_70577; // @[Switch.scala 41:52:@31736.4]
  wire  output_43_22; // @[Switch.scala 41:38:@31737.4]
  wire  _T_70580; // @[Switch.scala 41:52:@31739.4]
  wire  output_43_23; // @[Switch.scala 41:38:@31740.4]
  wire  _T_70583; // @[Switch.scala 41:52:@31742.4]
  wire  output_43_24; // @[Switch.scala 41:38:@31743.4]
  wire  _T_70586; // @[Switch.scala 41:52:@31745.4]
  wire  output_43_25; // @[Switch.scala 41:38:@31746.4]
  wire  _T_70589; // @[Switch.scala 41:52:@31748.4]
  wire  output_43_26; // @[Switch.scala 41:38:@31749.4]
  wire  _T_70592; // @[Switch.scala 41:52:@31751.4]
  wire  output_43_27; // @[Switch.scala 41:38:@31752.4]
  wire  _T_70595; // @[Switch.scala 41:52:@31754.4]
  wire  output_43_28; // @[Switch.scala 41:38:@31755.4]
  wire  _T_70598; // @[Switch.scala 41:52:@31757.4]
  wire  output_43_29; // @[Switch.scala 41:38:@31758.4]
  wire  _T_70601; // @[Switch.scala 41:52:@31760.4]
  wire  output_43_30; // @[Switch.scala 41:38:@31761.4]
  wire  _T_70604; // @[Switch.scala 41:52:@31763.4]
  wire  output_43_31; // @[Switch.scala 41:38:@31764.4]
  wire  _T_70607; // @[Switch.scala 41:52:@31766.4]
  wire  output_43_32; // @[Switch.scala 41:38:@31767.4]
  wire  _T_70610; // @[Switch.scala 41:52:@31769.4]
  wire  output_43_33; // @[Switch.scala 41:38:@31770.4]
  wire  _T_70613; // @[Switch.scala 41:52:@31772.4]
  wire  output_43_34; // @[Switch.scala 41:38:@31773.4]
  wire  _T_70616; // @[Switch.scala 41:52:@31775.4]
  wire  output_43_35; // @[Switch.scala 41:38:@31776.4]
  wire  _T_70619; // @[Switch.scala 41:52:@31778.4]
  wire  output_43_36; // @[Switch.scala 41:38:@31779.4]
  wire  _T_70622; // @[Switch.scala 41:52:@31781.4]
  wire  output_43_37; // @[Switch.scala 41:38:@31782.4]
  wire  _T_70625; // @[Switch.scala 41:52:@31784.4]
  wire  output_43_38; // @[Switch.scala 41:38:@31785.4]
  wire  _T_70628; // @[Switch.scala 41:52:@31787.4]
  wire  output_43_39; // @[Switch.scala 41:38:@31788.4]
  wire  _T_70631; // @[Switch.scala 41:52:@31790.4]
  wire  output_43_40; // @[Switch.scala 41:38:@31791.4]
  wire  _T_70634; // @[Switch.scala 41:52:@31793.4]
  wire  output_43_41; // @[Switch.scala 41:38:@31794.4]
  wire  _T_70637; // @[Switch.scala 41:52:@31796.4]
  wire  output_43_42; // @[Switch.scala 41:38:@31797.4]
  wire  _T_70640; // @[Switch.scala 41:52:@31799.4]
  wire  output_43_43; // @[Switch.scala 41:38:@31800.4]
  wire  _T_70643; // @[Switch.scala 41:52:@31802.4]
  wire  output_43_44; // @[Switch.scala 41:38:@31803.4]
  wire  _T_70646; // @[Switch.scala 41:52:@31805.4]
  wire  output_43_45; // @[Switch.scala 41:38:@31806.4]
  wire  _T_70649; // @[Switch.scala 41:52:@31808.4]
  wire  output_43_46; // @[Switch.scala 41:38:@31809.4]
  wire  _T_70652; // @[Switch.scala 41:52:@31811.4]
  wire  output_43_47; // @[Switch.scala 41:38:@31812.4]
  wire  _T_70655; // @[Switch.scala 41:52:@31814.4]
  wire  output_43_48; // @[Switch.scala 41:38:@31815.4]
  wire  _T_70658; // @[Switch.scala 41:52:@31817.4]
  wire  output_43_49; // @[Switch.scala 41:38:@31818.4]
  wire  _T_70661; // @[Switch.scala 41:52:@31820.4]
  wire  output_43_50; // @[Switch.scala 41:38:@31821.4]
  wire  _T_70664; // @[Switch.scala 41:52:@31823.4]
  wire  output_43_51; // @[Switch.scala 41:38:@31824.4]
  wire  _T_70667; // @[Switch.scala 41:52:@31826.4]
  wire  output_43_52; // @[Switch.scala 41:38:@31827.4]
  wire  _T_70670; // @[Switch.scala 41:52:@31829.4]
  wire  output_43_53; // @[Switch.scala 41:38:@31830.4]
  wire  _T_70673; // @[Switch.scala 41:52:@31832.4]
  wire  output_43_54; // @[Switch.scala 41:38:@31833.4]
  wire  _T_70676; // @[Switch.scala 41:52:@31835.4]
  wire  output_43_55; // @[Switch.scala 41:38:@31836.4]
  wire  _T_70679; // @[Switch.scala 41:52:@31838.4]
  wire  output_43_56; // @[Switch.scala 41:38:@31839.4]
  wire  _T_70682; // @[Switch.scala 41:52:@31841.4]
  wire  output_43_57; // @[Switch.scala 41:38:@31842.4]
  wire  _T_70685; // @[Switch.scala 41:52:@31844.4]
  wire  output_43_58; // @[Switch.scala 41:38:@31845.4]
  wire  _T_70688; // @[Switch.scala 41:52:@31847.4]
  wire  output_43_59; // @[Switch.scala 41:38:@31848.4]
  wire  _T_70691; // @[Switch.scala 41:52:@31850.4]
  wire  output_43_60; // @[Switch.scala 41:38:@31851.4]
  wire  _T_70694; // @[Switch.scala 41:52:@31853.4]
  wire  output_43_61; // @[Switch.scala 41:38:@31854.4]
  wire  _T_70697; // @[Switch.scala 41:52:@31856.4]
  wire  output_43_62; // @[Switch.scala 41:38:@31857.4]
  wire  _T_70700; // @[Switch.scala 41:52:@31859.4]
  wire  output_43_63; // @[Switch.scala 41:38:@31860.4]
  wire [7:0] _T_70708; // @[Switch.scala 43:31:@31868.4]
  wire [15:0] _T_70716; // @[Switch.scala 43:31:@31876.4]
  wire [7:0] _T_70723; // @[Switch.scala 43:31:@31883.4]
  wire [31:0] _T_70732; // @[Switch.scala 43:31:@31892.4]
  wire [7:0] _T_70739; // @[Switch.scala 43:31:@31899.4]
  wire [15:0] _T_70747; // @[Switch.scala 43:31:@31907.4]
  wire [7:0] _T_70754; // @[Switch.scala 43:31:@31914.4]
  wire [31:0] _T_70763; // @[Switch.scala 43:31:@31923.4]
  wire [63:0] _T_70764; // @[Switch.scala 43:31:@31924.4]
  wire  _T_70768; // @[Switch.scala 41:52:@31927.4]
  wire  output_44_0; // @[Switch.scala 41:38:@31928.4]
  wire  _T_70771; // @[Switch.scala 41:52:@31930.4]
  wire  output_44_1; // @[Switch.scala 41:38:@31931.4]
  wire  _T_70774; // @[Switch.scala 41:52:@31933.4]
  wire  output_44_2; // @[Switch.scala 41:38:@31934.4]
  wire  _T_70777; // @[Switch.scala 41:52:@31936.4]
  wire  output_44_3; // @[Switch.scala 41:38:@31937.4]
  wire  _T_70780; // @[Switch.scala 41:52:@31939.4]
  wire  output_44_4; // @[Switch.scala 41:38:@31940.4]
  wire  _T_70783; // @[Switch.scala 41:52:@31942.4]
  wire  output_44_5; // @[Switch.scala 41:38:@31943.4]
  wire  _T_70786; // @[Switch.scala 41:52:@31945.4]
  wire  output_44_6; // @[Switch.scala 41:38:@31946.4]
  wire  _T_70789; // @[Switch.scala 41:52:@31948.4]
  wire  output_44_7; // @[Switch.scala 41:38:@31949.4]
  wire  _T_70792; // @[Switch.scala 41:52:@31951.4]
  wire  output_44_8; // @[Switch.scala 41:38:@31952.4]
  wire  _T_70795; // @[Switch.scala 41:52:@31954.4]
  wire  output_44_9; // @[Switch.scala 41:38:@31955.4]
  wire  _T_70798; // @[Switch.scala 41:52:@31957.4]
  wire  output_44_10; // @[Switch.scala 41:38:@31958.4]
  wire  _T_70801; // @[Switch.scala 41:52:@31960.4]
  wire  output_44_11; // @[Switch.scala 41:38:@31961.4]
  wire  _T_70804; // @[Switch.scala 41:52:@31963.4]
  wire  output_44_12; // @[Switch.scala 41:38:@31964.4]
  wire  _T_70807; // @[Switch.scala 41:52:@31966.4]
  wire  output_44_13; // @[Switch.scala 41:38:@31967.4]
  wire  _T_70810; // @[Switch.scala 41:52:@31969.4]
  wire  output_44_14; // @[Switch.scala 41:38:@31970.4]
  wire  _T_70813; // @[Switch.scala 41:52:@31972.4]
  wire  output_44_15; // @[Switch.scala 41:38:@31973.4]
  wire  _T_70816; // @[Switch.scala 41:52:@31975.4]
  wire  output_44_16; // @[Switch.scala 41:38:@31976.4]
  wire  _T_70819; // @[Switch.scala 41:52:@31978.4]
  wire  output_44_17; // @[Switch.scala 41:38:@31979.4]
  wire  _T_70822; // @[Switch.scala 41:52:@31981.4]
  wire  output_44_18; // @[Switch.scala 41:38:@31982.4]
  wire  _T_70825; // @[Switch.scala 41:52:@31984.4]
  wire  output_44_19; // @[Switch.scala 41:38:@31985.4]
  wire  _T_70828; // @[Switch.scala 41:52:@31987.4]
  wire  output_44_20; // @[Switch.scala 41:38:@31988.4]
  wire  _T_70831; // @[Switch.scala 41:52:@31990.4]
  wire  output_44_21; // @[Switch.scala 41:38:@31991.4]
  wire  _T_70834; // @[Switch.scala 41:52:@31993.4]
  wire  output_44_22; // @[Switch.scala 41:38:@31994.4]
  wire  _T_70837; // @[Switch.scala 41:52:@31996.4]
  wire  output_44_23; // @[Switch.scala 41:38:@31997.4]
  wire  _T_70840; // @[Switch.scala 41:52:@31999.4]
  wire  output_44_24; // @[Switch.scala 41:38:@32000.4]
  wire  _T_70843; // @[Switch.scala 41:52:@32002.4]
  wire  output_44_25; // @[Switch.scala 41:38:@32003.4]
  wire  _T_70846; // @[Switch.scala 41:52:@32005.4]
  wire  output_44_26; // @[Switch.scala 41:38:@32006.4]
  wire  _T_70849; // @[Switch.scala 41:52:@32008.4]
  wire  output_44_27; // @[Switch.scala 41:38:@32009.4]
  wire  _T_70852; // @[Switch.scala 41:52:@32011.4]
  wire  output_44_28; // @[Switch.scala 41:38:@32012.4]
  wire  _T_70855; // @[Switch.scala 41:52:@32014.4]
  wire  output_44_29; // @[Switch.scala 41:38:@32015.4]
  wire  _T_70858; // @[Switch.scala 41:52:@32017.4]
  wire  output_44_30; // @[Switch.scala 41:38:@32018.4]
  wire  _T_70861; // @[Switch.scala 41:52:@32020.4]
  wire  output_44_31; // @[Switch.scala 41:38:@32021.4]
  wire  _T_70864; // @[Switch.scala 41:52:@32023.4]
  wire  output_44_32; // @[Switch.scala 41:38:@32024.4]
  wire  _T_70867; // @[Switch.scala 41:52:@32026.4]
  wire  output_44_33; // @[Switch.scala 41:38:@32027.4]
  wire  _T_70870; // @[Switch.scala 41:52:@32029.4]
  wire  output_44_34; // @[Switch.scala 41:38:@32030.4]
  wire  _T_70873; // @[Switch.scala 41:52:@32032.4]
  wire  output_44_35; // @[Switch.scala 41:38:@32033.4]
  wire  _T_70876; // @[Switch.scala 41:52:@32035.4]
  wire  output_44_36; // @[Switch.scala 41:38:@32036.4]
  wire  _T_70879; // @[Switch.scala 41:52:@32038.4]
  wire  output_44_37; // @[Switch.scala 41:38:@32039.4]
  wire  _T_70882; // @[Switch.scala 41:52:@32041.4]
  wire  output_44_38; // @[Switch.scala 41:38:@32042.4]
  wire  _T_70885; // @[Switch.scala 41:52:@32044.4]
  wire  output_44_39; // @[Switch.scala 41:38:@32045.4]
  wire  _T_70888; // @[Switch.scala 41:52:@32047.4]
  wire  output_44_40; // @[Switch.scala 41:38:@32048.4]
  wire  _T_70891; // @[Switch.scala 41:52:@32050.4]
  wire  output_44_41; // @[Switch.scala 41:38:@32051.4]
  wire  _T_70894; // @[Switch.scala 41:52:@32053.4]
  wire  output_44_42; // @[Switch.scala 41:38:@32054.4]
  wire  _T_70897; // @[Switch.scala 41:52:@32056.4]
  wire  output_44_43; // @[Switch.scala 41:38:@32057.4]
  wire  _T_70900; // @[Switch.scala 41:52:@32059.4]
  wire  output_44_44; // @[Switch.scala 41:38:@32060.4]
  wire  _T_70903; // @[Switch.scala 41:52:@32062.4]
  wire  output_44_45; // @[Switch.scala 41:38:@32063.4]
  wire  _T_70906; // @[Switch.scala 41:52:@32065.4]
  wire  output_44_46; // @[Switch.scala 41:38:@32066.4]
  wire  _T_70909; // @[Switch.scala 41:52:@32068.4]
  wire  output_44_47; // @[Switch.scala 41:38:@32069.4]
  wire  _T_70912; // @[Switch.scala 41:52:@32071.4]
  wire  output_44_48; // @[Switch.scala 41:38:@32072.4]
  wire  _T_70915; // @[Switch.scala 41:52:@32074.4]
  wire  output_44_49; // @[Switch.scala 41:38:@32075.4]
  wire  _T_70918; // @[Switch.scala 41:52:@32077.4]
  wire  output_44_50; // @[Switch.scala 41:38:@32078.4]
  wire  _T_70921; // @[Switch.scala 41:52:@32080.4]
  wire  output_44_51; // @[Switch.scala 41:38:@32081.4]
  wire  _T_70924; // @[Switch.scala 41:52:@32083.4]
  wire  output_44_52; // @[Switch.scala 41:38:@32084.4]
  wire  _T_70927; // @[Switch.scala 41:52:@32086.4]
  wire  output_44_53; // @[Switch.scala 41:38:@32087.4]
  wire  _T_70930; // @[Switch.scala 41:52:@32089.4]
  wire  output_44_54; // @[Switch.scala 41:38:@32090.4]
  wire  _T_70933; // @[Switch.scala 41:52:@32092.4]
  wire  output_44_55; // @[Switch.scala 41:38:@32093.4]
  wire  _T_70936; // @[Switch.scala 41:52:@32095.4]
  wire  output_44_56; // @[Switch.scala 41:38:@32096.4]
  wire  _T_70939; // @[Switch.scala 41:52:@32098.4]
  wire  output_44_57; // @[Switch.scala 41:38:@32099.4]
  wire  _T_70942; // @[Switch.scala 41:52:@32101.4]
  wire  output_44_58; // @[Switch.scala 41:38:@32102.4]
  wire  _T_70945; // @[Switch.scala 41:52:@32104.4]
  wire  output_44_59; // @[Switch.scala 41:38:@32105.4]
  wire  _T_70948; // @[Switch.scala 41:52:@32107.4]
  wire  output_44_60; // @[Switch.scala 41:38:@32108.4]
  wire  _T_70951; // @[Switch.scala 41:52:@32110.4]
  wire  output_44_61; // @[Switch.scala 41:38:@32111.4]
  wire  _T_70954; // @[Switch.scala 41:52:@32113.4]
  wire  output_44_62; // @[Switch.scala 41:38:@32114.4]
  wire  _T_70957; // @[Switch.scala 41:52:@32116.4]
  wire  output_44_63; // @[Switch.scala 41:38:@32117.4]
  wire [7:0] _T_70965; // @[Switch.scala 43:31:@32125.4]
  wire [15:0] _T_70973; // @[Switch.scala 43:31:@32133.4]
  wire [7:0] _T_70980; // @[Switch.scala 43:31:@32140.4]
  wire [31:0] _T_70989; // @[Switch.scala 43:31:@32149.4]
  wire [7:0] _T_70996; // @[Switch.scala 43:31:@32156.4]
  wire [15:0] _T_71004; // @[Switch.scala 43:31:@32164.4]
  wire [7:0] _T_71011; // @[Switch.scala 43:31:@32171.4]
  wire [31:0] _T_71020; // @[Switch.scala 43:31:@32180.4]
  wire [63:0] _T_71021; // @[Switch.scala 43:31:@32181.4]
  wire  _T_71025; // @[Switch.scala 41:52:@32184.4]
  wire  output_45_0; // @[Switch.scala 41:38:@32185.4]
  wire  _T_71028; // @[Switch.scala 41:52:@32187.4]
  wire  output_45_1; // @[Switch.scala 41:38:@32188.4]
  wire  _T_71031; // @[Switch.scala 41:52:@32190.4]
  wire  output_45_2; // @[Switch.scala 41:38:@32191.4]
  wire  _T_71034; // @[Switch.scala 41:52:@32193.4]
  wire  output_45_3; // @[Switch.scala 41:38:@32194.4]
  wire  _T_71037; // @[Switch.scala 41:52:@32196.4]
  wire  output_45_4; // @[Switch.scala 41:38:@32197.4]
  wire  _T_71040; // @[Switch.scala 41:52:@32199.4]
  wire  output_45_5; // @[Switch.scala 41:38:@32200.4]
  wire  _T_71043; // @[Switch.scala 41:52:@32202.4]
  wire  output_45_6; // @[Switch.scala 41:38:@32203.4]
  wire  _T_71046; // @[Switch.scala 41:52:@32205.4]
  wire  output_45_7; // @[Switch.scala 41:38:@32206.4]
  wire  _T_71049; // @[Switch.scala 41:52:@32208.4]
  wire  output_45_8; // @[Switch.scala 41:38:@32209.4]
  wire  _T_71052; // @[Switch.scala 41:52:@32211.4]
  wire  output_45_9; // @[Switch.scala 41:38:@32212.4]
  wire  _T_71055; // @[Switch.scala 41:52:@32214.4]
  wire  output_45_10; // @[Switch.scala 41:38:@32215.4]
  wire  _T_71058; // @[Switch.scala 41:52:@32217.4]
  wire  output_45_11; // @[Switch.scala 41:38:@32218.4]
  wire  _T_71061; // @[Switch.scala 41:52:@32220.4]
  wire  output_45_12; // @[Switch.scala 41:38:@32221.4]
  wire  _T_71064; // @[Switch.scala 41:52:@32223.4]
  wire  output_45_13; // @[Switch.scala 41:38:@32224.4]
  wire  _T_71067; // @[Switch.scala 41:52:@32226.4]
  wire  output_45_14; // @[Switch.scala 41:38:@32227.4]
  wire  _T_71070; // @[Switch.scala 41:52:@32229.4]
  wire  output_45_15; // @[Switch.scala 41:38:@32230.4]
  wire  _T_71073; // @[Switch.scala 41:52:@32232.4]
  wire  output_45_16; // @[Switch.scala 41:38:@32233.4]
  wire  _T_71076; // @[Switch.scala 41:52:@32235.4]
  wire  output_45_17; // @[Switch.scala 41:38:@32236.4]
  wire  _T_71079; // @[Switch.scala 41:52:@32238.4]
  wire  output_45_18; // @[Switch.scala 41:38:@32239.4]
  wire  _T_71082; // @[Switch.scala 41:52:@32241.4]
  wire  output_45_19; // @[Switch.scala 41:38:@32242.4]
  wire  _T_71085; // @[Switch.scala 41:52:@32244.4]
  wire  output_45_20; // @[Switch.scala 41:38:@32245.4]
  wire  _T_71088; // @[Switch.scala 41:52:@32247.4]
  wire  output_45_21; // @[Switch.scala 41:38:@32248.4]
  wire  _T_71091; // @[Switch.scala 41:52:@32250.4]
  wire  output_45_22; // @[Switch.scala 41:38:@32251.4]
  wire  _T_71094; // @[Switch.scala 41:52:@32253.4]
  wire  output_45_23; // @[Switch.scala 41:38:@32254.4]
  wire  _T_71097; // @[Switch.scala 41:52:@32256.4]
  wire  output_45_24; // @[Switch.scala 41:38:@32257.4]
  wire  _T_71100; // @[Switch.scala 41:52:@32259.4]
  wire  output_45_25; // @[Switch.scala 41:38:@32260.4]
  wire  _T_71103; // @[Switch.scala 41:52:@32262.4]
  wire  output_45_26; // @[Switch.scala 41:38:@32263.4]
  wire  _T_71106; // @[Switch.scala 41:52:@32265.4]
  wire  output_45_27; // @[Switch.scala 41:38:@32266.4]
  wire  _T_71109; // @[Switch.scala 41:52:@32268.4]
  wire  output_45_28; // @[Switch.scala 41:38:@32269.4]
  wire  _T_71112; // @[Switch.scala 41:52:@32271.4]
  wire  output_45_29; // @[Switch.scala 41:38:@32272.4]
  wire  _T_71115; // @[Switch.scala 41:52:@32274.4]
  wire  output_45_30; // @[Switch.scala 41:38:@32275.4]
  wire  _T_71118; // @[Switch.scala 41:52:@32277.4]
  wire  output_45_31; // @[Switch.scala 41:38:@32278.4]
  wire  _T_71121; // @[Switch.scala 41:52:@32280.4]
  wire  output_45_32; // @[Switch.scala 41:38:@32281.4]
  wire  _T_71124; // @[Switch.scala 41:52:@32283.4]
  wire  output_45_33; // @[Switch.scala 41:38:@32284.4]
  wire  _T_71127; // @[Switch.scala 41:52:@32286.4]
  wire  output_45_34; // @[Switch.scala 41:38:@32287.4]
  wire  _T_71130; // @[Switch.scala 41:52:@32289.4]
  wire  output_45_35; // @[Switch.scala 41:38:@32290.4]
  wire  _T_71133; // @[Switch.scala 41:52:@32292.4]
  wire  output_45_36; // @[Switch.scala 41:38:@32293.4]
  wire  _T_71136; // @[Switch.scala 41:52:@32295.4]
  wire  output_45_37; // @[Switch.scala 41:38:@32296.4]
  wire  _T_71139; // @[Switch.scala 41:52:@32298.4]
  wire  output_45_38; // @[Switch.scala 41:38:@32299.4]
  wire  _T_71142; // @[Switch.scala 41:52:@32301.4]
  wire  output_45_39; // @[Switch.scala 41:38:@32302.4]
  wire  _T_71145; // @[Switch.scala 41:52:@32304.4]
  wire  output_45_40; // @[Switch.scala 41:38:@32305.4]
  wire  _T_71148; // @[Switch.scala 41:52:@32307.4]
  wire  output_45_41; // @[Switch.scala 41:38:@32308.4]
  wire  _T_71151; // @[Switch.scala 41:52:@32310.4]
  wire  output_45_42; // @[Switch.scala 41:38:@32311.4]
  wire  _T_71154; // @[Switch.scala 41:52:@32313.4]
  wire  output_45_43; // @[Switch.scala 41:38:@32314.4]
  wire  _T_71157; // @[Switch.scala 41:52:@32316.4]
  wire  output_45_44; // @[Switch.scala 41:38:@32317.4]
  wire  _T_71160; // @[Switch.scala 41:52:@32319.4]
  wire  output_45_45; // @[Switch.scala 41:38:@32320.4]
  wire  _T_71163; // @[Switch.scala 41:52:@32322.4]
  wire  output_45_46; // @[Switch.scala 41:38:@32323.4]
  wire  _T_71166; // @[Switch.scala 41:52:@32325.4]
  wire  output_45_47; // @[Switch.scala 41:38:@32326.4]
  wire  _T_71169; // @[Switch.scala 41:52:@32328.4]
  wire  output_45_48; // @[Switch.scala 41:38:@32329.4]
  wire  _T_71172; // @[Switch.scala 41:52:@32331.4]
  wire  output_45_49; // @[Switch.scala 41:38:@32332.4]
  wire  _T_71175; // @[Switch.scala 41:52:@32334.4]
  wire  output_45_50; // @[Switch.scala 41:38:@32335.4]
  wire  _T_71178; // @[Switch.scala 41:52:@32337.4]
  wire  output_45_51; // @[Switch.scala 41:38:@32338.4]
  wire  _T_71181; // @[Switch.scala 41:52:@32340.4]
  wire  output_45_52; // @[Switch.scala 41:38:@32341.4]
  wire  _T_71184; // @[Switch.scala 41:52:@32343.4]
  wire  output_45_53; // @[Switch.scala 41:38:@32344.4]
  wire  _T_71187; // @[Switch.scala 41:52:@32346.4]
  wire  output_45_54; // @[Switch.scala 41:38:@32347.4]
  wire  _T_71190; // @[Switch.scala 41:52:@32349.4]
  wire  output_45_55; // @[Switch.scala 41:38:@32350.4]
  wire  _T_71193; // @[Switch.scala 41:52:@32352.4]
  wire  output_45_56; // @[Switch.scala 41:38:@32353.4]
  wire  _T_71196; // @[Switch.scala 41:52:@32355.4]
  wire  output_45_57; // @[Switch.scala 41:38:@32356.4]
  wire  _T_71199; // @[Switch.scala 41:52:@32358.4]
  wire  output_45_58; // @[Switch.scala 41:38:@32359.4]
  wire  _T_71202; // @[Switch.scala 41:52:@32361.4]
  wire  output_45_59; // @[Switch.scala 41:38:@32362.4]
  wire  _T_71205; // @[Switch.scala 41:52:@32364.4]
  wire  output_45_60; // @[Switch.scala 41:38:@32365.4]
  wire  _T_71208; // @[Switch.scala 41:52:@32367.4]
  wire  output_45_61; // @[Switch.scala 41:38:@32368.4]
  wire  _T_71211; // @[Switch.scala 41:52:@32370.4]
  wire  output_45_62; // @[Switch.scala 41:38:@32371.4]
  wire  _T_71214; // @[Switch.scala 41:52:@32373.4]
  wire  output_45_63; // @[Switch.scala 41:38:@32374.4]
  wire [7:0] _T_71222; // @[Switch.scala 43:31:@32382.4]
  wire [15:0] _T_71230; // @[Switch.scala 43:31:@32390.4]
  wire [7:0] _T_71237; // @[Switch.scala 43:31:@32397.4]
  wire [31:0] _T_71246; // @[Switch.scala 43:31:@32406.4]
  wire [7:0] _T_71253; // @[Switch.scala 43:31:@32413.4]
  wire [15:0] _T_71261; // @[Switch.scala 43:31:@32421.4]
  wire [7:0] _T_71268; // @[Switch.scala 43:31:@32428.4]
  wire [31:0] _T_71277; // @[Switch.scala 43:31:@32437.4]
  wire [63:0] _T_71278; // @[Switch.scala 43:31:@32438.4]
  wire  _T_71282; // @[Switch.scala 41:52:@32441.4]
  wire  output_46_0; // @[Switch.scala 41:38:@32442.4]
  wire  _T_71285; // @[Switch.scala 41:52:@32444.4]
  wire  output_46_1; // @[Switch.scala 41:38:@32445.4]
  wire  _T_71288; // @[Switch.scala 41:52:@32447.4]
  wire  output_46_2; // @[Switch.scala 41:38:@32448.4]
  wire  _T_71291; // @[Switch.scala 41:52:@32450.4]
  wire  output_46_3; // @[Switch.scala 41:38:@32451.4]
  wire  _T_71294; // @[Switch.scala 41:52:@32453.4]
  wire  output_46_4; // @[Switch.scala 41:38:@32454.4]
  wire  _T_71297; // @[Switch.scala 41:52:@32456.4]
  wire  output_46_5; // @[Switch.scala 41:38:@32457.4]
  wire  _T_71300; // @[Switch.scala 41:52:@32459.4]
  wire  output_46_6; // @[Switch.scala 41:38:@32460.4]
  wire  _T_71303; // @[Switch.scala 41:52:@32462.4]
  wire  output_46_7; // @[Switch.scala 41:38:@32463.4]
  wire  _T_71306; // @[Switch.scala 41:52:@32465.4]
  wire  output_46_8; // @[Switch.scala 41:38:@32466.4]
  wire  _T_71309; // @[Switch.scala 41:52:@32468.4]
  wire  output_46_9; // @[Switch.scala 41:38:@32469.4]
  wire  _T_71312; // @[Switch.scala 41:52:@32471.4]
  wire  output_46_10; // @[Switch.scala 41:38:@32472.4]
  wire  _T_71315; // @[Switch.scala 41:52:@32474.4]
  wire  output_46_11; // @[Switch.scala 41:38:@32475.4]
  wire  _T_71318; // @[Switch.scala 41:52:@32477.4]
  wire  output_46_12; // @[Switch.scala 41:38:@32478.4]
  wire  _T_71321; // @[Switch.scala 41:52:@32480.4]
  wire  output_46_13; // @[Switch.scala 41:38:@32481.4]
  wire  _T_71324; // @[Switch.scala 41:52:@32483.4]
  wire  output_46_14; // @[Switch.scala 41:38:@32484.4]
  wire  _T_71327; // @[Switch.scala 41:52:@32486.4]
  wire  output_46_15; // @[Switch.scala 41:38:@32487.4]
  wire  _T_71330; // @[Switch.scala 41:52:@32489.4]
  wire  output_46_16; // @[Switch.scala 41:38:@32490.4]
  wire  _T_71333; // @[Switch.scala 41:52:@32492.4]
  wire  output_46_17; // @[Switch.scala 41:38:@32493.4]
  wire  _T_71336; // @[Switch.scala 41:52:@32495.4]
  wire  output_46_18; // @[Switch.scala 41:38:@32496.4]
  wire  _T_71339; // @[Switch.scala 41:52:@32498.4]
  wire  output_46_19; // @[Switch.scala 41:38:@32499.4]
  wire  _T_71342; // @[Switch.scala 41:52:@32501.4]
  wire  output_46_20; // @[Switch.scala 41:38:@32502.4]
  wire  _T_71345; // @[Switch.scala 41:52:@32504.4]
  wire  output_46_21; // @[Switch.scala 41:38:@32505.4]
  wire  _T_71348; // @[Switch.scala 41:52:@32507.4]
  wire  output_46_22; // @[Switch.scala 41:38:@32508.4]
  wire  _T_71351; // @[Switch.scala 41:52:@32510.4]
  wire  output_46_23; // @[Switch.scala 41:38:@32511.4]
  wire  _T_71354; // @[Switch.scala 41:52:@32513.4]
  wire  output_46_24; // @[Switch.scala 41:38:@32514.4]
  wire  _T_71357; // @[Switch.scala 41:52:@32516.4]
  wire  output_46_25; // @[Switch.scala 41:38:@32517.4]
  wire  _T_71360; // @[Switch.scala 41:52:@32519.4]
  wire  output_46_26; // @[Switch.scala 41:38:@32520.4]
  wire  _T_71363; // @[Switch.scala 41:52:@32522.4]
  wire  output_46_27; // @[Switch.scala 41:38:@32523.4]
  wire  _T_71366; // @[Switch.scala 41:52:@32525.4]
  wire  output_46_28; // @[Switch.scala 41:38:@32526.4]
  wire  _T_71369; // @[Switch.scala 41:52:@32528.4]
  wire  output_46_29; // @[Switch.scala 41:38:@32529.4]
  wire  _T_71372; // @[Switch.scala 41:52:@32531.4]
  wire  output_46_30; // @[Switch.scala 41:38:@32532.4]
  wire  _T_71375; // @[Switch.scala 41:52:@32534.4]
  wire  output_46_31; // @[Switch.scala 41:38:@32535.4]
  wire  _T_71378; // @[Switch.scala 41:52:@32537.4]
  wire  output_46_32; // @[Switch.scala 41:38:@32538.4]
  wire  _T_71381; // @[Switch.scala 41:52:@32540.4]
  wire  output_46_33; // @[Switch.scala 41:38:@32541.4]
  wire  _T_71384; // @[Switch.scala 41:52:@32543.4]
  wire  output_46_34; // @[Switch.scala 41:38:@32544.4]
  wire  _T_71387; // @[Switch.scala 41:52:@32546.4]
  wire  output_46_35; // @[Switch.scala 41:38:@32547.4]
  wire  _T_71390; // @[Switch.scala 41:52:@32549.4]
  wire  output_46_36; // @[Switch.scala 41:38:@32550.4]
  wire  _T_71393; // @[Switch.scala 41:52:@32552.4]
  wire  output_46_37; // @[Switch.scala 41:38:@32553.4]
  wire  _T_71396; // @[Switch.scala 41:52:@32555.4]
  wire  output_46_38; // @[Switch.scala 41:38:@32556.4]
  wire  _T_71399; // @[Switch.scala 41:52:@32558.4]
  wire  output_46_39; // @[Switch.scala 41:38:@32559.4]
  wire  _T_71402; // @[Switch.scala 41:52:@32561.4]
  wire  output_46_40; // @[Switch.scala 41:38:@32562.4]
  wire  _T_71405; // @[Switch.scala 41:52:@32564.4]
  wire  output_46_41; // @[Switch.scala 41:38:@32565.4]
  wire  _T_71408; // @[Switch.scala 41:52:@32567.4]
  wire  output_46_42; // @[Switch.scala 41:38:@32568.4]
  wire  _T_71411; // @[Switch.scala 41:52:@32570.4]
  wire  output_46_43; // @[Switch.scala 41:38:@32571.4]
  wire  _T_71414; // @[Switch.scala 41:52:@32573.4]
  wire  output_46_44; // @[Switch.scala 41:38:@32574.4]
  wire  _T_71417; // @[Switch.scala 41:52:@32576.4]
  wire  output_46_45; // @[Switch.scala 41:38:@32577.4]
  wire  _T_71420; // @[Switch.scala 41:52:@32579.4]
  wire  output_46_46; // @[Switch.scala 41:38:@32580.4]
  wire  _T_71423; // @[Switch.scala 41:52:@32582.4]
  wire  output_46_47; // @[Switch.scala 41:38:@32583.4]
  wire  _T_71426; // @[Switch.scala 41:52:@32585.4]
  wire  output_46_48; // @[Switch.scala 41:38:@32586.4]
  wire  _T_71429; // @[Switch.scala 41:52:@32588.4]
  wire  output_46_49; // @[Switch.scala 41:38:@32589.4]
  wire  _T_71432; // @[Switch.scala 41:52:@32591.4]
  wire  output_46_50; // @[Switch.scala 41:38:@32592.4]
  wire  _T_71435; // @[Switch.scala 41:52:@32594.4]
  wire  output_46_51; // @[Switch.scala 41:38:@32595.4]
  wire  _T_71438; // @[Switch.scala 41:52:@32597.4]
  wire  output_46_52; // @[Switch.scala 41:38:@32598.4]
  wire  _T_71441; // @[Switch.scala 41:52:@32600.4]
  wire  output_46_53; // @[Switch.scala 41:38:@32601.4]
  wire  _T_71444; // @[Switch.scala 41:52:@32603.4]
  wire  output_46_54; // @[Switch.scala 41:38:@32604.4]
  wire  _T_71447; // @[Switch.scala 41:52:@32606.4]
  wire  output_46_55; // @[Switch.scala 41:38:@32607.4]
  wire  _T_71450; // @[Switch.scala 41:52:@32609.4]
  wire  output_46_56; // @[Switch.scala 41:38:@32610.4]
  wire  _T_71453; // @[Switch.scala 41:52:@32612.4]
  wire  output_46_57; // @[Switch.scala 41:38:@32613.4]
  wire  _T_71456; // @[Switch.scala 41:52:@32615.4]
  wire  output_46_58; // @[Switch.scala 41:38:@32616.4]
  wire  _T_71459; // @[Switch.scala 41:52:@32618.4]
  wire  output_46_59; // @[Switch.scala 41:38:@32619.4]
  wire  _T_71462; // @[Switch.scala 41:52:@32621.4]
  wire  output_46_60; // @[Switch.scala 41:38:@32622.4]
  wire  _T_71465; // @[Switch.scala 41:52:@32624.4]
  wire  output_46_61; // @[Switch.scala 41:38:@32625.4]
  wire  _T_71468; // @[Switch.scala 41:52:@32627.4]
  wire  output_46_62; // @[Switch.scala 41:38:@32628.4]
  wire  _T_71471; // @[Switch.scala 41:52:@32630.4]
  wire  output_46_63; // @[Switch.scala 41:38:@32631.4]
  wire [7:0] _T_71479; // @[Switch.scala 43:31:@32639.4]
  wire [15:0] _T_71487; // @[Switch.scala 43:31:@32647.4]
  wire [7:0] _T_71494; // @[Switch.scala 43:31:@32654.4]
  wire [31:0] _T_71503; // @[Switch.scala 43:31:@32663.4]
  wire [7:0] _T_71510; // @[Switch.scala 43:31:@32670.4]
  wire [15:0] _T_71518; // @[Switch.scala 43:31:@32678.4]
  wire [7:0] _T_71525; // @[Switch.scala 43:31:@32685.4]
  wire [31:0] _T_71534; // @[Switch.scala 43:31:@32694.4]
  wire [63:0] _T_71535; // @[Switch.scala 43:31:@32695.4]
  wire  _T_71539; // @[Switch.scala 41:52:@32698.4]
  wire  output_47_0; // @[Switch.scala 41:38:@32699.4]
  wire  _T_71542; // @[Switch.scala 41:52:@32701.4]
  wire  output_47_1; // @[Switch.scala 41:38:@32702.4]
  wire  _T_71545; // @[Switch.scala 41:52:@32704.4]
  wire  output_47_2; // @[Switch.scala 41:38:@32705.4]
  wire  _T_71548; // @[Switch.scala 41:52:@32707.4]
  wire  output_47_3; // @[Switch.scala 41:38:@32708.4]
  wire  _T_71551; // @[Switch.scala 41:52:@32710.4]
  wire  output_47_4; // @[Switch.scala 41:38:@32711.4]
  wire  _T_71554; // @[Switch.scala 41:52:@32713.4]
  wire  output_47_5; // @[Switch.scala 41:38:@32714.4]
  wire  _T_71557; // @[Switch.scala 41:52:@32716.4]
  wire  output_47_6; // @[Switch.scala 41:38:@32717.4]
  wire  _T_71560; // @[Switch.scala 41:52:@32719.4]
  wire  output_47_7; // @[Switch.scala 41:38:@32720.4]
  wire  _T_71563; // @[Switch.scala 41:52:@32722.4]
  wire  output_47_8; // @[Switch.scala 41:38:@32723.4]
  wire  _T_71566; // @[Switch.scala 41:52:@32725.4]
  wire  output_47_9; // @[Switch.scala 41:38:@32726.4]
  wire  _T_71569; // @[Switch.scala 41:52:@32728.4]
  wire  output_47_10; // @[Switch.scala 41:38:@32729.4]
  wire  _T_71572; // @[Switch.scala 41:52:@32731.4]
  wire  output_47_11; // @[Switch.scala 41:38:@32732.4]
  wire  _T_71575; // @[Switch.scala 41:52:@32734.4]
  wire  output_47_12; // @[Switch.scala 41:38:@32735.4]
  wire  _T_71578; // @[Switch.scala 41:52:@32737.4]
  wire  output_47_13; // @[Switch.scala 41:38:@32738.4]
  wire  _T_71581; // @[Switch.scala 41:52:@32740.4]
  wire  output_47_14; // @[Switch.scala 41:38:@32741.4]
  wire  _T_71584; // @[Switch.scala 41:52:@32743.4]
  wire  output_47_15; // @[Switch.scala 41:38:@32744.4]
  wire  _T_71587; // @[Switch.scala 41:52:@32746.4]
  wire  output_47_16; // @[Switch.scala 41:38:@32747.4]
  wire  _T_71590; // @[Switch.scala 41:52:@32749.4]
  wire  output_47_17; // @[Switch.scala 41:38:@32750.4]
  wire  _T_71593; // @[Switch.scala 41:52:@32752.4]
  wire  output_47_18; // @[Switch.scala 41:38:@32753.4]
  wire  _T_71596; // @[Switch.scala 41:52:@32755.4]
  wire  output_47_19; // @[Switch.scala 41:38:@32756.4]
  wire  _T_71599; // @[Switch.scala 41:52:@32758.4]
  wire  output_47_20; // @[Switch.scala 41:38:@32759.4]
  wire  _T_71602; // @[Switch.scala 41:52:@32761.4]
  wire  output_47_21; // @[Switch.scala 41:38:@32762.4]
  wire  _T_71605; // @[Switch.scala 41:52:@32764.4]
  wire  output_47_22; // @[Switch.scala 41:38:@32765.4]
  wire  _T_71608; // @[Switch.scala 41:52:@32767.4]
  wire  output_47_23; // @[Switch.scala 41:38:@32768.4]
  wire  _T_71611; // @[Switch.scala 41:52:@32770.4]
  wire  output_47_24; // @[Switch.scala 41:38:@32771.4]
  wire  _T_71614; // @[Switch.scala 41:52:@32773.4]
  wire  output_47_25; // @[Switch.scala 41:38:@32774.4]
  wire  _T_71617; // @[Switch.scala 41:52:@32776.4]
  wire  output_47_26; // @[Switch.scala 41:38:@32777.4]
  wire  _T_71620; // @[Switch.scala 41:52:@32779.4]
  wire  output_47_27; // @[Switch.scala 41:38:@32780.4]
  wire  _T_71623; // @[Switch.scala 41:52:@32782.4]
  wire  output_47_28; // @[Switch.scala 41:38:@32783.4]
  wire  _T_71626; // @[Switch.scala 41:52:@32785.4]
  wire  output_47_29; // @[Switch.scala 41:38:@32786.4]
  wire  _T_71629; // @[Switch.scala 41:52:@32788.4]
  wire  output_47_30; // @[Switch.scala 41:38:@32789.4]
  wire  _T_71632; // @[Switch.scala 41:52:@32791.4]
  wire  output_47_31; // @[Switch.scala 41:38:@32792.4]
  wire  _T_71635; // @[Switch.scala 41:52:@32794.4]
  wire  output_47_32; // @[Switch.scala 41:38:@32795.4]
  wire  _T_71638; // @[Switch.scala 41:52:@32797.4]
  wire  output_47_33; // @[Switch.scala 41:38:@32798.4]
  wire  _T_71641; // @[Switch.scala 41:52:@32800.4]
  wire  output_47_34; // @[Switch.scala 41:38:@32801.4]
  wire  _T_71644; // @[Switch.scala 41:52:@32803.4]
  wire  output_47_35; // @[Switch.scala 41:38:@32804.4]
  wire  _T_71647; // @[Switch.scala 41:52:@32806.4]
  wire  output_47_36; // @[Switch.scala 41:38:@32807.4]
  wire  _T_71650; // @[Switch.scala 41:52:@32809.4]
  wire  output_47_37; // @[Switch.scala 41:38:@32810.4]
  wire  _T_71653; // @[Switch.scala 41:52:@32812.4]
  wire  output_47_38; // @[Switch.scala 41:38:@32813.4]
  wire  _T_71656; // @[Switch.scala 41:52:@32815.4]
  wire  output_47_39; // @[Switch.scala 41:38:@32816.4]
  wire  _T_71659; // @[Switch.scala 41:52:@32818.4]
  wire  output_47_40; // @[Switch.scala 41:38:@32819.4]
  wire  _T_71662; // @[Switch.scala 41:52:@32821.4]
  wire  output_47_41; // @[Switch.scala 41:38:@32822.4]
  wire  _T_71665; // @[Switch.scala 41:52:@32824.4]
  wire  output_47_42; // @[Switch.scala 41:38:@32825.4]
  wire  _T_71668; // @[Switch.scala 41:52:@32827.4]
  wire  output_47_43; // @[Switch.scala 41:38:@32828.4]
  wire  _T_71671; // @[Switch.scala 41:52:@32830.4]
  wire  output_47_44; // @[Switch.scala 41:38:@32831.4]
  wire  _T_71674; // @[Switch.scala 41:52:@32833.4]
  wire  output_47_45; // @[Switch.scala 41:38:@32834.4]
  wire  _T_71677; // @[Switch.scala 41:52:@32836.4]
  wire  output_47_46; // @[Switch.scala 41:38:@32837.4]
  wire  _T_71680; // @[Switch.scala 41:52:@32839.4]
  wire  output_47_47; // @[Switch.scala 41:38:@32840.4]
  wire  _T_71683; // @[Switch.scala 41:52:@32842.4]
  wire  output_47_48; // @[Switch.scala 41:38:@32843.4]
  wire  _T_71686; // @[Switch.scala 41:52:@32845.4]
  wire  output_47_49; // @[Switch.scala 41:38:@32846.4]
  wire  _T_71689; // @[Switch.scala 41:52:@32848.4]
  wire  output_47_50; // @[Switch.scala 41:38:@32849.4]
  wire  _T_71692; // @[Switch.scala 41:52:@32851.4]
  wire  output_47_51; // @[Switch.scala 41:38:@32852.4]
  wire  _T_71695; // @[Switch.scala 41:52:@32854.4]
  wire  output_47_52; // @[Switch.scala 41:38:@32855.4]
  wire  _T_71698; // @[Switch.scala 41:52:@32857.4]
  wire  output_47_53; // @[Switch.scala 41:38:@32858.4]
  wire  _T_71701; // @[Switch.scala 41:52:@32860.4]
  wire  output_47_54; // @[Switch.scala 41:38:@32861.4]
  wire  _T_71704; // @[Switch.scala 41:52:@32863.4]
  wire  output_47_55; // @[Switch.scala 41:38:@32864.4]
  wire  _T_71707; // @[Switch.scala 41:52:@32866.4]
  wire  output_47_56; // @[Switch.scala 41:38:@32867.4]
  wire  _T_71710; // @[Switch.scala 41:52:@32869.4]
  wire  output_47_57; // @[Switch.scala 41:38:@32870.4]
  wire  _T_71713; // @[Switch.scala 41:52:@32872.4]
  wire  output_47_58; // @[Switch.scala 41:38:@32873.4]
  wire  _T_71716; // @[Switch.scala 41:52:@32875.4]
  wire  output_47_59; // @[Switch.scala 41:38:@32876.4]
  wire  _T_71719; // @[Switch.scala 41:52:@32878.4]
  wire  output_47_60; // @[Switch.scala 41:38:@32879.4]
  wire  _T_71722; // @[Switch.scala 41:52:@32881.4]
  wire  output_47_61; // @[Switch.scala 41:38:@32882.4]
  wire  _T_71725; // @[Switch.scala 41:52:@32884.4]
  wire  output_47_62; // @[Switch.scala 41:38:@32885.4]
  wire  _T_71728; // @[Switch.scala 41:52:@32887.4]
  wire  output_47_63; // @[Switch.scala 41:38:@32888.4]
  wire [7:0] _T_71736; // @[Switch.scala 43:31:@32896.4]
  wire [15:0] _T_71744; // @[Switch.scala 43:31:@32904.4]
  wire [7:0] _T_71751; // @[Switch.scala 43:31:@32911.4]
  wire [31:0] _T_71760; // @[Switch.scala 43:31:@32920.4]
  wire [7:0] _T_71767; // @[Switch.scala 43:31:@32927.4]
  wire [15:0] _T_71775; // @[Switch.scala 43:31:@32935.4]
  wire [7:0] _T_71782; // @[Switch.scala 43:31:@32942.4]
  wire [31:0] _T_71791; // @[Switch.scala 43:31:@32951.4]
  wire [63:0] _T_71792; // @[Switch.scala 43:31:@32952.4]
  wire  _T_71796; // @[Switch.scala 41:52:@32955.4]
  wire  output_48_0; // @[Switch.scala 41:38:@32956.4]
  wire  _T_71799; // @[Switch.scala 41:52:@32958.4]
  wire  output_48_1; // @[Switch.scala 41:38:@32959.4]
  wire  _T_71802; // @[Switch.scala 41:52:@32961.4]
  wire  output_48_2; // @[Switch.scala 41:38:@32962.4]
  wire  _T_71805; // @[Switch.scala 41:52:@32964.4]
  wire  output_48_3; // @[Switch.scala 41:38:@32965.4]
  wire  _T_71808; // @[Switch.scala 41:52:@32967.4]
  wire  output_48_4; // @[Switch.scala 41:38:@32968.4]
  wire  _T_71811; // @[Switch.scala 41:52:@32970.4]
  wire  output_48_5; // @[Switch.scala 41:38:@32971.4]
  wire  _T_71814; // @[Switch.scala 41:52:@32973.4]
  wire  output_48_6; // @[Switch.scala 41:38:@32974.4]
  wire  _T_71817; // @[Switch.scala 41:52:@32976.4]
  wire  output_48_7; // @[Switch.scala 41:38:@32977.4]
  wire  _T_71820; // @[Switch.scala 41:52:@32979.4]
  wire  output_48_8; // @[Switch.scala 41:38:@32980.4]
  wire  _T_71823; // @[Switch.scala 41:52:@32982.4]
  wire  output_48_9; // @[Switch.scala 41:38:@32983.4]
  wire  _T_71826; // @[Switch.scala 41:52:@32985.4]
  wire  output_48_10; // @[Switch.scala 41:38:@32986.4]
  wire  _T_71829; // @[Switch.scala 41:52:@32988.4]
  wire  output_48_11; // @[Switch.scala 41:38:@32989.4]
  wire  _T_71832; // @[Switch.scala 41:52:@32991.4]
  wire  output_48_12; // @[Switch.scala 41:38:@32992.4]
  wire  _T_71835; // @[Switch.scala 41:52:@32994.4]
  wire  output_48_13; // @[Switch.scala 41:38:@32995.4]
  wire  _T_71838; // @[Switch.scala 41:52:@32997.4]
  wire  output_48_14; // @[Switch.scala 41:38:@32998.4]
  wire  _T_71841; // @[Switch.scala 41:52:@33000.4]
  wire  output_48_15; // @[Switch.scala 41:38:@33001.4]
  wire  _T_71844; // @[Switch.scala 41:52:@33003.4]
  wire  output_48_16; // @[Switch.scala 41:38:@33004.4]
  wire  _T_71847; // @[Switch.scala 41:52:@33006.4]
  wire  output_48_17; // @[Switch.scala 41:38:@33007.4]
  wire  _T_71850; // @[Switch.scala 41:52:@33009.4]
  wire  output_48_18; // @[Switch.scala 41:38:@33010.4]
  wire  _T_71853; // @[Switch.scala 41:52:@33012.4]
  wire  output_48_19; // @[Switch.scala 41:38:@33013.4]
  wire  _T_71856; // @[Switch.scala 41:52:@33015.4]
  wire  output_48_20; // @[Switch.scala 41:38:@33016.4]
  wire  _T_71859; // @[Switch.scala 41:52:@33018.4]
  wire  output_48_21; // @[Switch.scala 41:38:@33019.4]
  wire  _T_71862; // @[Switch.scala 41:52:@33021.4]
  wire  output_48_22; // @[Switch.scala 41:38:@33022.4]
  wire  _T_71865; // @[Switch.scala 41:52:@33024.4]
  wire  output_48_23; // @[Switch.scala 41:38:@33025.4]
  wire  _T_71868; // @[Switch.scala 41:52:@33027.4]
  wire  output_48_24; // @[Switch.scala 41:38:@33028.4]
  wire  _T_71871; // @[Switch.scala 41:52:@33030.4]
  wire  output_48_25; // @[Switch.scala 41:38:@33031.4]
  wire  _T_71874; // @[Switch.scala 41:52:@33033.4]
  wire  output_48_26; // @[Switch.scala 41:38:@33034.4]
  wire  _T_71877; // @[Switch.scala 41:52:@33036.4]
  wire  output_48_27; // @[Switch.scala 41:38:@33037.4]
  wire  _T_71880; // @[Switch.scala 41:52:@33039.4]
  wire  output_48_28; // @[Switch.scala 41:38:@33040.4]
  wire  _T_71883; // @[Switch.scala 41:52:@33042.4]
  wire  output_48_29; // @[Switch.scala 41:38:@33043.4]
  wire  _T_71886; // @[Switch.scala 41:52:@33045.4]
  wire  output_48_30; // @[Switch.scala 41:38:@33046.4]
  wire  _T_71889; // @[Switch.scala 41:52:@33048.4]
  wire  output_48_31; // @[Switch.scala 41:38:@33049.4]
  wire  _T_71892; // @[Switch.scala 41:52:@33051.4]
  wire  output_48_32; // @[Switch.scala 41:38:@33052.4]
  wire  _T_71895; // @[Switch.scala 41:52:@33054.4]
  wire  output_48_33; // @[Switch.scala 41:38:@33055.4]
  wire  _T_71898; // @[Switch.scala 41:52:@33057.4]
  wire  output_48_34; // @[Switch.scala 41:38:@33058.4]
  wire  _T_71901; // @[Switch.scala 41:52:@33060.4]
  wire  output_48_35; // @[Switch.scala 41:38:@33061.4]
  wire  _T_71904; // @[Switch.scala 41:52:@33063.4]
  wire  output_48_36; // @[Switch.scala 41:38:@33064.4]
  wire  _T_71907; // @[Switch.scala 41:52:@33066.4]
  wire  output_48_37; // @[Switch.scala 41:38:@33067.4]
  wire  _T_71910; // @[Switch.scala 41:52:@33069.4]
  wire  output_48_38; // @[Switch.scala 41:38:@33070.4]
  wire  _T_71913; // @[Switch.scala 41:52:@33072.4]
  wire  output_48_39; // @[Switch.scala 41:38:@33073.4]
  wire  _T_71916; // @[Switch.scala 41:52:@33075.4]
  wire  output_48_40; // @[Switch.scala 41:38:@33076.4]
  wire  _T_71919; // @[Switch.scala 41:52:@33078.4]
  wire  output_48_41; // @[Switch.scala 41:38:@33079.4]
  wire  _T_71922; // @[Switch.scala 41:52:@33081.4]
  wire  output_48_42; // @[Switch.scala 41:38:@33082.4]
  wire  _T_71925; // @[Switch.scala 41:52:@33084.4]
  wire  output_48_43; // @[Switch.scala 41:38:@33085.4]
  wire  _T_71928; // @[Switch.scala 41:52:@33087.4]
  wire  output_48_44; // @[Switch.scala 41:38:@33088.4]
  wire  _T_71931; // @[Switch.scala 41:52:@33090.4]
  wire  output_48_45; // @[Switch.scala 41:38:@33091.4]
  wire  _T_71934; // @[Switch.scala 41:52:@33093.4]
  wire  output_48_46; // @[Switch.scala 41:38:@33094.4]
  wire  _T_71937; // @[Switch.scala 41:52:@33096.4]
  wire  output_48_47; // @[Switch.scala 41:38:@33097.4]
  wire  _T_71940; // @[Switch.scala 41:52:@33099.4]
  wire  output_48_48; // @[Switch.scala 41:38:@33100.4]
  wire  _T_71943; // @[Switch.scala 41:52:@33102.4]
  wire  output_48_49; // @[Switch.scala 41:38:@33103.4]
  wire  _T_71946; // @[Switch.scala 41:52:@33105.4]
  wire  output_48_50; // @[Switch.scala 41:38:@33106.4]
  wire  _T_71949; // @[Switch.scala 41:52:@33108.4]
  wire  output_48_51; // @[Switch.scala 41:38:@33109.4]
  wire  _T_71952; // @[Switch.scala 41:52:@33111.4]
  wire  output_48_52; // @[Switch.scala 41:38:@33112.4]
  wire  _T_71955; // @[Switch.scala 41:52:@33114.4]
  wire  output_48_53; // @[Switch.scala 41:38:@33115.4]
  wire  _T_71958; // @[Switch.scala 41:52:@33117.4]
  wire  output_48_54; // @[Switch.scala 41:38:@33118.4]
  wire  _T_71961; // @[Switch.scala 41:52:@33120.4]
  wire  output_48_55; // @[Switch.scala 41:38:@33121.4]
  wire  _T_71964; // @[Switch.scala 41:52:@33123.4]
  wire  output_48_56; // @[Switch.scala 41:38:@33124.4]
  wire  _T_71967; // @[Switch.scala 41:52:@33126.4]
  wire  output_48_57; // @[Switch.scala 41:38:@33127.4]
  wire  _T_71970; // @[Switch.scala 41:52:@33129.4]
  wire  output_48_58; // @[Switch.scala 41:38:@33130.4]
  wire  _T_71973; // @[Switch.scala 41:52:@33132.4]
  wire  output_48_59; // @[Switch.scala 41:38:@33133.4]
  wire  _T_71976; // @[Switch.scala 41:52:@33135.4]
  wire  output_48_60; // @[Switch.scala 41:38:@33136.4]
  wire  _T_71979; // @[Switch.scala 41:52:@33138.4]
  wire  output_48_61; // @[Switch.scala 41:38:@33139.4]
  wire  _T_71982; // @[Switch.scala 41:52:@33141.4]
  wire  output_48_62; // @[Switch.scala 41:38:@33142.4]
  wire  _T_71985; // @[Switch.scala 41:52:@33144.4]
  wire  output_48_63; // @[Switch.scala 41:38:@33145.4]
  wire [7:0] _T_71993; // @[Switch.scala 43:31:@33153.4]
  wire [15:0] _T_72001; // @[Switch.scala 43:31:@33161.4]
  wire [7:0] _T_72008; // @[Switch.scala 43:31:@33168.4]
  wire [31:0] _T_72017; // @[Switch.scala 43:31:@33177.4]
  wire [7:0] _T_72024; // @[Switch.scala 43:31:@33184.4]
  wire [15:0] _T_72032; // @[Switch.scala 43:31:@33192.4]
  wire [7:0] _T_72039; // @[Switch.scala 43:31:@33199.4]
  wire [31:0] _T_72048; // @[Switch.scala 43:31:@33208.4]
  wire [63:0] _T_72049; // @[Switch.scala 43:31:@33209.4]
  wire  _T_72053; // @[Switch.scala 41:52:@33212.4]
  wire  output_49_0; // @[Switch.scala 41:38:@33213.4]
  wire  _T_72056; // @[Switch.scala 41:52:@33215.4]
  wire  output_49_1; // @[Switch.scala 41:38:@33216.4]
  wire  _T_72059; // @[Switch.scala 41:52:@33218.4]
  wire  output_49_2; // @[Switch.scala 41:38:@33219.4]
  wire  _T_72062; // @[Switch.scala 41:52:@33221.4]
  wire  output_49_3; // @[Switch.scala 41:38:@33222.4]
  wire  _T_72065; // @[Switch.scala 41:52:@33224.4]
  wire  output_49_4; // @[Switch.scala 41:38:@33225.4]
  wire  _T_72068; // @[Switch.scala 41:52:@33227.4]
  wire  output_49_5; // @[Switch.scala 41:38:@33228.4]
  wire  _T_72071; // @[Switch.scala 41:52:@33230.4]
  wire  output_49_6; // @[Switch.scala 41:38:@33231.4]
  wire  _T_72074; // @[Switch.scala 41:52:@33233.4]
  wire  output_49_7; // @[Switch.scala 41:38:@33234.4]
  wire  _T_72077; // @[Switch.scala 41:52:@33236.4]
  wire  output_49_8; // @[Switch.scala 41:38:@33237.4]
  wire  _T_72080; // @[Switch.scala 41:52:@33239.4]
  wire  output_49_9; // @[Switch.scala 41:38:@33240.4]
  wire  _T_72083; // @[Switch.scala 41:52:@33242.4]
  wire  output_49_10; // @[Switch.scala 41:38:@33243.4]
  wire  _T_72086; // @[Switch.scala 41:52:@33245.4]
  wire  output_49_11; // @[Switch.scala 41:38:@33246.4]
  wire  _T_72089; // @[Switch.scala 41:52:@33248.4]
  wire  output_49_12; // @[Switch.scala 41:38:@33249.4]
  wire  _T_72092; // @[Switch.scala 41:52:@33251.4]
  wire  output_49_13; // @[Switch.scala 41:38:@33252.4]
  wire  _T_72095; // @[Switch.scala 41:52:@33254.4]
  wire  output_49_14; // @[Switch.scala 41:38:@33255.4]
  wire  _T_72098; // @[Switch.scala 41:52:@33257.4]
  wire  output_49_15; // @[Switch.scala 41:38:@33258.4]
  wire  _T_72101; // @[Switch.scala 41:52:@33260.4]
  wire  output_49_16; // @[Switch.scala 41:38:@33261.4]
  wire  _T_72104; // @[Switch.scala 41:52:@33263.4]
  wire  output_49_17; // @[Switch.scala 41:38:@33264.4]
  wire  _T_72107; // @[Switch.scala 41:52:@33266.4]
  wire  output_49_18; // @[Switch.scala 41:38:@33267.4]
  wire  _T_72110; // @[Switch.scala 41:52:@33269.4]
  wire  output_49_19; // @[Switch.scala 41:38:@33270.4]
  wire  _T_72113; // @[Switch.scala 41:52:@33272.4]
  wire  output_49_20; // @[Switch.scala 41:38:@33273.4]
  wire  _T_72116; // @[Switch.scala 41:52:@33275.4]
  wire  output_49_21; // @[Switch.scala 41:38:@33276.4]
  wire  _T_72119; // @[Switch.scala 41:52:@33278.4]
  wire  output_49_22; // @[Switch.scala 41:38:@33279.4]
  wire  _T_72122; // @[Switch.scala 41:52:@33281.4]
  wire  output_49_23; // @[Switch.scala 41:38:@33282.4]
  wire  _T_72125; // @[Switch.scala 41:52:@33284.4]
  wire  output_49_24; // @[Switch.scala 41:38:@33285.4]
  wire  _T_72128; // @[Switch.scala 41:52:@33287.4]
  wire  output_49_25; // @[Switch.scala 41:38:@33288.4]
  wire  _T_72131; // @[Switch.scala 41:52:@33290.4]
  wire  output_49_26; // @[Switch.scala 41:38:@33291.4]
  wire  _T_72134; // @[Switch.scala 41:52:@33293.4]
  wire  output_49_27; // @[Switch.scala 41:38:@33294.4]
  wire  _T_72137; // @[Switch.scala 41:52:@33296.4]
  wire  output_49_28; // @[Switch.scala 41:38:@33297.4]
  wire  _T_72140; // @[Switch.scala 41:52:@33299.4]
  wire  output_49_29; // @[Switch.scala 41:38:@33300.4]
  wire  _T_72143; // @[Switch.scala 41:52:@33302.4]
  wire  output_49_30; // @[Switch.scala 41:38:@33303.4]
  wire  _T_72146; // @[Switch.scala 41:52:@33305.4]
  wire  output_49_31; // @[Switch.scala 41:38:@33306.4]
  wire  _T_72149; // @[Switch.scala 41:52:@33308.4]
  wire  output_49_32; // @[Switch.scala 41:38:@33309.4]
  wire  _T_72152; // @[Switch.scala 41:52:@33311.4]
  wire  output_49_33; // @[Switch.scala 41:38:@33312.4]
  wire  _T_72155; // @[Switch.scala 41:52:@33314.4]
  wire  output_49_34; // @[Switch.scala 41:38:@33315.4]
  wire  _T_72158; // @[Switch.scala 41:52:@33317.4]
  wire  output_49_35; // @[Switch.scala 41:38:@33318.4]
  wire  _T_72161; // @[Switch.scala 41:52:@33320.4]
  wire  output_49_36; // @[Switch.scala 41:38:@33321.4]
  wire  _T_72164; // @[Switch.scala 41:52:@33323.4]
  wire  output_49_37; // @[Switch.scala 41:38:@33324.4]
  wire  _T_72167; // @[Switch.scala 41:52:@33326.4]
  wire  output_49_38; // @[Switch.scala 41:38:@33327.4]
  wire  _T_72170; // @[Switch.scala 41:52:@33329.4]
  wire  output_49_39; // @[Switch.scala 41:38:@33330.4]
  wire  _T_72173; // @[Switch.scala 41:52:@33332.4]
  wire  output_49_40; // @[Switch.scala 41:38:@33333.4]
  wire  _T_72176; // @[Switch.scala 41:52:@33335.4]
  wire  output_49_41; // @[Switch.scala 41:38:@33336.4]
  wire  _T_72179; // @[Switch.scala 41:52:@33338.4]
  wire  output_49_42; // @[Switch.scala 41:38:@33339.4]
  wire  _T_72182; // @[Switch.scala 41:52:@33341.4]
  wire  output_49_43; // @[Switch.scala 41:38:@33342.4]
  wire  _T_72185; // @[Switch.scala 41:52:@33344.4]
  wire  output_49_44; // @[Switch.scala 41:38:@33345.4]
  wire  _T_72188; // @[Switch.scala 41:52:@33347.4]
  wire  output_49_45; // @[Switch.scala 41:38:@33348.4]
  wire  _T_72191; // @[Switch.scala 41:52:@33350.4]
  wire  output_49_46; // @[Switch.scala 41:38:@33351.4]
  wire  _T_72194; // @[Switch.scala 41:52:@33353.4]
  wire  output_49_47; // @[Switch.scala 41:38:@33354.4]
  wire  _T_72197; // @[Switch.scala 41:52:@33356.4]
  wire  output_49_48; // @[Switch.scala 41:38:@33357.4]
  wire  _T_72200; // @[Switch.scala 41:52:@33359.4]
  wire  output_49_49; // @[Switch.scala 41:38:@33360.4]
  wire  _T_72203; // @[Switch.scala 41:52:@33362.4]
  wire  output_49_50; // @[Switch.scala 41:38:@33363.4]
  wire  _T_72206; // @[Switch.scala 41:52:@33365.4]
  wire  output_49_51; // @[Switch.scala 41:38:@33366.4]
  wire  _T_72209; // @[Switch.scala 41:52:@33368.4]
  wire  output_49_52; // @[Switch.scala 41:38:@33369.4]
  wire  _T_72212; // @[Switch.scala 41:52:@33371.4]
  wire  output_49_53; // @[Switch.scala 41:38:@33372.4]
  wire  _T_72215; // @[Switch.scala 41:52:@33374.4]
  wire  output_49_54; // @[Switch.scala 41:38:@33375.4]
  wire  _T_72218; // @[Switch.scala 41:52:@33377.4]
  wire  output_49_55; // @[Switch.scala 41:38:@33378.4]
  wire  _T_72221; // @[Switch.scala 41:52:@33380.4]
  wire  output_49_56; // @[Switch.scala 41:38:@33381.4]
  wire  _T_72224; // @[Switch.scala 41:52:@33383.4]
  wire  output_49_57; // @[Switch.scala 41:38:@33384.4]
  wire  _T_72227; // @[Switch.scala 41:52:@33386.4]
  wire  output_49_58; // @[Switch.scala 41:38:@33387.4]
  wire  _T_72230; // @[Switch.scala 41:52:@33389.4]
  wire  output_49_59; // @[Switch.scala 41:38:@33390.4]
  wire  _T_72233; // @[Switch.scala 41:52:@33392.4]
  wire  output_49_60; // @[Switch.scala 41:38:@33393.4]
  wire  _T_72236; // @[Switch.scala 41:52:@33395.4]
  wire  output_49_61; // @[Switch.scala 41:38:@33396.4]
  wire  _T_72239; // @[Switch.scala 41:52:@33398.4]
  wire  output_49_62; // @[Switch.scala 41:38:@33399.4]
  wire  _T_72242; // @[Switch.scala 41:52:@33401.4]
  wire  output_49_63; // @[Switch.scala 41:38:@33402.4]
  wire [7:0] _T_72250; // @[Switch.scala 43:31:@33410.4]
  wire [15:0] _T_72258; // @[Switch.scala 43:31:@33418.4]
  wire [7:0] _T_72265; // @[Switch.scala 43:31:@33425.4]
  wire [31:0] _T_72274; // @[Switch.scala 43:31:@33434.4]
  wire [7:0] _T_72281; // @[Switch.scala 43:31:@33441.4]
  wire [15:0] _T_72289; // @[Switch.scala 43:31:@33449.4]
  wire [7:0] _T_72296; // @[Switch.scala 43:31:@33456.4]
  wire [31:0] _T_72305; // @[Switch.scala 43:31:@33465.4]
  wire [63:0] _T_72306; // @[Switch.scala 43:31:@33466.4]
  wire  _T_72310; // @[Switch.scala 41:52:@33469.4]
  wire  output_50_0; // @[Switch.scala 41:38:@33470.4]
  wire  _T_72313; // @[Switch.scala 41:52:@33472.4]
  wire  output_50_1; // @[Switch.scala 41:38:@33473.4]
  wire  _T_72316; // @[Switch.scala 41:52:@33475.4]
  wire  output_50_2; // @[Switch.scala 41:38:@33476.4]
  wire  _T_72319; // @[Switch.scala 41:52:@33478.4]
  wire  output_50_3; // @[Switch.scala 41:38:@33479.4]
  wire  _T_72322; // @[Switch.scala 41:52:@33481.4]
  wire  output_50_4; // @[Switch.scala 41:38:@33482.4]
  wire  _T_72325; // @[Switch.scala 41:52:@33484.4]
  wire  output_50_5; // @[Switch.scala 41:38:@33485.4]
  wire  _T_72328; // @[Switch.scala 41:52:@33487.4]
  wire  output_50_6; // @[Switch.scala 41:38:@33488.4]
  wire  _T_72331; // @[Switch.scala 41:52:@33490.4]
  wire  output_50_7; // @[Switch.scala 41:38:@33491.4]
  wire  _T_72334; // @[Switch.scala 41:52:@33493.4]
  wire  output_50_8; // @[Switch.scala 41:38:@33494.4]
  wire  _T_72337; // @[Switch.scala 41:52:@33496.4]
  wire  output_50_9; // @[Switch.scala 41:38:@33497.4]
  wire  _T_72340; // @[Switch.scala 41:52:@33499.4]
  wire  output_50_10; // @[Switch.scala 41:38:@33500.4]
  wire  _T_72343; // @[Switch.scala 41:52:@33502.4]
  wire  output_50_11; // @[Switch.scala 41:38:@33503.4]
  wire  _T_72346; // @[Switch.scala 41:52:@33505.4]
  wire  output_50_12; // @[Switch.scala 41:38:@33506.4]
  wire  _T_72349; // @[Switch.scala 41:52:@33508.4]
  wire  output_50_13; // @[Switch.scala 41:38:@33509.4]
  wire  _T_72352; // @[Switch.scala 41:52:@33511.4]
  wire  output_50_14; // @[Switch.scala 41:38:@33512.4]
  wire  _T_72355; // @[Switch.scala 41:52:@33514.4]
  wire  output_50_15; // @[Switch.scala 41:38:@33515.4]
  wire  _T_72358; // @[Switch.scala 41:52:@33517.4]
  wire  output_50_16; // @[Switch.scala 41:38:@33518.4]
  wire  _T_72361; // @[Switch.scala 41:52:@33520.4]
  wire  output_50_17; // @[Switch.scala 41:38:@33521.4]
  wire  _T_72364; // @[Switch.scala 41:52:@33523.4]
  wire  output_50_18; // @[Switch.scala 41:38:@33524.4]
  wire  _T_72367; // @[Switch.scala 41:52:@33526.4]
  wire  output_50_19; // @[Switch.scala 41:38:@33527.4]
  wire  _T_72370; // @[Switch.scala 41:52:@33529.4]
  wire  output_50_20; // @[Switch.scala 41:38:@33530.4]
  wire  _T_72373; // @[Switch.scala 41:52:@33532.4]
  wire  output_50_21; // @[Switch.scala 41:38:@33533.4]
  wire  _T_72376; // @[Switch.scala 41:52:@33535.4]
  wire  output_50_22; // @[Switch.scala 41:38:@33536.4]
  wire  _T_72379; // @[Switch.scala 41:52:@33538.4]
  wire  output_50_23; // @[Switch.scala 41:38:@33539.4]
  wire  _T_72382; // @[Switch.scala 41:52:@33541.4]
  wire  output_50_24; // @[Switch.scala 41:38:@33542.4]
  wire  _T_72385; // @[Switch.scala 41:52:@33544.4]
  wire  output_50_25; // @[Switch.scala 41:38:@33545.4]
  wire  _T_72388; // @[Switch.scala 41:52:@33547.4]
  wire  output_50_26; // @[Switch.scala 41:38:@33548.4]
  wire  _T_72391; // @[Switch.scala 41:52:@33550.4]
  wire  output_50_27; // @[Switch.scala 41:38:@33551.4]
  wire  _T_72394; // @[Switch.scala 41:52:@33553.4]
  wire  output_50_28; // @[Switch.scala 41:38:@33554.4]
  wire  _T_72397; // @[Switch.scala 41:52:@33556.4]
  wire  output_50_29; // @[Switch.scala 41:38:@33557.4]
  wire  _T_72400; // @[Switch.scala 41:52:@33559.4]
  wire  output_50_30; // @[Switch.scala 41:38:@33560.4]
  wire  _T_72403; // @[Switch.scala 41:52:@33562.4]
  wire  output_50_31; // @[Switch.scala 41:38:@33563.4]
  wire  _T_72406; // @[Switch.scala 41:52:@33565.4]
  wire  output_50_32; // @[Switch.scala 41:38:@33566.4]
  wire  _T_72409; // @[Switch.scala 41:52:@33568.4]
  wire  output_50_33; // @[Switch.scala 41:38:@33569.4]
  wire  _T_72412; // @[Switch.scala 41:52:@33571.4]
  wire  output_50_34; // @[Switch.scala 41:38:@33572.4]
  wire  _T_72415; // @[Switch.scala 41:52:@33574.4]
  wire  output_50_35; // @[Switch.scala 41:38:@33575.4]
  wire  _T_72418; // @[Switch.scala 41:52:@33577.4]
  wire  output_50_36; // @[Switch.scala 41:38:@33578.4]
  wire  _T_72421; // @[Switch.scala 41:52:@33580.4]
  wire  output_50_37; // @[Switch.scala 41:38:@33581.4]
  wire  _T_72424; // @[Switch.scala 41:52:@33583.4]
  wire  output_50_38; // @[Switch.scala 41:38:@33584.4]
  wire  _T_72427; // @[Switch.scala 41:52:@33586.4]
  wire  output_50_39; // @[Switch.scala 41:38:@33587.4]
  wire  _T_72430; // @[Switch.scala 41:52:@33589.4]
  wire  output_50_40; // @[Switch.scala 41:38:@33590.4]
  wire  _T_72433; // @[Switch.scala 41:52:@33592.4]
  wire  output_50_41; // @[Switch.scala 41:38:@33593.4]
  wire  _T_72436; // @[Switch.scala 41:52:@33595.4]
  wire  output_50_42; // @[Switch.scala 41:38:@33596.4]
  wire  _T_72439; // @[Switch.scala 41:52:@33598.4]
  wire  output_50_43; // @[Switch.scala 41:38:@33599.4]
  wire  _T_72442; // @[Switch.scala 41:52:@33601.4]
  wire  output_50_44; // @[Switch.scala 41:38:@33602.4]
  wire  _T_72445; // @[Switch.scala 41:52:@33604.4]
  wire  output_50_45; // @[Switch.scala 41:38:@33605.4]
  wire  _T_72448; // @[Switch.scala 41:52:@33607.4]
  wire  output_50_46; // @[Switch.scala 41:38:@33608.4]
  wire  _T_72451; // @[Switch.scala 41:52:@33610.4]
  wire  output_50_47; // @[Switch.scala 41:38:@33611.4]
  wire  _T_72454; // @[Switch.scala 41:52:@33613.4]
  wire  output_50_48; // @[Switch.scala 41:38:@33614.4]
  wire  _T_72457; // @[Switch.scala 41:52:@33616.4]
  wire  output_50_49; // @[Switch.scala 41:38:@33617.4]
  wire  _T_72460; // @[Switch.scala 41:52:@33619.4]
  wire  output_50_50; // @[Switch.scala 41:38:@33620.4]
  wire  _T_72463; // @[Switch.scala 41:52:@33622.4]
  wire  output_50_51; // @[Switch.scala 41:38:@33623.4]
  wire  _T_72466; // @[Switch.scala 41:52:@33625.4]
  wire  output_50_52; // @[Switch.scala 41:38:@33626.4]
  wire  _T_72469; // @[Switch.scala 41:52:@33628.4]
  wire  output_50_53; // @[Switch.scala 41:38:@33629.4]
  wire  _T_72472; // @[Switch.scala 41:52:@33631.4]
  wire  output_50_54; // @[Switch.scala 41:38:@33632.4]
  wire  _T_72475; // @[Switch.scala 41:52:@33634.4]
  wire  output_50_55; // @[Switch.scala 41:38:@33635.4]
  wire  _T_72478; // @[Switch.scala 41:52:@33637.4]
  wire  output_50_56; // @[Switch.scala 41:38:@33638.4]
  wire  _T_72481; // @[Switch.scala 41:52:@33640.4]
  wire  output_50_57; // @[Switch.scala 41:38:@33641.4]
  wire  _T_72484; // @[Switch.scala 41:52:@33643.4]
  wire  output_50_58; // @[Switch.scala 41:38:@33644.4]
  wire  _T_72487; // @[Switch.scala 41:52:@33646.4]
  wire  output_50_59; // @[Switch.scala 41:38:@33647.4]
  wire  _T_72490; // @[Switch.scala 41:52:@33649.4]
  wire  output_50_60; // @[Switch.scala 41:38:@33650.4]
  wire  _T_72493; // @[Switch.scala 41:52:@33652.4]
  wire  output_50_61; // @[Switch.scala 41:38:@33653.4]
  wire  _T_72496; // @[Switch.scala 41:52:@33655.4]
  wire  output_50_62; // @[Switch.scala 41:38:@33656.4]
  wire  _T_72499; // @[Switch.scala 41:52:@33658.4]
  wire  output_50_63; // @[Switch.scala 41:38:@33659.4]
  wire [7:0] _T_72507; // @[Switch.scala 43:31:@33667.4]
  wire [15:0] _T_72515; // @[Switch.scala 43:31:@33675.4]
  wire [7:0] _T_72522; // @[Switch.scala 43:31:@33682.4]
  wire [31:0] _T_72531; // @[Switch.scala 43:31:@33691.4]
  wire [7:0] _T_72538; // @[Switch.scala 43:31:@33698.4]
  wire [15:0] _T_72546; // @[Switch.scala 43:31:@33706.4]
  wire [7:0] _T_72553; // @[Switch.scala 43:31:@33713.4]
  wire [31:0] _T_72562; // @[Switch.scala 43:31:@33722.4]
  wire [63:0] _T_72563; // @[Switch.scala 43:31:@33723.4]
  wire  _T_72567; // @[Switch.scala 41:52:@33726.4]
  wire  output_51_0; // @[Switch.scala 41:38:@33727.4]
  wire  _T_72570; // @[Switch.scala 41:52:@33729.4]
  wire  output_51_1; // @[Switch.scala 41:38:@33730.4]
  wire  _T_72573; // @[Switch.scala 41:52:@33732.4]
  wire  output_51_2; // @[Switch.scala 41:38:@33733.4]
  wire  _T_72576; // @[Switch.scala 41:52:@33735.4]
  wire  output_51_3; // @[Switch.scala 41:38:@33736.4]
  wire  _T_72579; // @[Switch.scala 41:52:@33738.4]
  wire  output_51_4; // @[Switch.scala 41:38:@33739.4]
  wire  _T_72582; // @[Switch.scala 41:52:@33741.4]
  wire  output_51_5; // @[Switch.scala 41:38:@33742.4]
  wire  _T_72585; // @[Switch.scala 41:52:@33744.4]
  wire  output_51_6; // @[Switch.scala 41:38:@33745.4]
  wire  _T_72588; // @[Switch.scala 41:52:@33747.4]
  wire  output_51_7; // @[Switch.scala 41:38:@33748.4]
  wire  _T_72591; // @[Switch.scala 41:52:@33750.4]
  wire  output_51_8; // @[Switch.scala 41:38:@33751.4]
  wire  _T_72594; // @[Switch.scala 41:52:@33753.4]
  wire  output_51_9; // @[Switch.scala 41:38:@33754.4]
  wire  _T_72597; // @[Switch.scala 41:52:@33756.4]
  wire  output_51_10; // @[Switch.scala 41:38:@33757.4]
  wire  _T_72600; // @[Switch.scala 41:52:@33759.4]
  wire  output_51_11; // @[Switch.scala 41:38:@33760.4]
  wire  _T_72603; // @[Switch.scala 41:52:@33762.4]
  wire  output_51_12; // @[Switch.scala 41:38:@33763.4]
  wire  _T_72606; // @[Switch.scala 41:52:@33765.4]
  wire  output_51_13; // @[Switch.scala 41:38:@33766.4]
  wire  _T_72609; // @[Switch.scala 41:52:@33768.4]
  wire  output_51_14; // @[Switch.scala 41:38:@33769.4]
  wire  _T_72612; // @[Switch.scala 41:52:@33771.4]
  wire  output_51_15; // @[Switch.scala 41:38:@33772.4]
  wire  _T_72615; // @[Switch.scala 41:52:@33774.4]
  wire  output_51_16; // @[Switch.scala 41:38:@33775.4]
  wire  _T_72618; // @[Switch.scala 41:52:@33777.4]
  wire  output_51_17; // @[Switch.scala 41:38:@33778.4]
  wire  _T_72621; // @[Switch.scala 41:52:@33780.4]
  wire  output_51_18; // @[Switch.scala 41:38:@33781.4]
  wire  _T_72624; // @[Switch.scala 41:52:@33783.4]
  wire  output_51_19; // @[Switch.scala 41:38:@33784.4]
  wire  _T_72627; // @[Switch.scala 41:52:@33786.4]
  wire  output_51_20; // @[Switch.scala 41:38:@33787.4]
  wire  _T_72630; // @[Switch.scala 41:52:@33789.4]
  wire  output_51_21; // @[Switch.scala 41:38:@33790.4]
  wire  _T_72633; // @[Switch.scala 41:52:@33792.4]
  wire  output_51_22; // @[Switch.scala 41:38:@33793.4]
  wire  _T_72636; // @[Switch.scala 41:52:@33795.4]
  wire  output_51_23; // @[Switch.scala 41:38:@33796.4]
  wire  _T_72639; // @[Switch.scala 41:52:@33798.4]
  wire  output_51_24; // @[Switch.scala 41:38:@33799.4]
  wire  _T_72642; // @[Switch.scala 41:52:@33801.4]
  wire  output_51_25; // @[Switch.scala 41:38:@33802.4]
  wire  _T_72645; // @[Switch.scala 41:52:@33804.4]
  wire  output_51_26; // @[Switch.scala 41:38:@33805.4]
  wire  _T_72648; // @[Switch.scala 41:52:@33807.4]
  wire  output_51_27; // @[Switch.scala 41:38:@33808.4]
  wire  _T_72651; // @[Switch.scala 41:52:@33810.4]
  wire  output_51_28; // @[Switch.scala 41:38:@33811.4]
  wire  _T_72654; // @[Switch.scala 41:52:@33813.4]
  wire  output_51_29; // @[Switch.scala 41:38:@33814.4]
  wire  _T_72657; // @[Switch.scala 41:52:@33816.4]
  wire  output_51_30; // @[Switch.scala 41:38:@33817.4]
  wire  _T_72660; // @[Switch.scala 41:52:@33819.4]
  wire  output_51_31; // @[Switch.scala 41:38:@33820.4]
  wire  _T_72663; // @[Switch.scala 41:52:@33822.4]
  wire  output_51_32; // @[Switch.scala 41:38:@33823.4]
  wire  _T_72666; // @[Switch.scala 41:52:@33825.4]
  wire  output_51_33; // @[Switch.scala 41:38:@33826.4]
  wire  _T_72669; // @[Switch.scala 41:52:@33828.4]
  wire  output_51_34; // @[Switch.scala 41:38:@33829.4]
  wire  _T_72672; // @[Switch.scala 41:52:@33831.4]
  wire  output_51_35; // @[Switch.scala 41:38:@33832.4]
  wire  _T_72675; // @[Switch.scala 41:52:@33834.4]
  wire  output_51_36; // @[Switch.scala 41:38:@33835.4]
  wire  _T_72678; // @[Switch.scala 41:52:@33837.4]
  wire  output_51_37; // @[Switch.scala 41:38:@33838.4]
  wire  _T_72681; // @[Switch.scala 41:52:@33840.4]
  wire  output_51_38; // @[Switch.scala 41:38:@33841.4]
  wire  _T_72684; // @[Switch.scala 41:52:@33843.4]
  wire  output_51_39; // @[Switch.scala 41:38:@33844.4]
  wire  _T_72687; // @[Switch.scala 41:52:@33846.4]
  wire  output_51_40; // @[Switch.scala 41:38:@33847.4]
  wire  _T_72690; // @[Switch.scala 41:52:@33849.4]
  wire  output_51_41; // @[Switch.scala 41:38:@33850.4]
  wire  _T_72693; // @[Switch.scala 41:52:@33852.4]
  wire  output_51_42; // @[Switch.scala 41:38:@33853.4]
  wire  _T_72696; // @[Switch.scala 41:52:@33855.4]
  wire  output_51_43; // @[Switch.scala 41:38:@33856.4]
  wire  _T_72699; // @[Switch.scala 41:52:@33858.4]
  wire  output_51_44; // @[Switch.scala 41:38:@33859.4]
  wire  _T_72702; // @[Switch.scala 41:52:@33861.4]
  wire  output_51_45; // @[Switch.scala 41:38:@33862.4]
  wire  _T_72705; // @[Switch.scala 41:52:@33864.4]
  wire  output_51_46; // @[Switch.scala 41:38:@33865.4]
  wire  _T_72708; // @[Switch.scala 41:52:@33867.4]
  wire  output_51_47; // @[Switch.scala 41:38:@33868.4]
  wire  _T_72711; // @[Switch.scala 41:52:@33870.4]
  wire  output_51_48; // @[Switch.scala 41:38:@33871.4]
  wire  _T_72714; // @[Switch.scala 41:52:@33873.4]
  wire  output_51_49; // @[Switch.scala 41:38:@33874.4]
  wire  _T_72717; // @[Switch.scala 41:52:@33876.4]
  wire  output_51_50; // @[Switch.scala 41:38:@33877.4]
  wire  _T_72720; // @[Switch.scala 41:52:@33879.4]
  wire  output_51_51; // @[Switch.scala 41:38:@33880.4]
  wire  _T_72723; // @[Switch.scala 41:52:@33882.4]
  wire  output_51_52; // @[Switch.scala 41:38:@33883.4]
  wire  _T_72726; // @[Switch.scala 41:52:@33885.4]
  wire  output_51_53; // @[Switch.scala 41:38:@33886.4]
  wire  _T_72729; // @[Switch.scala 41:52:@33888.4]
  wire  output_51_54; // @[Switch.scala 41:38:@33889.4]
  wire  _T_72732; // @[Switch.scala 41:52:@33891.4]
  wire  output_51_55; // @[Switch.scala 41:38:@33892.4]
  wire  _T_72735; // @[Switch.scala 41:52:@33894.4]
  wire  output_51_56; // @[Switch.scala 41:38:@33895.4]
  wire  _T_72738; // @[Switch.scala 41:52:@33897.4]
  wire  output_51_57; // @[Switch.scala 41:38:@33898.4]
  wire  _T_72741; // @[Switch.scala 41:52:@33900.4]
  wire  output_51_58; // @[Switch.scala 41:38:@33901.4]
  wire  _T_72744; // @[Switch.scala 41:52:@33903.4]
  wire  output_51_59; // @[Switch.scala 41:38:@33904.4]
  wire  _T_72747; // @[Switch.scala 41:52:@33906.4]
  wire  output_51_60; // @[Switch.scala 41:38:@33907.4]
  wire  _T_72750; // @[Switch.scala 41:52:@33909.4]
  wire  output_51_61; // @[Switch.scala 41:38:@33910.4]
  wire  _T_72753; // @[Switch.scala 41:52:@33912.4]
  wire  output_51_62; // @[Switch.scala 41:38:@33913.4]
  wire  _T_72756; // @[Switch.scala 41:52:@33915.4]
  wire  output_51_63; // @[Switch.scala 41:38:@33916.4]
  wire [7:0] _T_72764; // @[Switch.scala 43:31:@33924.4]
  wire [15:0] _T_72772; // @[Switch.scala 43:31:@33932.4]
  wire [7:0] _T_72779; // @[Switch.scala 43:31:@33939.4]
  wire [31:0] _T_72788; // @[Switch.scala 43:31:@33948.4]
  wire [7:0] _T_72795; // @[Switch.scala 43:31:@33955.4]
  wire [15:0] _T_72803; // @[Switch.scala 43:31:@33963.4]
  wire [7:0] _T_72810; // @[Switch.scala 43:31:@33970.4]
  wire [31:0] _T_72819; // @[Switch.scala 43:31:@33979.4]
  wire [63:0] _T_72820; // @[Switch.scala 43:31:@33980.4]
  wire  _T_72824; // @[Switch.scala 41:52:@33983.4]
  wire  output_52_0; // @[Switch.scala 41:38:@33984.4]
  wire  _T_72827; // @[Switch.scala 41:52:@33986.4]
  wire  output_52_1; // @[Switch.scala 41:38:@33987.4]
  wire  _T_72830; // @[Switch.scala 41:52:@33989.4]
  wire  output_52_2; // @[Switch.scala 41:38:@33990.4]
  wire  _T_72833; // @[Switch.scala 41:52:@33992.4]
  wire  output_52_3; // @[Switch.scala 41:38:@33993.4]
  wire  _T_72836; // @[Switch.scala 41:52:@33995.4]
  wire  output_52_4; // @[Switch.scala 41:38:@33996.4]
  wire  _T_72839; // @[Switch.scala 41:52:@33998.4]
  wire  output_52_5; // @[Switch.scala 41:38:@33999.4]
  wire  _T_72842; // @[Switch.scala 41:52:@34001.4]
  wire  output_52_6; // @[Switch.scala 41:38:@34002.4]
  wire  _T_72845; // @[Switch.scala 41:52:@34004.4]
  wire  output_52_7; // @[Switch.scala 41:38:@34005.4]
  wire  _T_72848; // @[Switch.scala 41:52:@34007.4]
  wire  output_52_8; // @[Switch.scala 41:38:@34008.4]
  wire  _T_72851; // @[Switch.scala 41:52:@34010.4]
  wire  output_52_9; // @[Switch.scala 41:38:@34011.4]
  wire  _T_72854; // @[Switch.scala 41:52:@34013.4]
  wire  output_52_10; // @[Switch.scala 41:38:@34014.4]
  wire  _T_72857; // @[Switch.scala 41:52:@34016.4]
  wire  output_52_11; // @[Switch.scala 41:38:@34017.4]
  wire  _T_72860; // @[Switch.scala 41:52:@34019.4]
  wire  output_52_12; // @[Switch.scala 41:38:@34020.4]
  wire  _T_72863; // @[Switch.scala 41:52:@34022.4]
  wire  output_52_13; // @[Switch.scala 41:38:@34023.4]
  wire  _T_72866; // @[Switch.scala 41:52:@34025.4]
  wire  output_52_14; // @[Switch.scala 41:38:@34026.4]
  wire  _T_72869; // @[Switch.scala 41:52:@34028.4]
  wire  output_52_15; // @[Switch.scala 41:38:@34029.4]
  wire  _T_72872; // @[Switch.scala 41:52:@34031.4]
  wire  output_52_16; // @[Switch.scala 41:38:@34032.4]
  wire  _T_72875; // @[Switch.scala 41:52:@34034.4]
  wire  output_52_17; // @[Switch.scala 41:38:@34035.4]
  wire  _T_72878; // @[Switch.scala 41:52:@34037.4]
  wire  output_52_18; // @[Switch.scala 41:38:@34038.4]
  wire  _T_72881; // @[Switch.scala 41:52:@34040.4]
  wire  output_52_19; // @[Switch.scala 41:38:@34041.4]
  wire  _T_72884; // @[Switch.scala 41:52:@34043.4]
  wire  output_52_20; // @[Switch.scala 41:38:@34044.4]
  wire  _T_72887; // @[Switch.scala 41:52:@34046.4]
  wire  output_52_21; // @[Switch.scala 41:38:@34047.4]
  wire  _T_72890; // @[Switch.scala 41:52:@34049.4]
  wire  output_52_22; // @[Switch.scala 41:38:@34050.4]
  wire  _T_72893; // @[Switch.scala 41:52:@34052.4]
  wire  output_52_23; // @[Switch.scala 41:38:@34053.4]
  wire  _T_72896; // @[Switch.scala 41:52:@34055.4]
  wire  output_52_24; // @[Switch.scala 41:38:@34056.4]
  wire  _T_72899; // @[Switch.scala 41:52:@34058.4]
  wire  output_52_25; // @[Switch.scala 41:38:@34059.4]
  wire  _T_72902; // @[Switch.scala 41:52:@34061.4]
  wire  output_52_26; // @[Switch.scala 41:38:@34062.4]
  wire  _T_72905; // @[Switch.scala 41:52:@34064.4]
  wire  output_52_27; // @[Switch.scala 41:38:@34065.4]
  wire  _T_72908; // @[Switch.scala 41:52:@34067.4]
  wire  output_52_28; // @[Switch.scala 41:38:@34068.4]
  wire  _T_72911; // @[Switch.scala 41:52:@34070.4]
  wire  output_52_29; // @[Switch.scala 41:38:@34071.4]
  wire  _T_72914; // @[Switch.scala 41:52:@34073.4]
  wire  output_52_30; // @[Switch.scala 41:38:@34074.4]
  wire  _T_72917; // @[Switch.scala 41:52:@34076.4]
  wire  output_52_31; // @[Switch.scala 41:38:@34077.4]
  wire  _T_72920; // @[Switch.scala 41:52:@34079.4]
  wire  output_52_32; // @[Switch.scala 41:38:@34080.4]
  wire  _T_72923; // @[Switch.scala 41:52:@34082.4]
  wire  output_52_33; // @[Switch.scala 41:38:@34083.4]
  wire  _T_72926; // @[Switch.scala 41:52:@34085.4]
  wire  output_52_34; // @[Switch.scala 41:38:@34086.4]
  wire  _T_72929; // @[Switch.scala 41:52:@34088.4]
  wire  output_52_35; // @[Switch.scala 41:38:@34089.4]
  wire  _T_72932; // @[Switch.scala 41:52:@34091.4]
  wire  output_52_36; // @[Switch.scala 41:38:@34092.4]
  wire  _T_72935; // @[Switch.scala 41:52:@34094.4]
  wire  output_52_37; // @[Switch.scala 41:38:@34095.4]
  wire  _T_72938; // @[Switch.scala 41:52:@34097.4]
  wire  output_52_38; // @[Switch.scala 41:38:@34098.4]
  wire  _T_72941; // @[Switch.scala 41:52:@34100.4]
  wire  output_52_39; // @[Switch.scala 41:38:@34101.4]
  wire  _T_72944; // @[Switch.scala 41:52:@34103.4]
  wire  output_52_40; // @[Switch.scala 41:38:@34104.4]
  wire  _T_72947; // @[Switch.scala 41:52:@34106.4]
  wire  output_52_41; // @[Switch.scala 41:38:@34107.4]
  wire  _T_72950; // @[Switch.scala 41:52:@34109.4]
  wire  output_52_42; // @[Switch.scala 41:38:@34110.4]
  wire  _T_72953; // @[Switch.scala 41:52:@34112.4]
  wire  output_52_43; // @[Switch.scala 41:38:@34113.4]
  wire  _T_72956; // @[Switch.scala 41:52:@34115.4]
  wire  output_52_44; // @[Switch.scala 41:38:@34116.4]
  wire  _T_72959; // @[Switch.scala 41:52:@34118.4]
  wire  output_52_45; // @[Switch.scala 41:38:@34119.4]
  wire  _T_72962; // @[Switch.scala 41:52:@34121.4]
  wire  output_52_46; // @[Switch.scala 41:38:@34122.4]
  wire  _T_72965; // @[Switch.scala 41:52:@34124.4]
  wire  output_52_47; // @[Switch.scala 41:38:@34125.4]
  wire  _T_72968; // @[Switch.scala 41:52:@34127.4]
  wire  output_52_48; // @[Switch.scala 41:38:@34128.4]
  wire  _T_72971; // @[Switch.scala 41:52:@34130.4]
  wire  output_52_49; // @[Switch.scala 41:38:@34131.4]
  wire  _T_72974; // @[Switch.scala 41:52:@34133.4]
  wire  output_52_50; // @[Switch.scala 41:38:@34134.4]
  wire  _T_72977; // @[Switch.scala 41:52:@34136.4]
  wire  output_52_51; // @[Switch.scala 41:38:@34137.4]
  wire  _T_72980; // @[Switch.scala 41:52:@34139.4]
  wire  output_52_52; // @[Switch.scala 41:38:@34140.4]
  wire  _T_72983; // @[Switch.scala 41:52:@34142.4]
  wire  output_52_53; // @[Switch.scala 41:38:@34143.4]
  wire  _T_72986; // @[Switch.scala 41:52:@34145.4]
  wire  output_52_54; // @[Switch.scala 41:38:@34146.4]
  wire  _T_72989; // @[Switch.scala 41:52:@34148.4]
  wire  output_52_55; // @[Switch.scala 41:38:@34149.4]
  wire  _T_72992; // @[Switch.scala 41:52:@34151.4]
  wire  output_52_56; // @[Switch.scala 41:38:@34152.4]
  wire  _T_72995; // @[Switch.scala 41:52:@34154.4]
  wire  output_52_57; // @[Switch.scala 41:38:@34155.4]
  wire  _T_72998; // @[Switch.scala 41:52:@34157.4]
  wire  output_52_58; // @[Switch.scala 41:38:@34158.4]
  wire  _T_73001; // @[Switch.scala 41:52:@34160.4]
  wire  output_52_59; // @[Switch.scala 41:38:@34161.4]
  wire  _T_73004; // @[Switch.scala 41:52:@34163.4]
  wire  output_52_60; // @[Switch.scala 41:38:@34164.4]
  wire  _T_73007; // @[Switch.scala 41:52:@34166.4]
  wire  output_52_61; // @[Switch.scala 41:38:@34167.4]
  wire  _T_73010; // @[Switch.scala 41:52:@34169.4]
  wire  output_52_62; // @[Switch.scala 41:38:@34170.4]
  wire  _T_73013; // @[Switch.scala 41:52:@34172.4]
  wire  output_52_63; // @[Switch.scala 41:38:@34173.4]
  wire [7:0] _T_73021; // @[Switch.scala 43:31:@34181.4]
  wire [15:0] _T_73029; // @[Switch.scala 43:31:@34189.4]
  wire [7:0] _T_73036; // @[Switch.scala 43:31:@34196.4]
  wire [31:0] _T_73045; // @[Switch.scala 43:31:@34205.4]
  wire [7:0] _T_73052; // @[Switch.scala 43:31:@34212.4]
  wire [15:0] _T_73060; // @[Switch.scala 43:31:@34220.4]
  wire [7:0] _T_73067; // @[Switch.scala 43:31:@34227.4]
  wire [31:0] _T_73076; // @[Switch.scala 43:31:@34236.4]
  wire [63:0] _T_73077; // @[Switch.scala 43:31:@34237.4]
  wire  _T_73081; // @[Switch.scala 41:52:@34240.4]
  wire  output_53_0; // @[Switch.scala 41:38:@34241.4]
  wire  _T_73084; // @[Switch.scala 41:52:@34243.4]
  wire  output_53_1; // @[Switch.scala 41:38:@34244.4]
  wire  _T_73087; // @[Switch.scala 41:52:@34246.4]
  wire  output_53_2; // @[Switch.scala 41:38:@34247.4]
  wire  _T_73090; // @[Switch.scala 41:52:@34249.4]
  wire  output_53_3; // @[Switch.scala 41:38:@34250.4]
  wire  _T_73093; // @[Switch.scala 41:52:@34252.4]
  wire  output_53_4; // @[Switch.scala 41:38:@34253.4]
  wire  _T_73096; // @[Switch.scala 41:52:@34255.4]
  wire  output_53_5; // @[Switch.scala 41:38:@34256.4]
  wire  _T_73099; // @[Switch.scala 41:52:@34258.4]
  wire  output_53_6; // @[Switch.scala 41:38:@34259.4]
  wire  _T_73102; // @[Switch.scala 41:52:@34261.4]
  wire  output_53_7; // @[Switch.scala 41:38:@34262.4]
  wire  _T_73105; // @[Switch.scala 41:52:@34264.4]
  wire  output_53_8; // @[Switch.scala 41:38:@34265.4]
  wire  _T_73108; // @[Switch.scala 41:52:@34267.4]
  wire  output_53_9; // @[Switch.scala 41:38:@34268.4]
  wire  _T_73111; // @[Switch.scala 41:52:@34270.4]
  wire  output_53_10; // @[Switch.scala 41:38:@34271.4]
  wire  _T_73114; // @[Switch.scala 41:52:@34273.4]
  wire  output_53_11; // @[Switch.scala 41:38:@34274.4]
  wire  _T_73117; // @[Switch.scala 41:52:@34276.4]
  wire  output_53_12; // @[Switch.scala 41:38:@34277.4]
  wire  _T_73120; // @[Switch.scala 41:52:@34279.4]
  wire  output_53_13; // @[Switch.scala 41:38:@34280.4]
  wire  _T_73123; // @[Switch.scala 41:52:@34282.4]
  wire  output_53_14; // @[Switch.scala 41:38:@34283.4]
  wire  _T_73126; // @[Switch.scala 41:52:@34285.4]
  wire  output_53_15; // @[Switch.scala 41:38:@34286.4]
  wire  _T_73129; // @[Switch.scala 41:52:@34288.4]
  wire  output_53_16; // @[Switch.scala 41:38:@34289.4]
  wire  _T_73132; // @[Switch.scala 41:52:@34291.4]
  wire  output_53_17; // @[Switch.scala 41:38:@34292.4]
  wire  _T_73135; // @[Switch.scala 41:52:@34294.4]
  wire  output_53_18; // @[Switch.scala 41:38:@34295.4]
  wire  _T_73138; // @[Switch.scala 41:52:@34297.4]
  wire  output_53_19; // @[Switch.scala 41:38:@34298.4]
  wire  _T_73141; // @[Switch.scala 41:52:@34300.4]
  wire  output_53_20; // @[Switch.scala 41:38:@34301.4]
  wire  _T_73144; // @[Switch.scala 41:52:@34303.4]
  wire  output_53_21; // @[Switch.scala 41:38:@34304.4]
  wire  _T_73147; // @[Switch.scala 41:52:@34306.4]
  wire  output_53_22; // @[Switch.scala 41:38:@34307.4]
  wire  _T_73150; // @[Switch.scala 41:52:@34309.4]
  wire  output_53_23; // @[Switch.scala 41:38:@34310.4]
  wire  _T_73153; // @[Switch.scala 41:52:@34312.4]
  wire  output_53_24; // @[Switch.scala 41:38:@34313.4]
  wire  _T_73156; // @[Switch.scala 41:52:@34315.4]
  wire  output_53_25; // @[Switch.scala 41:38:@34316.4]
  wire  _T_73159; // @[Switch.scala 41:52:@34318.4]
  wire  output_53_26; // @[Switch.scala 41:38:@34319.4]
  wire  _T_73162; // @[Switch.scala 41:52:@34321.4]
  wire  output_53_27; // @[Switch.scala 41:38:@34322.4]
  wire  _T_73165; // @[Switch.scala 41:52:@34324.4]
  wire  output_53_28; // @[Switch.scala 41:38:@34325.4]
  wire  _T_73168; // @[Switch.scala 41:52:@34327.4]
  wire  output_53_29; // @[Switch.scala 41:38:@34328.4]
  wire  _T_73171; // @[Switch.scala 41:52:@34330.4]
  wire  output_53_30; // @[Switch.scala 41:38:@34331.4]
  wire  _T_73174; // @[Switch.scala 41:52:@34333.4]
  wire  output_53_31; // @[Switch.scala 41:38:@34334.4]
  wire  _T_73177; // @[Switch.scala 41:52:@34336.4]
  wire  output_53_32; // @[Switch.scala 41:38:@34337.4]
  wire  _T_73180; // @[Switch.scala 41:52:@34339.4]
  wire  output_53_33; // @[Switch.scala 41:38:@34340.4]
  wire  _T_73183; // @[Switch.scala 41:52:@34342.4]
  wire  output_53_34; // @[Switch.scala 41:38:@34343.4]
  wire  _T_73186; // @[Switch.scala 41:52:@34345.4]
  wire  output_53_35; // @[Switch.scala 41:38:@34346.4]
  wire  _T_73189; // @[Switch.scala 41:52:@34348.4]
  wire  output_53_36; // @[Switch.scala 41:38:@34349.4]
  wire  _T_73192; // @[Switch.scala 41:52:@34351.4]
  wire  output_53_37; // @[Switch.scala 41:38:@34352.4]
  wire  _T_73195; // @[Switch.scala 41:52:@34354.4]
  wire  output_53_38; // @[Switch.scala 41:38:@34355.4]
  wire  _T_73198; // @[Switch.scala 41:52:@34357.4]
  wire  output_53_39; // @[Switch.scala 41:38:@34358.4]
  wire  _T_73201; // @[Switch.scala 41:52:@34360.4]
  wire  output_53_40; // @[Switch.scala 41:38:@34361.4]
  wire  _T_73204; // @[Switch.scala 41:52:@34363.4]
  wire  output_53_41; // @[Switch.scala 41:38:@34364.4]
  wire  _T_73207; // @[Switch.scala 41:52:@34366.4]
  wire  output_53_42; // @[Switch.scala 41:38:@34367.4]
  wire  _T_73210; // @[Switch.scala 41:52:@34369.4]
  wire  output_53_43; // @[Switch.scala 41:38:@34370.4]
  wire  _T_73213; // @[Switch.scala 41:52:@34372.4]
  wire  output_53_44; // @[Switch.scala 41:38:@34373.4]
  wire  _T_73216; // @[Switch.scala 41:52:@34375.4]
  wire  output_53_45; // @[Switch.scala 41:38:@34376.4]
  wire  _T_73219; // @[Switch.scala 41:52:@34378.4]
  wire  output_53_46; // @[Switch.scala 41:38:@34379.4]
  wire  _T_73222; // @[Switch.scala 41:52:@34381.4]
  wire  output_53_47; // @[Switch.scala 41:38:@34382.4]
  wire  _T_73225; // @[Switch.scala 41:52:@34384.4]
  wire  output_53_48; // @[Switch.scala 41:38:@34385.4]
  wire  _T_73228; // @[Switch.scala 41:52:@34387.4]
  wire  output_53_49; // @[Switch.scala 41:38:@34388.4]
  wire  _T_73231; // @[Switch.scala 41:52:@34390.4]
  wire  output_53_50; // @[Switch.scala 41:38:@34391.4]
  wire  _T_73234; // @[Switch.scala 41:52:@34393.4]
  wire  output_53_51; // @[Switch.scala 41:38:@34394.4]
  wire  _T_73237; // @[Switch.scala 41:52:@34396.4]
  wire  output_53_52; // @[Switch.scala 41:38:@34397.4]
  wire  _T_73240; // @[Switch.scala 41:52:@34399.4]
  wire  output_53_53; // @[Switch.scala 41:38:@34400.4]
  wire  _T_73243; // @[Switch.scala 41:52:@34402.4]
  wire  output_53_54; // @[Switch.scala 41:38:@34403.4]
  wire  _T_73246; // @[Switch.scala 41:52:@34405.4]
  wire  output_53_55; // @[Switch.scala 41:38:@34406.4]
  wire  _T_73249; // @[Switch.scala 41:52:@34408.4]
  wire  output_53_56; // @[Switch.scala 41:38:@34409.4]
  wire  _T_73252; // @[Switch.scala 41:52:@34411.4]
  wire  output_53_57; // @[Switch.scala 41:38:@34412.4]
  wire  _T_73255; // @[Switch.scala 41:52:@34414.4]
  wire  output_53_58; // @[Switch.scala 41:38:@34415.4]
  wire  _T_73258; // @[Switch.scala 41:52:@34417.4]
  wire  output_53_59; // @[Switch.scala 41:38:@34418.4]
  wire  _T_73261; // @[Switch.scala 41:52:@34420.4]
  wire  output_53_60; // @[Switch.scala 41:38:@34421.4]
  wire  _T_73264; // @[Switch.scala 41:52:@34423.4]
  wire  output_53_61; // @[Switch.scala 41:38:@34424.4]
  wire  _T_73267; // @[Switch.scala 41:52:@34426.4]
  wire  output_53_62; // @[Switch.scala 41:38:@34427.4]
  wire  _T_73270; // @[Switch.scala 41:52:@34429.4]
  wire  output_53_63; // @[Switch.scala 41:38:@34430.4]
  wire [7:0] _T_73278; // @[Switch.scala 43:31:@34438.4]
  wire [15:0] _T_73286; // @[Switch.scala 43:31:@34446.4]
  wire [7:0] _T_73293; // @[Switch.scala 43:31:@34453.4]
  wire [31:0] _T_73302; // @[Switch.scala 43:31:@34462.4]
  wire [7:0] _T_73309; // @[Switch.scala 43:31:@34469.4]
  wire [15:0] _T_73317; // @[Switch.scala 43:31:@34477.4]
  wire [7:0] _T_73324; // @[Switch.scala 43:31:@34484.4]
  wire [31:0] _T_73333; // @[Switch.scala 43:31:@34493.4]
  wire [63:0] _T_73334; // @[Switch.scala 43:31:@34494.4]
  wire  _T_73338; // @[Switch.scala 41:52:@34497.4]
  wire  output_54_0; // @[Switch.scala 41:38:@34498.4]
  wire  _T_73341; // @[Switch.scala 41:52:@34500.4]
  wire  output_54_1; // @[Switch.scala 41:38:@34501.4]
  wire  _T_73344; // @[Switch.scala 41:52:@34503.4]
  wire  output_54_2; // @[Switch.scala 41:38:@34504.4]
  wire  _T_73347; // @[Switch.scala 41:52:@34506.4]
  wire  output_54_3; // @[Switch.scala 41:38:@34507.4]
  wire  _T_73350; // @[Switch.scala 41:52:@34509.4]
  wire  output_54_4; // @[Switch.scala 41:38:@34510.4]
  wire  _T_73353; // @[Switch.scala 41:52:@34512.4]
  wire  output_54_5; // @[Switch.scala 41:38:@34513.4]
  wire  _T_73356; // @[Switch.scala 41:52:@34515.4]
  wire  output_54_6; // @[Switch.scala 41:38:@34516.4]
  wire  _T_73359; // @[Switch.scala 41:52:@34518.4]
  wire  output_54_7; // @[Switch.scala 41:38:@34519.4]
  wire  _T_73362; // @[Switch.scala 41:52:@34521.4]
  wire  output_54_8; // @[Switch.scala 41:38:@34522.4]
  wire  _T_73365; // @[Switch.scala 41:52:@34524.4]
  wire  output_54_9; // @[Switch.scala 41:38:@34525.4]
  wire  _T_73368; // @[Switch.scala 41:52:@34527.4]
  wire  output_54_10; // @[Switch.scala 41:38:@34528.4]
  wire  _T_73371; // @[Switch.scala 41:52:@34530.4]
  wire  output_54_11; // @[Switch.scala 41:38:@34531.4]
  wire  _T_73374; // @[Switch.scala 41:52:@34533.4]
  wire  output_54_12; // @[Switch.scala 41:38:@34534.4]
  wire  _T_73377; // @[Switch.scala 41:52:@34536.4]
  wire  output_54_13; // @[Switch.scala 41:38:@34537.4]
  wire  _T_73380; // @[Switch.scala 41:52:@34539.4]
  wire  output_54_14; // @[Switch.scala 41:38:@34540.4]
  wire  _T_73383; // @[Switch.scala 41:52:@34542.4]
  wire  output_54_15; // @[Switch.scala 41:38:@34543.4]
  wire  _T_73386; // @[Switch.scala 41:52:@34545.4]
  wire  output_54_16; // @[Switch.scala 41:38:@34546.4]
  wire  _T_73389; // @[Switch.scala 41:52:@34548.4]
  wire  output_54_17; // @[Switch.scala 41:38:@34549.4]
  wire  _T_73392; // @[Switch.scala 41:52:@34551.4]
  wire  output_54_18; // @[Switch.scala 41:38:@34552.4]
  wire  _T_73395; // @[Switch.scala 41:52:@34554.4]
  wire  output_54_19; // @[Switch.scala 41:38:@34555.4]
  wire  _T_73398; // @[Switch.scala 41:52:@34557.4]
  wire  output_54_20; // @[Switch.scala 41:38:@34558.4]
  wire  _T_73401; // @[Switch.scala 41:52:@34560.4]
  wire  output_54_21; // @[Switch.scala 41:38:@34561.4]
  wire  _T_73404; // @[Switch.scala 41:52:@34563.4]
  wire  output_54_22; // @[Switch.scala 41:38:@34564.4]
  wire  _T_73407; // @[Switch.scala 41:52:@34566.4]
  wire  output_54_23; // @[Switch.scala 41:38:@34567.4]
  wire  _T_73410; // @[Switch.scala 41:52:@34569.4]
  wire  output_54_24; // @[Switch.scala 41:38:@34570.4]
  wire  _T_73413; // @[Switch.scala 41:52:@34572.4]
  wire  output_54_25; // @[Switch.scala 41:38:@34573.4]
  wire  _T_73416; // @[Switch.scala 41:52:@34575.4]
  wire  output_54_26; // @[Switch.scala 41:38:@34576.4]
  wire  _T_73419; // @[Switch.scala 41:52:@34578.4]
  wire  output_54_27; // @[Switch.scala 41:38:@34579.4]
  wire  _T_73422; // @[Switch.scala 41:52:@34581.4]
  wire  output_54_28; // @[Switch.scala 41:38:@34582.4]
  wire  _T_73425; // @[Switch.scala 41:52:@34584.4]
  wire  output_54_29; // @[Switch.scala 41:38:@34585.4]
  wire  _T_73428; // @[Switch.scala 41:52:@34587.4]
  wire  output_54_30; // @[Switch.scala 41:38:@34588.4]
  wire  _T_73431; // @[Switch.scala 41:52:@34590.4]
  wire  output_54_31; // @[Switch.scala 41:38:@34591.4]
  wire  _T_73434; // @[Switch.scala 41:52:@34593.4]
  wire  output_54_32; // @[Switch.scala 41:38:@34594.4]
  wire  _T_73437; // @[Switch.scala 41:52:@34596.4]
  wire  output_54_33; // @[Switch.scala 41:38:@34597.4]
  wire  _T_73440; // @[Switch.scala 41:52:@34599.4]
  wire  output_54_34; // @[Switch.scala 41:38:@34600.4]
  wire  _T_73443; // @[Switch.scala 41:52:@34602.4]
  wire  output_54_35; // @[Switch.scala 41:38:@34603.4]
  wire  _T_73446; // @[Switch.scala 41:52:@34605.4]
  wire  output_54_36; // @[Switch.scala 41:38:@34606.4]
  wire  _T_73449; // @[Switch.scala 41:52:@34608.4]
  wire  output_54_37; // @[Switch.scala 41:38:@34609.4]
  wire  _T_73452; // @[Switch.scala 41:52:@34611.4]
  wire  output_54_38; // @[Switch.scala 41:38:@34612.4]
  wire  _T_73455; // @[Switch.scala 41:52:@34614.4]
  wire  output_54_39; // @[Switch.scala 41:38:@34615.4]
  wire  _T_73458; // @[Switch.scala 41:52:@34617.4]
  wire  output_54_40; // @[Switch.scala 41:38:@34618.4]
  wire  _T_73461; // @[Switch.scala 41:52:@34620.4]
  wire  output_54_41; // @[Switch.scala 41:38:@34621.4]
  wire  _T_73464; // @[Switch.scala 41:52:@34623.4]
  wire  output_54_42; // @[Switch.scala 41:38:@34624.4]
  wire  _T_73467; // @[Switch.scala 41:52:@34626.4]
  wire  output_54_43; // @[Switch.scala 41:38:@34627.4]
  wire  _T_73470; // @[Switch.scala 41:52:@34629.4]
  wire  output_54_44; // @[Switch.scala 41:38:@34630.4]
  wire  _T_73473; // @[Switch.scala 41:52:@34632.4]
  wire  output_54_45; // @[Switch.scala 41:38:@34633.4]
  wire  _T_73476; // @[Switch.scala 41:52:@34635.4]
  wire  output_54_46; // @[Switch.scala 41:38:@34636.4]
  wire  _T_73479; // @[Switch.scala 41:52:@34638.4]
  wire  output_54_47; // @[Switch.scala 41:38:@34639.4]
  wire  _T_73482; // @[Switch.scala 41:52:@34641.4]
  wire  output_54_48; // @[Switch.scala 41:38:@34642.4]
  wire  _T_73485; // @[Switch.scala 41:52:@34644.4]
  wire  output_54_49; // @[Switch.scala 41:38:@34645.4]
  wire  _T_73488; // @[Switch.scala 41:52:@34647.4]
  wire  output_54_50; // @[Switch.scala 41:38:@34648.4]
  wire  _T_73491; // @[Switch.scala 41:52:@34650.4]
  wire  output_54_51; // @[Switch.scala 41:38:@34651.4]
  wire  _T_73494; // @[Switch.scala 41:52:@34653.4]
  wire  output_54_52; // @[Switch.scala 41:38:@34654.4]
  wire  _T_73497; // @[Switch.scala 41:52:@34656.4]
  wire  output_54_53; // @[Switch.scala 41:38:@34657.4]
  wire  _T_73500; // @[Switch.scala 41:52:@34659.4]
  wire  output_54_54; // @[Switch.scala 41:38:@34660.4]
  wire  _T_73503; // @[Switch.scala 41:52:@34662.4]
  wire  output_54_55; // @[Switch.scala 41:38:@34663.4]
  wire  _T_73506; // @[Switch.scala 41:52:@34665.4]
  wire  output_54_56; // @[Switch.scala 41:38:@34666.4]
  wire  _T_73509; // @[Switch.scala 41:52:@34668.4]
  wire  output_54_57; // @[Switch.scala 41:38:@34669.4]
  wire  _T_73512; // @[Switch.scala 41:52:@34671.4]
  wire  output_54_58; // @[Switch.scala 41:38:@34672.4]
  wire  _T_73515; // @[Switch.scala 41:52:@34674.4]
  wire  output_54_59; // @[Switch.scala 41:38:@34675.4]
  wire  _T_73518; // @[Switch.scala 41:52:@34677.4]
  wire  output_54_60; // @[Switch.scala 41:38:@34678.4]
  wire  _T_73521; // @[Switch.scala 41:52:@34680.4]
  wire  output_54_61; // @[Switch.scala 41:38:@34681.4]
  wire  _T_73524; // @[Switch.scala 41:52:@34683.4]
  wire  output_54_62; // @[Switch.scala 41:38:@34684.4]
  wire  _T_73527; // @[Switch.scala 41:52:@34686.4]
  wire  output_54_63; // @[Switch.scala 41:38:@34687.4]
  wire [7:0] _T_73535; // @[Switch.scala 43:31:@34695.4]
  wire [15:0] _T_73543; // @[Switch.scala 43:31:@34703.4]
  wire [7:0] _T_73550; // @[Switch.scala 43:31:@34710.4]
  wire [31:0] _T_73559; // @[Switch.scala 43:31:@34719.4]
  wire [7:0] _T_73566; // @[Switch.scala 43:31:@34726.4]
  wire [15:0] _T_73574; // @[Switch.scala 43:31:@34734.4]
  wire [7:0] _T_73581; // @[Switch.scala 43:31:@34741.4]
  wire [31:0] _T_73590; // @[Switch.scala 43:31:@34750.4]
  wire [63:0] _T_73591; // @[Switch.scala 43:31:@34751.4]
  wire  _T_73595; // @[Switch.scala 41:52:@34754.4]
  wire  output_55_0; // @[Switch.scala 41:38:@34755.4]
  wire  _T_73598; // @[Switch.scala 41:52:@34757.4]
  wire  output_55_1; // @[Switch.scala 41:38:@34758.4]
  wire  _T_73601; // @[Switch.scala 41:52:@34760.4]
  wire  output_55_2; // @[Switch.scala 41:38:@34761.4]
  wire  _T_73604; // @[Switch.scala 41:52:@34763.4]
  wire  output_55_3; // @[Switch.scala 41:38:@34764.4]
  wire  _T_73607; // @[Switch.scala 41:52:@34766.4]
  wire  output_55_4; // @[Switch.scala 41:38:@34767.4]
  wire  _T_73610; // @[Switch.scala 41:52:@34769.4]
  wire  output_55_5; // @[Switch.scala 41:38:@34770.4]
  wire  _T_73613; // @[Switch.scala 41:52:@34772.4]
  wire  output_55_6; // @[Switch.scala 41:38:@34773.4]
  wire  _T_73616; // @[Switch.scala 41:52:@34775.4]
  wire  output_55_7; // @[Switch.scala 41:38:@34776.4]
  wire  _T_73619; // @[Switch.scala 41:52:@34778.4]
  wire  output_55_8; // @[Switch.scala 41:38:@34779.4]
  wire  _T_73622; // @[Switch.scala 41:52:@34781.4]
  wire  output_55_9; // @[Switch.scala 41:38:@34782.4]
  wire  _T_73625; // @[Switch.scala 41:52:@34784.4]
  wire  output_55_10; // @[Switch.scala 41:38:@34785.4]
  wire  _T_73628; // @[Switch.scala 41:52:@34787.4]
  wire  output_55_11; // @[Switch.scala 41:38:@34788.4]
  wire  _T_73631; // @[Switch.scala 41:52:@34790.4]
  wire  output_55_12; // @[Switch.scala 41:38:@34791.4]
  wire  _T_73634; // @[Switch.scala 41:52:@34793.4]
  wire  output_55_13; // @[Switch.scala 41:38:@34794.4]
  wire  _T_73637; // @[Switch.scala 41:52:@34796.4]
  wire  output_55_14; // @[Switch.scala 41:38:@34797.4]
  wire  _T_73640; // @[Switch.scala 41:52:@34799.4]
  wire  output_55_15; // @[Switch.scala 41:38:@34800.4]
  wire  _T_73643; // @[Switch.scala 41:52:@34802.4]
  wire  output_55_16; // @[Switch.scala 41:38:@34803.4]
  wire  _T_73646; // @[Switch.scala 41:52:@34805.4]
  wire  output_55_17; // @[Switch.scala 41:38:@34806.4]
  wire  _T_73649; // @[Switch.scala 41:52:@34808.4]
  wire  output_55_18; // @[Switch.scala 41:38:@34809.4]
  wire  _T_73652; // @[Switch.scala 41:52:@34811.4]
  wire  output_55_19; // @[Switch.scala 41:38:@34812.4]
  wire  _T_73655; // @[Switch.scala 41:52:@34814.4]
  wire  output_55_20; // @[Switch.scala 41:38:@34815.4]
  wire  _T_73658; // @[Switch.scala 41:52:@34817.4]
  wire  output_55_21; // @[Switch.scala 41:38:@34818.4]
  wire  _T_73661; // @[Switch.scala 41:52:@34820.4]
  wire  output_55_22; // @[Switch.scala 41:38:@34821.4]
  wire  _T_73664; // @[Switch.scala 41:52:@34823.4]
  wire  output_55_23; // @[Switch.scala 41:38:@34824.4]
  wire  _T_73667; // @[Switch.scala 41:52:@34826.4]
  wire  output_55_24; // @[Switch.scala 41:38:@34827.4]
  wire  _T_73670; // @[Switch.scala 41:52:@34829.4]
  wire  output_55_25; // @[Switch.scala 41:38:@34830.4]
  wire  _T_73673; // @[Switch.scala 41:52:@34832.4]
  wire  output_55_26; // @[Switch.scala 41:38:@34833.4]
  wire  _T_73676; // @[Switch.scala 41:52:@34835.4]
  wire  output_55_27; // @[Switch.scala 41:38:@34836.4]
  wire  _T_73679; // @[Switch.scala 41:52:@34838.4]
  wire  output_55_28; // @[Switch.scala 41:38:@34839.4]
  wire  _T_73682; // @[Switch.scala 41:52:@34841.4]
  wire  output_55_29; // @[Switch.scala 41:38:@34842.4]
  wire  _T_73685; // @[Switch.scala 41:52:@34844.4]
  wire  output_55_30; // @[Switch.scala 41:38:@34845.4]
  wire  _T_73688; // @[Switch.scala 41:52:@34847.4]
  wire  output_55_31; // @[Switch.scala 41:38:@34848.4]
  wire  _T_73691; // @[Switch.scala 41:52:@34850.4]
  wire  output_55_32; // @[Switch.scala 41:38:@34851.4]
  wire  _T_73694; // @[Switch.scala 41:52:@34853.4]
  wire  output_55_33; // @[Switch.scala 41:38:@34854.4]
  wire  _T_73697; // @[Switch.scala 41:52:@34856.4]
  wire  output_55_34; // @[Switch.scala 41:38:@34857.4]
  wire  _T_73700; // @[Switch.scala 41:52:@34859.4]
  wire  output_55_35; // @[Switch.scala 41:38:@34860.4]
  wire  _T_73703; // @[Switch.scala 41:52:@34862.4]
  wire  output_55_36; // @[Switch.scala 41:38:@34863.4]
  wire  _T_73706; // @[Switch.scala 41:52:@34865.4]
  wire  output_55_37; // @[Switch.scala 41:38:@34866.4]
  wire  _T_73709; // @[Switch.scala 41:52:@34868.4]
  wire  output_55_38; // @[Switch.scala 41:38:@34869.4]
  wire  _T_73712; // @[Switch.scala 41:52:@34871.4]
  wire  output_55_39; // @[Switch.scala 41:38:@34872.4]
  wire  _T_73715; // @[Switch.scala 41:52:@34874.4]
  wire  output_55_40; // @[Switch.scala 41:38:@34875.4]
  wire  _T_73718; // @[Switch.scala 41:52:@34877.4]
  wire  output_55_41; // @[Switch.scala 41:38:@34878.4]
  wire  _T_73721; // @[Switch.scala 41:52:@34880.4]
  wire  output_55_42; // @[Switch.scala 41:38:@34881.4]
  wire  _T_73724; // @[Switch.scala 41:52:@34883.4]
  wire  output_55_43; // @[Switch.scala 41:38:@34884.4]
  wire  _T_73727; // @[Switch.scala 41:52:@34886.4]
  wire  output_55_44; // @[Switch.scala 41:38:@34887.4]
  wire  _T_73730; // @[Switch.scala 41:52:@34889.4]
  wire  output_55_45; // @[Switch.scala 41:38:@34890.4]
  wire  _T_73733; // @[Switch.scala 41:52:@34892.4]
  wire  output_55_46; // @[Switch.scala 41:38:@34893.4]
  wire  _T_73736; // @[Switch.scala 41:52:@34895.4]
  wire  output_55_47; // @[Switch.scala 41:38:@34896.4]
  wire  _T_73739; // @[Switch.scala 41:52:@34898.4]
  wire  output_55_48; // @[Switch.scala 41:38:@34899.4]
  wire  _T_73742; // @[Switch.scala 41:52:@34901.4]
  wire  output_55_49; // @[Switch.scala 41:38:@34902.4]
  wire  _T_73745; // @[Switch.scala 41:52:@34904.4]
  wire  output_55_50; // @[Switch.scala 41:38:@34905.4]
  wire  _T_73748; // @[Switch.scala 41:52:@34907.4]
  wire  output_55_51; // @[Switch.scala 41:38:@34908.4]
  wire  _T_73751; // @[Switch.scala 41:52:@34910.4]
  wire  output_55_52; // @[Switch.scala 41:38:@34911.4]
  wire  _T_73754; // @[Switch.scala 41:52:@34913.4]
  wire  output_55_53; // @[Switch.scala 41:38:@34914.4]
  wire  _T_73757; // @[Switch.scala 41:52:@34916.4]
  wire  output_55_54; // @[Switch.scala 41:38:@34917.4]
  wire  _T_73760; // @[Switch.scala 41:52:@34919.4]
  wire  output_55_55; // @[Switch.scala 41:38:@34920.4]
  wire  _T_73763; // @[Switch.scala 41:52:@34922.4]
  wire  output_55_56; // @[Switch.scala 41:38:@34923.4]
  wire  _T_73766; // @[Switch.scala 41:52:@34925.4]
  wire  output_55_57; // @[Switch.scala 41:38:@34926.4]
  wire  _T_73769; // @[Switch.scala 41:52:@34928.4]
  wire  output_55_58; // @[Switch.scala 41:38:@34929.4]
  wire  _T_73772; // @[Switch.scala 41:52:@34931.4]
  wire  output_55_59; // @[Switch.scala 41:38:@34932.4]
  wire  _T_73775; // @[Switch.scala 41:52:@34934.4]
  wire  output_55_60; // @[Switch.scala 41:38:@34935.4]
  wire  _T_73778; // @[Switch.scala 41:52:@34937.4]
  wire  output_55_61; // @[Switch.scala 41:38:@34938.4]
  wire  _T_73781; // @[Switch.scala 41:52:@34940.4]
  wire  output_55_62; // @[Switch.scala 41:38:@34941.4]
  wire  _T_73784; // @[Switch.scala 41:52:@34943.4]
  wire  output_55_63; // @[Switch.scala 41:38:@34944.4]
  wire [7:0] _T_73792; // @[Switch.scala 43:31:@34952.4]
  wire [15:0] _T_73800; // @[Switch.scala 43:31:@34960.4]
  wire [7:0] _T_73807; // @[Switch.scala 43:31:@34967.4]
  wire [31:0] _T_73816; // @[Switch.scala 43:31:@34976.4]
  wire [7:0] _T_73823; // @[Switch.scala 43:31:@34983.4]
  wire [15:0] _T_73831; // @[Switch.scala 43:31:@34991.4]
  wire [7:0] _T_73838; // @[Switch.scala 43:31:@34998.4]
  wire [31:0] _T_73847; // @[Switch.scala 43:31:@35007.4]
  wire [63:0] _T_73848; // @[Switch.scala 43:31:@35008.4]
  wire  _T_73852; // @[Switch.scala 41:52:@35011.4]
  wire  output_56_0; // @[Switch.scala 41:38:@35012.4]
  wire  _T_73855; // @[Switch.scala 41:52:@35014.4]
  wire  output_56_1; // @[Switch.scala 41:38:@35015.4]
  wire  _T_73858; // @[Switch.scala 41:52:@35017.4]
  wire  output_56_2; // @[Switch.scala 41:38:@35018.4]
  wire  _T_73861; // @[Switch.scala 41:52:@35020.4]
  wire  output_56_3; // @[Switch.scala 41:38:@35021.4]
  wire  _T_73864; // @[Switch.scala 41:52:@35023.4]
  wire  output_56_4; // @[Switch.scala 41:38:@35024.4]
  wire  _T_73867; // @[Switch.scala 41:52:@35026.4]
  wire  output_56_5; // @[Switch.scala 41:38:@35027.4]
  wire  _T_73870; // @[Switch.scala 41:52:@35029.4]
  wire  output_56_6; // @[Switch.scala 41:38:@35030.4]
  wire  _T_73873; // @[Switch.scala 41:52:@35032.4]
  wire  output_56_7; // @[Switch.scala 41:38:@35033.4]
  wire  _T_73876; // @[Switch.scala 41:52:@35035.4]
  wire  output_56_8; // @[Switch.scala 41:38:@35036.4]
  wire  _T_73879; // @[Switch.scala 41:52:@35038.4]
  wire  output_56_9; // @[Switch.scala 41:38:@35039.4]
  wire  _T_73882; // @[Switch.scala 41:52:@35041.4]
  wire  output_56_10; // @[Switch.scala 41:38:@35042.4]
  wire  _T_73885; // @[Switch.scala 41:52:@35044.4]
  wire  output_56_11; // @[Switch.scala 41:38:@35045.4]
  wire  _T_73888; // @[Switch.scala 41:52:@35047.4]
  wire  output_56_12; // @[Switch.scala 41:38:@35048.4]
  wire  _T_73891; // @[Switch.scala 41:52:@35050.4]
  wire  output_56_13; // @[Switch.scala 41:38:@35051.4]
  wire  _T_73894; // @[Switch.scala 41:52:@35053.4]
  wire  output_56_14; // @[Switch.scala 41:38:@35054.4]
  wire  _T_73897; // @[Switch.scala 41:52:@35056.4]
  wire  output_56_15; // @[Switch.scala 41:38:@35057.4]
  wire  _T_73900; // @[Switch.scala 41:52:@35059.4]
  wire  output_56_16; // @[Switch.scala 41:38:@35060.4]
  wire  _T_73903; // @[Switch.scala 41:52:@35062.4]
  wire  output_56_17; // @[Switch.scala 41:38:@35063.4]
  wire  _T_73906; // @[Switch.scala 41:52:@35065.4]
  wire  output_56_18; // @[Switch.scala 41:38:@35066.4]
  wire  _T_73909; // @[Switch.scala 41:52:@35068.4]
  wire  output_56_19; // @[Switch.scala 41:38:@35069.4]
  wire  _T_73912; // @[Switch.scala 41:52:@35071.4]
  wire  output_56_20; // @[Switch.scala 41:38:@35072.4]
  wire  _T_73915; // @[Switch.scala 41:52:@35074.4]
  wire  output_56_21; // @[Switch.scala 41:38:@35075.4]
  wire  _T_73918; // @[Switch.scala 41:52:@35077.4]
  wire  output_56_22; // @[Switch.scala 41:38:@35078.4]
  wire  _T_73921; // @[Switch.scala 41:52:@35080.4]
  wire  output_56_23; // @[Switch.scala 41:38:@35081.4]
  wire  _T_73924; // @[Switch.scala 41:52:@35083.4]
  wire  output_56_24; // @[Switch.scala 41:38:@35084.4]
  wire  _T_73927; // @[Switch.scala 41:52:@35086.4]
  wire  output_56_25; // @[Switch.scala 41:38:@35087.4]
  wire  _T_73930; // @[Switch.scala 41:52:@35089.4]
  wire  output_56_26; // @[Switch.scala 41:38:@35090.4]
  wire  _T_73933; // @[Switch.scala 41:52:@35092.4]
  wire  output_56_27; // @[Switch.scala 41:38:@35093.4]
  wire  _T_73936; // @[Switch.scala 41:52:@35095.4]
  wire  output_56_28; // @[Switch.scala 41:38:@35096.4]
  wire  _T_73939; // @[Switch.scala 41:52:@35098.4]
  wire  output_56_29; // @[Switch.scala 41:38:@35099.4]
  wire  _T_73942; // @[Switch.scala 41:52:@35101.4]
  wire  output_56_30; // @[Switch.scala 41:38:@35102.4]
  wire  _T_73945; // @[Switch.scala 41:52:@35104.4]
  wire  output_56_31; // @[Switch.scala 41:38:@35105.4]
  wire  _T_73948; // @[Switch.scala 41:52:@35107.4]
  wire  output_56_32; // @[Switch.scala 41:38:@35108.4]
  wire  _T_73951; // @[Switch.scala 41:52:@35110.4]
  wire  output_56_33; // @[Switch.scala 41:38:@35111.4]
  wire  _T_73954; // @[Switch.scala 41:52:@35113.4]
  wire  output_56_34; // @[Switch.scala 41:38:@35114.4]
  wire  _T_73957; // @[Switch.scala 41:52:@35116.4]
  wire  output_56_35; // @[Switch.scala 41:38:@35117.4]
  wire  _T_73960; // @[Switch.scala 41:52:@35119.4]
  wire  output_56_36; // @[Switch.scala 41:38:@35120.4]
  wire  _T_73963; // @[Switch.scala 41:52:@35122.4]
  wire  output_56_37; // @[Switch.scala 41:38:@35123.4]
  wire  _T_73966; // @[Switch.scala 41:52:@35125.4]
  wire  output_56_38; // @[Switch.scala 41:38:@35126.4]
  wire  _T_73969; // @[Switch.scala 41:52:@35128.4]
  wire  output_56_39; // @[Switch.scala 41:38:@35129.4]
  wire  _T_73972; // @[Switch.scala 41:52:@35131.4]
  wire  output_56_40; // @[Switch.scala 41:38:@35132.4]
  wire  _T_73975; // @[Switch.scala 41:52:@35134.4]
  wire  output_56_41; // @[Switch.scala 41:38:@35135.4]
  wire  _T_73978; // @[Switch.scala 41:52:@35137.4]
  wire  output_56_42; // @[Switch.scala 41:38:@35138.4]
  wire  _T_73981; // @[Switch.scala 41:52:@35140.4]
  wire  output_56_43; // @[Switch.scala 41:38:@35141.4]
  wire  _T_73984; // @[Switch.scala 41:52:@35143.4]
  wire  output_56_44; // @[Switch.scala 41:38:@35144.4]
  wire  _T_73987; // @[Switch.scala 41:52:@35146.4]
  wire  output_56_45; // @[Switch.scala 41:38:@35147.4]
  wire  _T_73990; // @[Switch.scala 41:52:@35149.4]
  wire  output_56_46; // @[Switch.scala 41:38:@35150.4]
  wire  _T_73993; // @[Switch.scala 41:52:@35152.4]
  wire  output_56_47; // @[Switch.scala 41:38:@35153.4]
  wire  _T_73996; // @[Switch.scala 41:52:@35155.4]
  wire  output_56_48; // @[Switch.scala 41:38:@35156.4]
  wire  _T_73999; // @[Switch.scala 41:52:@35158.4]
  wire  output_56_49; // @[Switch.scala 41:38:@35159.4]
  wire  _T_74002; // @[Switch.scala 41:52:@35161.4]
  wire  output_56_50; // @[Switch.scala 41:38:@35162.4]
  wire  _T_74005; // @[Switch.scala 41:52:@35164.4]
  wire  output_56_51; // @[Switch.scala 41:38:@35165.4]
  wire  _T_74008; // @[Switch.scala 41:52:@35167.4]
  wire  output_56_52; // @[Switch.scala 41:38:@35168.4]
  wire  _T_74011; // @[Switch.scala 41:52:@35170.4]
  wire  output_56_53; // @[Switch.scala 41:38:@35171.4]
  wire  _T_74014; // @[Switch.scala 41:52:@35173.4]
  wire  output_56_54; // @[Switch.scala 41:38:@35174.4]
  wire  _T_74017; // @[Switch.scala 41:52:@35176.4]
  wire  output_56_55; // @[Switch.scala 41:38:@35177.4]
  wire  _T_74020; // @[Switch.scala 41:52:@35179.4]
  wire  output_56_56; // @[Switch.scala 41:38:@35180.4]
  wire  _T_74023; // @[Switch.scala 41:52:@35182.4]
  wire  output_56_57; // @[Switch.scala 41:38:@35183.4]
  wire  _T_74026; // @[Switch.scala 41:52:@35185.4]
  wire  output_56_58; // @[Switch.scala 41:38:@35186.4]
  wire  _T_74029; // @[Switch.scala 41:52:@35188.4]
  wire  output_56_59; // @[Switch.scala 41:38:@35189.4]
  wire  _T_74032; // @[Switch.scala 41:52:@35191.4]
  wire  output_56_60; // @[Switch.scala 41:38:@35192.4]
  wire  _T_74035; // @[Switch.scala 41:52:@35194.4]
  wire  output_56_61; // @[Switch.scala 41:38:@35195.4]
  wire  _T_74038; // @[Switch.scala 41:52:@35197.4]
  wire  output_56_62; // @[Switch.scala 41:38:@35198.4]
  wire  _T_74041; // @[Switch.scala 41:52:@35200.4]
  wire  output_56_63; // @[Switch.scala 41:38:@35201.4]
  wire [7:0] _T_74049; // @[Switch.scala 43:31:@35209.4]
  wire [15:0] _T_74057; // @[Switch.scala 43:31:@35217.4]
  wire [7:0] _T_74064; // @[Switch.scala 43:31:@35224.4]
  wire [31:0] _T_74073; // @[Switch.scala 43:31:@35233.4]
  wire [7:0] _T_74080; // @[Switch.scala 43:31:@35240.4]
  wire [15:0] _T_74088; // @[Switch.scala 43:31:@35248.4]
  wire [7:0] _T_74095; // @[Switch.scala 43:31:@35255.4]
  wire [31:0] _T_74104; // @[Switch.scala 43:31:@35264.4]
  wire [63:0] _T_74105; // @[Switch.scala 43:31:@35265.4]
  wire  _T_74109; // @[Switch.scala 41:52:@35268.4]
  wire  output_57_0; // @[Switch.scala 41:38:@35269.4]
  wire  _T_74112; // @[Switch.scala 41:52:@35271.4]
  wire  output_57_1; // @[Switch.scala 41:38:@35272.4]
  wire  _T_74115; // @[Switch.scala 41:52:@35274.4]
  wire  output_57_2; // @[Switch.scala 41:38:@35275.4]
  wire  _T_74118; // @[Switch.scala 41:52:@35277.4]
  wire  output_57_3; // @[Switch.scala 41:38:@35278.4]
  wire  _T_74121; // @[Switch.scala 41:52:@35280.4]
  wire  output_57_4; // @[Switch.scala 41:38:@35281.4]
  wire  _T_74124; // @[Switch.scala 41:52:@35283.4]
  wire  output_57_5; // @[Switch.scala 41:38:@35284.4]
  wire  _T_74127; // @[Switch.scala 41:52:@35286.4]
  wire  output_57_6; // @[Switch.scala 41:38:@35287.4]
  wire  _T_74130; // @[Switch.scala 41:52:@35289.4]
  wire  output_57_7; // @[Switch.scala 41:38:@35290.4]
  wire  _T_74133; // @[Switch.scala 41:52:@35292.4]
  wire  output_57_8; // @[Switch.scala 41:38:@35293.4]
  wire  _T_74136; // @[Switch.scala 41:52:@35295.4]
  wire  output_57_9; // @[Switch.scala 41:38:@35296.4]
  wire  _T_74139; // @[Switch.scala 41:52:@35298.4]
  wire  output_57_10; // @[Switch.scala 41:38:@35299.4]
  wire  _T_74142; // @[Switch.scala 41:52:@35301.4]
  wire  output_57_11; // @[Switch.scala 41:38:@35302.4]
  wire  _T_74145; // @[Switch.scala 41:52:@35304.4]
  wire  output_57_12; // @[Switch.scala 41:38:@35305.4]
  wire  _T_74148; // @[Switch.scala 41:52:@35307.4]
  wire  output_57_13; // @[Switch.scala 41:38:@35308.4]
  wire  _T_74151; // @[Switch.scala 41:52:@35310.4]
  wire  output_57_14; // @[Switch.scala 41:38:@35311.4]
  wire  _T_74154; // @[Switch.scala 41:52:@35313.4]
  wire  output_57_15; // @[Switch.scala 41:38:@35314.4]
  wire  _T_74157; // @[Switch.scala 41:52:@35316.4]
  wire  output_57_16; // @[Switch.scala 41:38:@35317.4]
  wire  _T_74160; // @[Switch.scala 41:52:@35319.4]
  wire  output_57_17; // @[Switch.scala 41:38:@35320.4]
  wire  _T_74163; // @[Switch.scala 41:52:@35322.4]
  wire  output_57_18; // @[Switch.scala 41:38:@35323.4]
  wire  _T_74166; // @[Switch.scala 41:52:@35325.4]
  wire  output_57_19; // @[Switch.scala 41:38:@35326.4]
  wire  _T_74169; // @[Switch.scala 41:52:@35328.4]
  wire  output_57_20; // @[Switch.scala 41:38:@35329.4]
  wire  _T_74172; // @[Switch.scala 41:52:@35331.4]
  wire  output_57_21; // @[Switch.scala 41:38:@35332.4]
  wire  _T_74175; // @[Switch.scala 41:52:@35334.4]
  wire  output_57_22; // @[Switch.scala 41:38:@35335.4]
  wire  _T_74178; // @[Switch.scala 41:52:@35337.4]
  wire  output_57_23; // @[Switch.scala 41:38:@35338.4]
  wire  _T_74181; // @[Switch.scala 41:52:@35340.4]
  wire  output_57_24; // @[Switch.scala 41:38:@35341.4]
  wire  _T_74184; // @[Switch.scala 41:52:@35343.4]
  wire  output_57_25; // @[Switch.scala 41:38:@35344.4]
  wire  _T_74187; // @[Switch.scala 41:52:@35346.4]
  wire  output_57_26; // @[Switch.scala 41:38:@35347.4]
  wire  _T_74190; // @[Switch.scala 41:52:@35349.4]
  wire  output_57_27; // @[Switch.scala 41:38:@35350.4]
  wire  _T_74193; // @[Switch.scala 41:52:@35352.4]
  wire  output_57_28; // @[Switch.scala 41:38:@35353.4]
  wire  _T_74196; // @[Switch.scala 41:52:@35355.4]
  wire  output_57_29; // @[Switch.scala 41:38:@35356.4]
  wire  _T_74199; // @[Switch.scala 41:52:@35358.4]
  wire  output_57_30; // @[Switch.scala 41:38:@35359.4]
  wire  _T_74202; // @[Switch.scala 41:52:@35361.4]
  wire  output_57_31; // @[Switch.scala 41:38:@35362.4]
  wire  _T_74205; // @[Switch.scala 41:52:@35364.4]
  wire  output_57_32; // @[Switch.scala 41:38:@35365.4]
  wire  _T_74208; // @[Switch.scala 41:52:@35367.4]
  wire  output_57_33; // @[Switch.scala 41:38:@35368.4]
  wire  _T_74211; // @[Switch.scala 41:52:@35370.4]
  wire  output_57_34; // @[Switch.scala 41:38:@35371.4]
  wire  _T_74214; // @[Switch.scala 41:52:@35373.4]
  wire  output_57_35; // @[Switch.scala 41:38:@35374.4]
  wire  _T_74217; // @[Switch.scala 41:52:@35376.4]
  wire  output_57_36; // @[Switch.scala 41:38:@35377.4]
  wire  _T_74220; // @[Switch.scala 41:52:@35379.4]
  wire  output_57_37; // @[Switch.scala 41:38:@35380.4]
  wire  _T_74223; // @[Switch.scala 41:52:@35382.4]
  wire  output_57_38; // @[Switch.scala 41:38:@35383.4]
  wire  _T_74226; // @[Switch.scala 41:52:@35385.4]
  wire  output_57_39; // @[Switch.scala 41:38:@35386.4]
  wire  _T_74229; // @[Switch.scala 41:52:@35388.4]
  wire  output_57_40; // @[Switch.scala 41:38:@35389.4]
  wire  _T_74232; // @[Switch.scala 41:52:@35391.4]
  wire  output_57_41; // @[Switch.scala 41:38:@35392.4]
  wire  _T_74235; // @[Switch.scala 41:52:@35394.4]
  wire  output_57_42; // @[Switch.scala 41:38:@35395.4]
  wire  _T_74238; // @[Switch.scala 41:52:@35397.4]
  wire  output_57_43; // @[Switch.scala 41:38:@35398.4]
  wire  _T_74241; // @[Switch.scala 41:52:@35400.4]
  wire  output_57_44; // @[Switch.scala 41:38:@35401.4]
  wire  _T_74244; // @[Switch.scala 41:52:@35403.4]
  wire  output_57_45; // @[Switch.scala 41:38:@35404.4]
  wire  _T_74247; // @[Switch.scala 41:52:@35406.4]
  wire  output_57_46; // @[Switch.scala 41:38:@35407.4]
  wire  _T_74250; // @[Switch.scala 41:52:@35409.4]
  wire  output_57_47; // @[Switch.scala 41:38:@35410.4]
  wire  _T_74253; // @[Switch.scala 41:52:@35412.4]
  wire  output_57_48; // @[Switch.scala 41:38:@35413.4]
  wire  _T_74256; // @[Switch.scala 41:52:@35415.4]
  wire  output_57_49; // @[Switch.scala 41:38:@35416.4]
  wire  _T_74259; // @[Switch.scala 41:52:@35418.4]
  wire  output_57_50; // @[Switch.scala 41:38:@35419.4]
  wire  _T_74262; // @[Switch.scala 41:52:@35421.4]
  wire  output_57_51; // @[Switch.scala 41:38:@35422.4]
  wire  _T_74265; // @[Switch.scala 41:52:@35424.4]
  wire  output_57_52; // @[Switch.scala 41:38:@35425.4]
  wire  _T_74268; // @[Switch.scala 41:52:@35427.4]
  wire  output_57_53; // @[Switch.scala 41:38:@35428.4]
  wire  _T_74271; // @[Switch.scala 41:52:@35430.4]
  wire  output_57_54; // @[Switch.scala 41:38:@35431.4]
  wire  _T_74274; // @[Switch.scala 41:52:@35433.4]
  wire  output_57_55; // @[Switch.scala 41:38:@35434.4]
  wire  _T_74277; // @[Switch.scala 41:52:@35436.4]
  wire  output_57_56; // @[Switch.scala 41:38:@35437.4]
  wire  _T_74280; // @[Switch.scala 41:52:@35439.4]
  wire  output_57_57; // @[Switch.scala 41:38:@35440.4]
  wire  _T_74283; // @[Switch.scala 41:52:@35442.4]
  wire  output_57_58; // @[Switch.scala 41:38:@35443.4]
  wire  _T_74286; // @[Switch.scala 41:52:@35445.4]
  wire  output_57_59; // @[Switch.scala 41:38:@35446.4]
  wire  _T_74289; // @[Switch.scala 41:52:@35448.4]
  wire  output_57_60; // @[Switch.scala 41:38:@35449.4]
  wire  _T_74292; // @[Switch.scala 41:52:@35451.4]
  wire  output_57_61; // @[Switch.scala 41:38:@35452.4]
  wire  _T_74295; // @[Switch.scala 41:52:@35454.4]
  wire  output_57_62; // @[Switch.scala 41:38:@35455.4]
  wire  _T_74298; // @[Switch.scala 41:52:@35457.4]
  wire  output_57_63; // @[Switch.scala 41:38:@35458.4]
  wire [7:0] _T_74306; // @[Switch.scala 43:31:@35466.4]
  wire [15:0] _T_74314; // @[Switch.scala 43:31:@35474.4]
  wire [7:0] _T_74321; // @[Switch.scala 43:31:@35481.4]
  wire [31:0] _T_74330; // @[Switch.scala 43:31:@35490.4]
  wire [7:0] _T_74337; // @[Switch.scala 43:31:@35497.4]
  wire [15:0] _T_74345; // @[Switch.scala 43:31:@35505.4]
  wire [7:0] _T_74352; // @[Switch.scala 43:31:@35512.4]
  wire [31:0] _T_74361; // @[Switch.scala 43:31:@35521.4]
  wire [63:0] _T_74362; // @[Switch.scala 43:31:@35522.4]
  wire  _T_74366; // @[Switch.scala 41:52:@35525.4]
  wire  output_58_0; // @[Switch.scala 41:38:@35526.4]
  wire  _T_74369; // @[Switch.scala 41:52:@35528.4]
  wire  output_58_1; // @[Switch.scala 41:38:@35529.4]
  wire  _T_74372; // @[Switch.scala 41:52:@35531.4]
  wire  output_58_2; // @[Switch.scala 41:38:@35532.4]
  wire  _T_74375; // @[Switch.scala 41:52:@35534.4]
  wire  output_58_3; // @[Switch.scala 41:38:@35535.4]
  wire  _T_74378; // @[Switch.scala 41:52:@35537.4]
  wire  output_58_4; // @[Switch.scala 41:38:@35538.4]
  wire  _T_74381; // @[Switch.scala 41:52:@35540.4]
  wire  output_58_5; // @[Switch.scala 41:38:@35541.4]
  wire  _T_74384; // @[Switch.scala 41:52:@35543.4]
  wire  output_58_6; // @[Switch.scala 41:38:@35544.4]
  wire  _T_74387; // @[Switch.scala 41:52:@35546.4]
  wire  output_58_7; // @[Switch.scala 41:38:@35547.4]
  wire  _T_74390; // @[Switch.scala 41:52:@35549.4]
  wire  output_58_8; // @[Switch.scala 41:38:@35550.4]
  wire  _T_74393; // @[Switch.scala 41:52:@35552.4]
  wire  output_58_9; // @[Switch.scala 41:38:@35553.4]
  wire  _T_74396; // @[Switch.scala 41:52:@35555.4]
  wire  output_58_10; // @[Switch.scala 41:38:@35556.4]
  wire  _T_74399; // @[Switch.scala 41:52:@35558.4]
  wire  output_58_11; // @[Switch.scala 41:38:@35559.4]
  wire  _T_74402; // @[Switch.scala 41:52:@35561.4]
  wire  output_58_12; // @[Switch.scala 41:38:@35562.4]
  wire  _T_74405; // @[Switch.scala 41:52:@35564.4]
  wire  output_58_13; // @[Switch.scala 41:38:@35565.4]
  wire  _T_74408; // @[Switch.scala 41:52:@35567.4]
  wire  output_58_14; // @[Switch.scala 41:38:@35568.4]
  wire  _T_74411; // @[Switch.scala 41:52:@35570.4]
  wire  output_58_15; // @[Switch.scala 41:38:@35571.4]
  wire  _T_74414; // @[Switch.scala 41:52:@35573.4]
  wire  output_58_16; // @[Switch.scala 41:38:@35574.4]
  wire  _T_74417; // @[Switch.scala 41:52:@35576.4]
  wire  output_58_17; // @[Switch.scala 41:38:@35577.4]
  wire  _T_74420; // @[Switch.scala 41:52:@35579.4]
  wire  output_58_18; // @[Switch.scala 41:38:@35580.4]
  wire  _T_74423; // @[Switch.scala 41:52:@35582.4]
  wire  output_58_19; // @[Switch.scala 41:38:@35583.4]
  wire  _T_74426; // @[Switch.scala 41:52:@35585.4]
  wire  output_58_20; // @[Switch.scala 41:38:@35586.4]
  wire  _T_74429; // @[Switch.scala 41:52:@35588.4]
  wire  output_58_21; // @[Switch.scala 41:38:@35589.4]
  wire  _T_74432; // @[Switch.scala 41:52:@35591.4]
  wire  output_58_22; // @[Switch.scala 41:38:@35592.4]
  wire  _T_74435; // @[Switch.scala 41:52:@35594.4]
  wire  output_58_23; // @[Switch.scala 41:38:@35595.4]
  wire  _T_74438; // @[Switch.scala 41:52:@35597.4]
  wire  output_58_24; // @[Switch.scala 41:38:@35598.4]
  wire  _T_74441; // @[Switch.scala 41:52:@35600.4]
  wire  output_58_25; // @[Switch.scala 41:38:@35601.4]
  wire  _T_74444; // @[Switch.scala 41:52:@35603.4]
  wire  output_58_26; // @[Switch.scala 41:38:@35604.4]
  wire  _T_74447; // @[Switch.scala 41:52:@35606.4]
  wire  output_58_27; // @[Switch.scala 41:38:@35607.4]
  wire  _T_74450; // @[Switch.scala 41:52:@35609.4]
  wire  output_58_28; // @[Switch.scala 41:38:@35610.4]
  wire  _T_74453; // @[Switch.scala 41:52:@35612.4]
  wire  output_58_29; // @[Switch.scala 41:38:@35613.4]
  wire  _T_74456; // @[Switch.scala 41:52:@35615.4]
  wire  output_58_30; // @[Switch.scala 41:38:@35616.4]
  wire  _T_74459; // @[Switch.scala 41:52:@35618.4]
  wire  output_58_31; // @[Switch.scala 41:38:@35619.4]
  wire  _T_74462; // @[Switch.scala 41:52:@35621.4]
  wire  output_58_32; // @[Switch.scala 41:38:@35622.4]
  wire  _T_74465; // @[Switch.scala 41:52:@35624.4]
  wire  output_58_33; // @[Switch.scala 41:38:@35625.4]
  wire  _T_74468; // @[Switch.scala 41:52:@35627.4]
  wire  output_58_34; // @[Switch.scala 41:38:@35628.4]
  wire  _T_74471; // @[Switch.scala 41:52:@35630.4]
  wire  output_58_35; // @[Switch.scala 41:38:@35631.4]
  wire  _T_74474; // @[Switch.scala 41:52:@35633.4]
  wire  output_58_36; // @[Switch.scala 41:38:@35634.4]
  wire  _T_74477; // @[Switch.scala 41:52:@35636.4]
  wire  output_58_37; // @[Switch.scala 41:38:@35637.4]
  wire  _T_74480; // @[Switch.scala 41:52:@35639.4]
  wire  output_58_38; // @[Switch.scala 41:38:@35640.4]
  wire  _T_74483; // @[Switch.scala 41:52:@35642.4]
  wire  output_58_39; // @[Switch.scala 41:38:@35643.4]
  wire  _T_74486; // @[Switch.scala 41:52:@35645.4]
  wire  output_58_40; // @[Switch.scala 41:38:@35646.4]
  wire  _T_74489; // @[Switch.scala 41:52:@35648.4]
  wire  output_58_41; // @[Switch.scala 41:38:@35649.4]
  wire  _T_74492; // @[Switch.scala 41:52:@35651.4]
  wire  output_58_42; // @[Switch.scala 41:38:@35652.4]
  wire  _T_74495; // @[Switch.scala 41:52:@35654.4]
  wire  output_58_43; // @[Switch.scala 41:38:@35655.4]
  wire  _T_74498; // @[Switch.scala 41:52:@35657.4]
  wire  output_58_44; // @[Switch.scala 41:38:@35658.4]
  wire  _T_74501; // @[Switch.scala 41:52:@35660.4]
  wire  output_58_45; // @[Switch.scala 41:38:@35661.4]
  wire  _T_74504; // @[Switch.scala 41:52:@35663.4]
  wire  output_58_46; // @[Switch.scala 41:38:@35664.4]
  wire  _T_74507; // @[Switch.scala 41:52:@35666.4]
  wire  output_58_47; // @[Switch.scala 41:38:@35667.4]
  wire  _T_74510; // @[Switch.scala 41:52:@35669.4]
  wire  output_58_48; // @[Switch.scala 41:38:@35670.4]
  wire  _T_74513; // @[Switch.scala 41:52:@35672.4]
  wire  output_58_49; // @[Switch.scala 41:38:@35673.4]
  wire  _T_74516; // @[Switch.scala 41:52:@35675.4]
  wire  output_58_50; // @[Switch.scala 41:38:@35676.4]
  wire  _T_74519; // @[Switch.scala 41:52:@35678.4]
  wire  output_58_51; // @[Switch.scala 41:38:@35679.4]
  wire  _T_74522; // @[Switch.scala 41:52:@35681.4]
  wire  output_58_52; // @[Switch.scala 41:38:@35682.4]
  wire  _T_74525; // @[Switch.scala 41:52:@35684.4]
  wire  output_58_53; // @[Switch.scala 41:38:@35685.4]
  wire  _T_74528; // @[Switch.scala 41:52:@35687.4]
  wire  output_58_54; // @[Switch.scala 41:38:@35688.4]
  wire  _T_74531; // @[Switch.scala 41:52:@35690.4]
  wire  output_58_55; // @[Switch.scala 41:38:@35691.4]
  wire  _T_74534; // @[Switch.scala 41:52:@35693.4]
  wire  output_58_56; // @[Switch.scala 41:38:@35694.4]
  wire  _T_74537; // @[Switch.scala 41:52:@35696.4]
  wire  output_58_57; // @[Switch.scala 41:38:@35697.4]
  wire  _T_74540; // @[Switch.scala 41:52:@35699.4]
  wire  output_58_58; // @[Switch.scala 41:38:@35700.4]
  wire  _T_74543; // @[Switch.scala 41:52:@35702.4]
  wire  output_58_59; // @[Switch.scala 41:38:@35703.4]
  wire  _T_74546; // @[Switch.scala 41:52:@35705.4]
  wire  output_58_60; // @[Switch.scala 41:38:@35706.4]
  wire  _T_74549; // @[Switch.scala 41:52:@35708.4]
  wire  output_58_61; // @[Switch.scala 41:38:@35709.4]
  wire  _T_74552; // @[Switch.scala 41:52:@35711.4]
  wire  output_58_62; // @[Switch.scala 41:38:@35712.4]
  wire  _T_74555; // @[Switch.scala 41:52:@35714.4]
  wire  output_58_63; // @[Switch.scala 41:38:@35715.4]
  wire [7:0] _T_74563; // @[Switch.scala 43:31:@35723.4]
  wire [15:0] _T_74571; // @[Switch.scala 43:31:@35731.4]
  wire [7:0] _T_74578; // @[Switch.scala 43:31:@35738.4]
  wire [31:0] _T_74587; // @[Switch.scala 43:31:@35747.4]
  wire [7:0] _T_74594; // @[Switch.scala 43:31:@35754.4]
  wire [15:0] _T_74602; // @[Switch.scala 43:31:@35762.4]
  wire [7:0] _T_74609; // @[Switch.scala 43:31:@35769.4]
  wire [31:0] _T_74618; // @[Switch.scala 43:31:@35778.4]
  wire [63:0] _T_74619; // @[Switch.scala 43:31:@35779.4]
  wire  _T_74623; // @[Switch.scala 41:52:@35782.4]
  wire  output_59_0; // @[Switch.scala 41:38:@35783.4]
  wire  _T_74626; // @[Switch.scala 41:52:@35785.4]
  wire  output_59_1; // @[Switch.scala 41:38:@35786.4]
  wire  _T_74629; // @[Switch.scala 41:52:@35788.4]
  wire  output_59_2; // @[Switch.scala 41:38:@35789.4]
  wire  _T_74632; // @[Switch.scala 41:52:@35791.4]
  wire  output_59_3; // @[Switch.scala 41:38:@35792.4]
  wire  _T_74635; // @[Switch.scala 41:52:@35794.4]
  wire  output_59_4; // @[Switch.scala 41:38:@35795.4]
  wire  _T_74638; // @[Switch.scala 41:52:@35797.4]
  wire  output_59_5; // @[Switch.scala 41:38:@35798.4]
  wire  _T_74641; // @[Switch.scala 41:52:@35800.4]
  wire  output_59_6; // @[Switch.scala 41:38:@35801.4]
  wire  _T_74644; // @[Switch.scala 41:52:@35803.4]
  wire  output_59_7; // @[Switch.scala 41:38:@35804.4]
  wire  _T_74647; // @[Switch.scala 41:52:@35806.4]
  wire  output_59_8; // @[Switch.scala 41:38:@35807.4]
  wire  _T_74650; // @[Switch.scala 41:52:@35809.4]
  wire  output_59_9; // @[Switch.scala 41:38:@35810.4]
  wire  _T_74653; // @[Switch.scala 41:52:@35812.4]
  wire  output_59_10; // @[Switch.scala 41:38:@35813.4]
  wire  _T_74656; // @[Switch.scala 41:52:@35815.4]
  wire  output_59_11; // @[Switch.scala 41:38:@35816.4]
  wire  _T_74659; // @[Switch.scala 41:52:@35818.4]
  wire  output_59_12; // @[Switch.scala 41:38:@35819.4]
  wire  _T_74662; // @[Switch.scala 41:52:@35821.4]
  wire  output_59_13; // @[Switch.scala 41:38:@35822.4]
  wire  _T_74665; // @[Switch.scala 41:52:@35824.4]
  wire  output_59_14; // @[Switch.scala 41:38:@35825.4]
  wire  _T_74668; // @[Switch.scala 41:52:@35827.4]
  wire  output_59_15; // @[Switch.scala 41:38:@35828.4]
  wire  _T_74671; // @[Switch.scala 41:52:@35830.4]
  wire  output_59_16; // @[Switch.scala 41:38:@35831.4]
  wire  _T_74674; // @[Switch.scala 41:52:@35833.4]
  wire  output_59_17; // @[Switch.scala 41:38:@35834.4]
  wire  _T_74677; // @[Switch.scala 41:52:@35836.4]
  wire  output_59_18; // @[Switch.scala 41:38:@35837.4]
  wire  _T_74680; // @[Switch.scala 41:52:@35839.4]
  wire  output_59_19; // @[Switch.scala 41:38:@35840.4]
  wire  _T_74683; // @[Switch.scala 41:52:@35842.4]
  wire  output_59_20; // @[Switch.scala 41:38:@35843.4]
  wire  _T_74686; // @[Switch.scala 41:52:@35845.4]
  wire  output_59_21; // @[Switch.scala 41:38:@35846.4]
  wire  _T_74689; // @[Switch.scala 41:52:@35848.4]
  wire  output_59_22; // @[Switch.scala 41:38:@35849.4]
  wire  _T_74692; // @[Switch.scala 41:52:@35851.4]
  wire  output_59_23; // @[Switch.scala 41:38:@35852.4]
  wire  _T_74695; // @[Switch.scala 41:52:@35854.4]
  wire  output_59_24; // @[Switch.scala 41:38:@35855.4]
  wire  _T_74698; // @[Switch.scala 41:52:@35857.4]
  wire  output_59_25; // @[Switch.scala 41:38:@35858.4]
  wire  _T_74701; // @[Switch.scala 41:52:@35860.4]
  wire  output_59_26; // @[Switch.scala 41:38:@35861.4]
  wire  _T_74704; // @[Switch.scala 41:52:@35863.4]
  wire  output_59_27; // @[Switch.scala 41:38:@35864.4]
  wire  _T_74707; // @[Switch.scala 41:52:@35866.4]
  wire  output_59_28; // @[Switch.scala 41:38:@35867.4]
  wire  _T_74710; // @[Switch.scala 41:52:@35869.4]
  wire  output_59_29; // @[Switch.scala 41:38:@35870.4]
  wire  _T_74713; // @[Switch.scala 41:52:@35872.4]
  wire  output_59_30; // @[Switch.scala 41:38:@35873.4]
  wire  _T_74716; // @[Switch.scala 41:52:@35875.4]
  wire  output_59_31; // @[Switch.scala 41:38:@35876.4]
  wire  _T_74719; // @[Switch.scala 41:52:@35878.4]
  wire  output_59_32; // @[Switch.scala 41:38:@35879.4]
  wire  _T_74722; // @[Switch.scala 41:52:@35881.4]
  wire  output_59_33; // @[Switch.scala 41:38:@35882.4]
  wire  _T_74725; // @[Switch.scala 41:52:@35884.4]
  wire  output_59_34; // @[Switch.scala 41:38:@35885.4]
  wire  _T_74728; // @[Switch.scala 41:52:@35887.4]
  wire  output_59_35; // @[Switch.scala 41:38:@35888.4]
  wire  _T_74731; // @[Switch.scala 41:52:@35890.4]
  wire  output_59_36; // @[Switch.scala 41:38:@35891.4]
  wire  _T_74734; // @[Switch.scala 41:52:@35893.4]
  wire  output_59_37; // @[Switch.scala 41:38:@35894.4]
  wire  _T_74737; // @[Switch.scala 41:52:@35896.4]
  wire  output_59_38; // @[Switch.scala 41:38:@35897.4]
  wire  _T_74740; // @[Switch.scala 41:52:@35899.4]
  wire  output_59_39; // @[Switch.scala 41:38:@35900.4]
  wire  _T_74743; // @[Switch.scala 41:52:@35902.4]
  wire  output_59_40; // @[Switch.scala 41:38:@35903.4]
  wire  _T_74746; // @[Switch.scala 41:52:@35905.4]
  wire  output_59_41; // @[Switch.scala 41:38:@35906.4]
  wire  _T_74749; // @[Switch.scala 41:52:@35908.4]
  wire  output_59_42; // @[Switch.scala 41:38:@35909.4]
  wire  _T_74752; // @[Switch.scala 41:52:@35911.4]
  wire  output_59_43; // @[Switch.scala 41:38:@35912.4]
  wire  _T_74755; // @[Switch.scala 41:52:@35914.4]
  wire  output_59_44; // @[Switch.scala 41:38:@35915.4]
  wire  _T_74758; // @[Switch.scala 41:52:@35917.4]
  wire  output_59_45; // @[Switch.scala 41:38:@35918.4]
  wire  _T_74761; // @[Switch.scala 41:52:@35920.4]
  wire  output_59_46; // @[Switch.scala 41:38:@35921.4]
  wire  _T_74764; // @[Switch.scala 41:52:@35923.4]
  wire  output_59_47; // @[Switch.scala 41:38:@35924.4]
  wire  _T_74767; // @[Switch.scala 41:52:@35926.4]
  wire  output_59_48; // @[Switch.scala 41:38:@35927.4]
  wire  _T_74770; // @[Switch.scala 41:52:@35929.4]
  wire  output_59_49; // @[Switch.scala 41:38:@35930.4]
  wire  _T_74773; // @[Switch.scala 41:52:@35932.4]
  wire  output_59_50; // @[Switch.scala 41:38:@35933.4]
  wire  _T_74776; // @[Switch.scala 41:52:@35935.4]
  wire  output_59_51; // @[Switch.scala 41:38:@35936.4]
  wire  _T_74779; // @[Switch.scala 41:52:@35938.4]
  wire  output_59_52; // @[Switch.scala 41:38:@35939.4]
  wire  _T_74782; // @[Switch.scala 41:52:@35941.4]
  wire  output_59_53; // @[Switch.scala 41:38:@35942.4]
  wire  _T_74785; // @[Switch.scala 41:52:@35944.4]
  wire  output_59_54; // @[Switch.scala 41:38:@35945.4]
  wire  _T_74788; // @[Switch.scala 41:52:@35947.4]
  wire  output_59_55; // @[Switch.scala 41:38:@35948.4]
  wire  _T_74791; // @[Switch.scala 41:52:@35950.4]
  wire  output_59_56; // @[Switch.scala 41:38:@35951.4]
  wire  _T_74794; // @[Switch.scala 41:52:@35953.4]
  wire  output_59_57; // @[Switch.scala 41:38:@35954.4]
  wire  _T_74797; // @[Switch.scala 41:52:@35956.4]
  wire  output_59_58; // @[Switch.scala 41:38:@35957.4]
  wire  _T_74800; // @[Switch.scala 41:52:@35959.4]
  wire  output_59_59; // @[Switch.scala 41:38:@35960.4]
  wire  _T_74803; // @[Switch.scala 41:52:@35962.4]
  wire  output_59_60; // @[Switch.scala 41:38:@35963.4]
  wire  _T_74806; // @[Switch.scala 41:52:@35965.4]
  wire  output_59_61; // @[Switch.scala 41:38:@35966.4]
  wire  _T_74809; // @[Switch.scala 41:52:@35968.4]
  wire  output_59_62; // @[Switch.scala 41:38:@35969.4]
  wire  _T_74812; // @[Switch.scala 41:52:@35971.4]
  wire  output_59_63; // @[Switch.scala 41:38:@35972.4]
  wire [7:0] _T_74820; // @[Switch.scala 43:31:@35980.4]
  wire [15:0] _T_74828; // @[Switch.scala 43:31:@35988.4]
  wire [7:0] _T_74835; // @[Switch.scala 43:31:@35995.4]
  wire [31:0] _T_74844; // @[Switch.scala 43:31:@36004.4]
  wire [7:0] _T_74851; // @[Switch.scala 43:31:@36011.4]
  wire [15:0] _T_74859; // @[Switch.scala 43:31:@36019.4]
  wire [7:0] _T_74866; // @[Switch.scala 43:31:@36026.4]
  wire [31:0] _T_74875; // @[Switch.scala 43:31:@36035.4]
  wire [63:0] _T_74876; // @[Switch.scala 43:31:@36036.4]
  wire  _T_74880; // @[Switch.scala 41:52:@36039.4]
  wire  output_60_0; // @[Switch.scala 41:38:@36040.4]
  wire  _T_74883; // @[Switch.scala 41:52:@36042.4]
  wire  output_60_1; // @[Switch.scala 41:38:@36043.4]
  wire  _T_74886; // @[Switch.scala 41:52:@36045.4]
  wire  output_60_2; // @[Switch.scala 41:38:@36046.4]
  wire  _T_74889; // @[Switch.scala 41:52:@36048.4]
  wire  output_60_3; // @[Switch.scala 41:38:@36049.4]
  wire  _T_74892; // @[Switch.scala 41:52:@36051.4]
  wire  output_60_4; // @[Switch.scala 41:38:@36052.4]
  wire  _T_74895; // @[Switch.scala 41:52:@36054.4]
  wire  output_60_5; // @[Switch.scala 41:38:@36055.4]
  wire  _T_74898; // @[Switch.scala 41:52:@36057.4]
  wire  output_60_6; // @[Switch.scala 41:38:@36058.4]
  wire  _T_74901; // @[Switch.scala 41:52:@36060.4]
  wire  output_60_7; // @[Switch.scala 41:38:@36061.4]
  wire  _T_74904; // @[Switch.scala 41:52:@36063.4]
  wire  output_60_8; // @[Switch.scala 41:38:@36064.4]
  wire  _T_74907; // @[Switch.scala 41:52:@36066.4]
  wire  output_60_9; // @[Switch.scala 41:38:@36067.4]
  wire  _T_74910; // @[Switch.scala 41:52:@36069.4]
  wire  output_60_10; // @[Switch.scala 41:38:@36070.4]
  wire  _T_74913; // @[Switch.scala 41:52:@36072.4]
  wire  output_60_11; // @[Switch.scala 41:38:@36073.4]
  wire  _T_74916; // @[Switch.scala 41:52:@36075.4]
  wire  output_60_12; // @[Switch.scala 41:38:@36076.4]
  wire  _T_74919; // @[Switch.scala 41:52:@36078.4]
  wire  output_60_13; // @[Switch.scala 41:38:@36079.4]
  wire  _T_74922; // @[Switch.scala 41:52:@36081.4]
  wire  output_60_14; // @[Switch.scala 41:38:@36082.4]
  wire  _T_74925; // @[Switch.scala 41:52:@36084.4]
  wire  output_60_15; // @[Switch.scala 41:38:@36085.4]
  wire  _T_74928; // @[Switch.scala 41:52:@36087.4]
  wire  output_60_16; // @[Switch.scala 41:38:@36088.4]
  wire  _T_74931; // @[Switch.scala 41:52:@36090.4]
  wire  output_60_17; // @[Switch.scala 41:38:@36091.4]
  wire  _T_74934; // @[Switch.scala 41:52:@36093.4]
  wire  output_60_18; // @[Switch.scala 41:38:@36094.4]
  wire  _T_74937; // @[Switch.scala 41:52:@36096.4]
  wire  output_60_19; // @[Switch.scala 41:38:@36097.4]
  wire  _T_74940; // @[Switch.scala 41:52:@36099.4]
  wire  output_60_20; // @[Switch.scala 41:38:@36100.4]
  wire  _T_74943; // @[Switch.scala 41:52:@36102.4]
  wire  output_60_21; // @[Switch.scala 41:38:@36103.4]
  wire  _T_74946; // @[Switch.scala 41:52:@36105.4]
  wire  output_60_22; // @[Switch.scala 41:38:@36106.4]
  wire  _T_74949; // @[Switch.scala 41:52:@36108.4]
  wire  output_60_23; // @[Switch.scala 41:38:@36109.4]
  wire  _T_74952; // @[Switch.scala 41:52:@36111.4]
  wire  output_60_24; // @[Switch.scala 41:38:@36112.4]
  wire  _T_74955; // @[Switch.scala 41:52:@36114.4]
  wire  output_60_25; // @[Switch.scala 41:38:@36115.4]
  wire  _T_74958; // @[Switch.scala 41:52:@36117.4]
  wire  output_60_26; // @[Switch.scala 41:38:@36118.4]
  wire  _T_74961; // @[Switch.scala 41:52:@36120.4]
  wire  output_60_27; // @[Switch.scala 41:38:@36121.4]
  wire  _T_74964; // @[Switch.scala 41:52:@36123.4]
  wire  output_60_28; // @[Switch.scala 41:38:@36124.4]
  wire  _T_74967; // @[Switch.scala 41:52:@36126.4]
  wire  output_60_29; // @[Switch.scala 41:38:@36127.4]
  wire  _T_74970; // @[Switch.scala 41:52:@36129.4]
  wire  output_60_30; // @[Switch.scala 41:38:@36130.4]
  wire  _T_74973; // @[Switch.scala 41:52:@36132.4]
  wire  output_60_31; // @[Switch.scala 41:38:@36133.4]
  wire  _T_74976; // @[Switch.scala 41:52:@36135.4]
  wire  output_60_32; // @[Switch.scala 41:38:@36136.4]
  wire  _T_74979; // @[Switch.scala 41:52:@36138.4]
  wire  output_60_33; // @[Switch.scala 41:38:@36139.4]
  wire  _T_74982; // @[Switch.scala 41:52:@36141.4]
  wire  output_60_34; // @[Switch.scala 41:38:@36142.4]
  wire  _T_74985; // @[Switch.scala 41:52:@36144.4]
  wire  output_60_35; // @[Switch.scala 41:38:@36145.4]
  wire  _T_74988; // @[Switch.scala 41:52:@36147.4]
  wire  output_60_36; // @[Switch.scala 41:38:@36148.4]
  wire  _T_74991; // @[Switch.scala 41:52:@36150.4]
  wire  output_60_37; // @[Switch.scala 41:38:@36151.4]
  wire  _T_74994; // @[Switch.scala 41:52:@36153.4]
  wire  output_60_38; // @[Switch.scala 41:38:@36154.4]
  wire  _T_74997; // @[Switch.scala 41:52:@36156.4]
  wire  output_60_39; // @[Switch.scala 41:38:@36157.4]
  wire  _T_75000; // @[Switch.scala 41:52:@36159.4]
  wire  output_60_40; // @[Switch.scala 41:38:@36160.4]
  wire  _T_75003; // @[Switch.scala 41:52:@36162.4]
  wire  output_60_41; // @[Switch.scala 41:38:@36163.4]
  wire  _T_75006; // @[Switch.scala 41:52:@36165.4]
  wire  output_60_42; // @[Switch.scala 41:38:@36166.4]
  wire  _T_75009; // @[Switch.scala 41:52:@36168.4]
  wire  output_60_43; // @[Switch.scala 41:38:@36169.4]
  wire  _T_75012; // @[Switch.scala 41:52:@36171.4]
  wire  output_60_44; // @[Switch.scala 41:38:@36172.4]
  wire  _T_75015; // @[Switch.scala 41:52:@36174.4]
  wire  output_60_45; // @[Switch.scala 41:38:@36175.4]
  wire  _T_75018; // @[Switch.scala 41:52:@36177.4]
  wire  output_60_46; // @[Switch.scala 41:38:@36178.4]
  wire  _T_75021; // @[Switch.scala 41:52:@36180.4]
  wire  output_60_47; // @[Switch.scala 41:38:@36181.4]
  wire  _T_75024; // @[Switch.scala 41:52:@36183.4]
  wire  output_60_48; // @[Switch.scala 41:38:@36184.4]
  wire  _T_75027; // @[Switch.scala 41:52:@36186.4]
  wire  output_60_49; // @[Switch.scala 41:38:@36187.4]
  wire  _T_75030; // @[Switch.scala 41:52:@36189.4]
  wire  output_60_50; // @[Switch.scala 41:38:@36190.4]
  wire  _T_75033; // @[Switch.scala 41:52:@36192.4]
  wire  output_60_51; // @[Switch.scala 41:38:@36193.4]
  wire  _T_75036; // @[Switch.scala 41:52:@36195.4]
  wire  output_60_52; // @[Switch.scala 41:38:@36196.4]
  wire  _T_75039; // @[Switch.scala 41:52:@36198.4]
  wire  output_60_53; // @[Switch.scala 41:38:@36199.4]
  wire  _T_75042; // @[Switch.scala 41:52:@36201.4]
  wire  output_60_54; // @[Switch.scala 41:38:@36202.4]
  wire  _T_75045; // @[Switch.scala 41:52:@36204.4]
  wire  output_60_55; // @[Switch.scala 41:38:@36205.4]
  wire  _T_75048; // @[Switch.scala 41:52:@36207.4]
  wire  output_60_56; // @[Switch.scala 41:38:@36208.4]
  wire  _T_75051; // @[Switch.scala 41:52:@36210.4]
  wire  output_60_57; // @[Switch.scala 41:38:@36211.4]
  wire  _T_75054; // @[Switch.scala 41:52:@36213.4]
  wire  output_60_58; // @[Switch.scala 41:38:@36214.4]
  wire  _T_75057; // @[Switch.scala 41:52:@36216.4]
  wire  output_60_59; // @[Switch.scala 41:38:@36217.4]
  wire  _T_75060; // @[Switch.scala 41:52:@36219.4]
  wire  output_60_60; // @[Switch.scala 41:38:@36220.4]
  wire  _T_75063; // @[Switch.scala 41:52:@36222.4]
  wire  output_60_61; // @[Switch.scala 41:38:@36223.4]
  wire  _T_75066; // @[Switch.scala 41:52:@36225.4]
  wire  output_60_62; // @[Switch.scala 41:38:@36226.4]
  wire  _T_75069; // @[Switch.scala 41:52:@36228.4]
  wire  output_60_63; // @[Switch.scala 41:38:@36229.4]
  wire [7:0] _T_75077; // @[Switch.scala 43:31:@36237.4]
  wire [15:0] _T_75085; // @[Switch.scala 43:31:@36245.4]
  wire [7:0] _T_75092; // @[Switch.scala 43:31:@36252.4]
  wire [31:0] _T_75101; // @[Switch.scala 43:31:@36261.4]
  wire [7:0] _T_75108; // @[Switch.scala 43:31:@36268.4]
  wire [15:0] _T_75116; // @[Switch.scala 43:31:@36276.4]
  wire [7:0] _T_75123; // @[Switch.scala 43:31:@36283.4]
  wire [31:0] _T_75132; // @[Switch.scala 43:31:@36292.4]
  wire [63:0] _T_75133; // @[Switch.scala 43:31:@36293.4]
  wire  _T_75137; // @[Switch.scala 41:52:@36296.4]
  wire  output_61_0; // @[Switch.scala 41:38:@36297.4]
  wire  _T_75140; // @[Switch.scala 41:52:@36299.4]
  wire  output_61_1; // @[Switch.scala 41:38:@36300.4]
  wire  _T_75143; // @[Switch.scala 41:52:@36302.4]
  wire  output_61_2; // @[Switch.scala 41:38:@36303.4]
  wire  _T_75146; // @[Switch.scala 41:52:@36305.4]
  wire  output_61_3; // @[Switch.scala 41:38:@36306.4]
  wire  _T_75149; // @[Switch.scala 41:52:@36308.4]
  wire  output_61_4; // @[Switch.scala 41:38:@36309.4]
  wire  _T_75152; // @[Switch.scala 41:52:@36311.4]
  wire  output_61_5; // @[Switch.scala 41:38:@36312.4]
  wire  _T_75155; // @[Switch.scala 41:52:@36314.4]
  wire  output_61_6; // @[Switch.scala 41:38:@36315.4]
  wire  _T_75158; // @[Switch.scala 41:52:@36317.4]
  wire  output_61_7; // @[Switch.scala 41:38:@36318.4]
  wire  _T_75161; // @[Switch.scala 41:52:@36320.4]
  wire  output_61_8; // @[Switch.scala 41:38:@36321.4]
  wire  _T_75164; // @[Switch.scala 41:52:@36323.4]
  wire  output_61_9; // @[Switch.scala 41:38:@36324.4]
  wire  _T_75167; // @[Switch.scala 41:52:@36326.4]
  wire  output_61_10; // @[Switch.scala 41:38:@36327.4]
  wire  _T_75170; // @[Switch.scala 41:52:@36329.4]
  wire  output_61_11; // @[Switch.scala 41:38:@36330.4]
  wire  _T_75173; // @[Switch.scala 41:52:@36332.4]
  wire  output_61_12; // @[Switch.scala 41:38:@36333.4]
  wire  _T_75176; // @[Switch.scala 41:52:@36335.4]
  wire  output_61_13; // @[Switch.scala 41:38:@36336.4]
  wire  _T_75179; // @[Switch.scala 41:52:@36338.4]
  wire  output_61_14; // @[Switch.scala 41:38:@36339.4]
  wire  _T_75182; // @[Switch.scala 41:52:@36341.4]
  wire  output_61_15; // @[Switch.scala 41:38:@36342.4]
  wire  _T_75185; // @[Switch.scala 41:52:@36344.4]
  wire  output_61_16; // @[Switch.scala 41:38:@36345.4]
  wire  _T_75188; // @[Switch.scala 41:52:@36347.4]
  wire  output_61_17; // @[Switch.scala 41:38:@36348.4]
  wire  _T_75191; // @[Switch.scala 41:52:@36350.4]
  wire  output_61_18; // @[Switch.scala 41:38:@36351.4]
  wire  _T_75194; // @[Switch.scala 41:52:@36353.4]
  wire  output_61_19; // @[Switch.scala 41:38:@36354.4]
  wire  _T_75197; // @[Switch.scala 41:52:@36356.4]
  wire  output_61_20; // @[Switch.scala 41:38:@36357.4]
  wire  _T_75200; // @[Switch.scala 41:52:@36359.4]
  wire  output_61_21; // @[Switch.scala 41:38:@36360.4]
  wire  _T_75203; // @[Switch.scala 41:52:@36362.4]
  wire  output_61_22; // @[Switch.scala 41:38:@36363.4]
  wire  _T_75206; // @[Switch.scala 41:52:@36365.4]
  wire  output_61_23; // @[Switch.scala 41:38:@36366.4]
  wire  _T_75209; // @[Switch.scala 41:52:@36368.4]
  wire  output_61_24; // @[Switch.scala 41:38:@36369.4]
  wire  _T_75212; // @[Switch.scala 41:52:@36371.4]
  wire  output_61_25; // @[Switch.scala 41:38:@36372.4]
  wire  _T_75215; // @[Switch.scala 41:52:@36374.4]
  wire  output_61_26; // @[Switch.scala 41:38:@36375.4]
  wire  _T_75218; // @[Switch.scala 41:52:@36377.4]
  wire  output_61_27; // @[Switch.scala 41:38:@36378.4]
  wire  _T_75221; // @[Switch.scala 41:52:@36380.4]
  wire  output_61_28; // @[Switch.scala 41:38:@36381.4]
  wire  _T_75224; // @[Switch.scala 41:52:@36383.4]
  wire  output_61_29; // @[Switch.scala 41:38:@36384.4]
  wire  _T_75227; // @[Switch.scala 41:52:@36386.4]
  wire  output_61_30; // @[Switch.scala 41:38:@36387.4]
  wire  _T_75230; // @[Switch.scala 41:52:@36389.4]
  wire  output_61_31; // @[Switch.scala 41:38:@36390.4]
  wire  _T_75233; // @[Switch.scala 41:52:@36392.4]
  wire  output_61_32; // @[Switch.scala 41:38:@36393.4]
  wire  _T_75236; // @[Switch.scala 41:52:@36395.4]
  wire  output_61_33; // @[Switch.scala 41:38:@36396.4]
  wire  _T_75239; // @[Switch.scala 41:52:@36398.4]
  wire  output_61_34; // @[Switch.scala 41:38:@36399.4]
  wire  _T_75242; // @[Switch.scala 41:52:@36401.4]
  wire  output_61_35; // @[Switch.scala 41:38:@36402.4]
  wire  _T_75245; // @[Switch.scala 41:52:@36404.4]
  wire  output_61_36; // @[Switch.scala 41:38:@36405.4]
  wire  _T_75248; // @[Switch.scala 41:52:@36407.4]
  wire  output_61_37; // @[Switch.scala 41:38:@36408.4]
  wire  _T_75251; // @[Switch.scala 41:52:@36410.4]
  wire  output_61_38; // @[Switch.scala 41:38:@36411.4]
  wire  _T_75254; // @[Switch.scala 41:52:@36413.4]
  wire  output_61_39; // @[Switch.scala 41:38:@36414.4]
  wire  _T_75257; // @[Switch.scala 41:52:@36416.4]
  wire  output_61_40; // @[Switch.scala 41:38:@36417.4]
  wire  _T_75260; // @[Switch.scala 41:52:@36419.4]
  wire  output_61_41; // @[Switch.scala 41:38:@36420.4]
  wire  _T_75263; // @[Switch.scala 41:52:@36422.4]
  wire  output_61_42; // @[Switch.scala 41:38:@36423.4]
  wire  _T_75266; // @[Switch.scala 41:52:@36425.4]
  wire  output_61_43; // @[Switch.scala 41:38:@36426.4]
  wire  _T_75269; // @[Switch.scala 41:52:@36428.4]
  wire  output_61_44; // @[Switch.scala 41:38:@36429.4]
  wire  _T_75272; // @[Switch.scala 41:52:@36431.4]
  wire  output_61_45; // @[Switch.scala 41:38:@36432.4]
  wire  _T_75275; // @[Switch.scala 41:52:@36434.4]
  wire  output_61_46; // @[Switch.scala 41:38:@36435.4]
  wire  _T_75278; // @[Switch.scala 41:52:@36437.4]
  wire  output_61_47; // @[Switch.scala 41:38:@36438.4]
  wire  _T_75281; // @[Switch.scala 41:52:@36440.4]
  wire  output_61_48; // @[Switch.scala 41:38:@36441.4]
  wire  _T_75284; // @[Switch.scala 41:52:@36443.4]
  wire  output_61_49; // @[Switch.scala 41:38:@36444.4]
  wire  _T_75287; // @[Switch.scala 41:52:@36446.4]
  wire  output_61_50; // @[Switch.scala 41:38:@36447.4]
  wire  _T_75290; // @[Switch.scala 41:52:@36449.4]
  wire  output_61_51; // @[Switch.scala 41:38:@36450.4]
  wire  _T_75293; // @[Switch.scala 41:52:@36452.4]
  wire  output_61_52; // @[Switch.scala 41:38:@36453.4]
  wire  _T_75296; // @[Switch.scala 41:52:@36455.4]
  wire  output_61_53; // @[Switch.scala 41:38:@36456.4]
  wire  _T_75299; // @[Switch.scala 41:52:@36458.4]
  wire  output_61_54; // @[Switch.scala 41:38:@36459.4]
  wire  _T_75302; // @[Switch.scala 41:52:@36461.4]
  wire  output_61_55; // @[Switch.scala 41:38:@36462.4]
  wire  _T_75305; // @[Switch.scala 41:52:@36464.4]
  wire  output_61_56; // @[Switch.scala 41:38:@36465.4]
  wire  _T_75308; // @[Switch.scala 41:52:@36467.4]
  wire  output_61_57; // @[Switch.scala 41:38:@36468.4]
  wire  _T_75311; // @[Switch.scala 41:52:@36470.4]
  wire  output_61_58; // @[Switch.scala 41:38:@36471.4]
  wire  _T_75314; // @[Switch.scala 41:52:@36473.4]
  wire  output_61_59; // @[Switch.scala 41:38:@36474.4]
  wire  _T_75317; // @[Switch.scala 41:52:@36476.4]
  wire  output_61_60; // @[Switch.scala 41:38:@36477.4]
  wire  _T_75320; // @[Switch.scala 41:52:@36479.4]
  wire  output_61_61; // @[Switch.scala 41:38:@36480.4]
  wire  _T_75323; // @[Switch.scala 41:52:@36482.4]
  wire  output_61_62; // @[Switch.scala 41:38:@36483.4]
  wire  _T_75326; // @[Switch.scala 41:52:@36485.4]
  wire  output_61_63; // @[Switch.scala 41:38:@36486.4]
  wire [7:0] _T_75334; // @[Switch.scala 43:31:@36494.4]
  wire [15:0] _T_75342; // @[Switch.scala 43:31:@36502.4]
  wire [7:0] _T_75349; // @[Switch.scala 43:31:@36509.4]
  wire [31:0] _T_75358; // @[Switch.scala 43:31:@36518.4]
  wire [7:0] _T_75365; // @[Switch.scala 43:31:@36525.4]
  wire [15:0] _T_75373; // @[Switch.scala 43:31:@36533.4]
  wire [7:0] _T_75380; // @[Switch.scala 43:31:@36540.4]
  wire [31:0] _T_75389; // @[Switch.scala 43:31:@36549.4]
  wire [63:0] _T_75390; // @[Switch.scala 43:31:@36550.4]
  wire  _T_75394; // @[Switch.scala 41:52:@36553.4]
  wire  output_62_0; // @[Switch.scala 41:38:@36554.4]
  wire  _T_75397; // @[Switch.scala 41:52:@36556.4]
  wire  output_62_1; // @[Switch.scala 41:38:@36557.4]
  wire  _T_75400; // @[Switch.scala 41:52:@36559.4]
  wire  output_62_2; // @[Switch.scala 41:38:@36560.4]
  wire  _T_75403; // @[Switch.scala 41:52:@36562.4]
  wire  output_62_3; // @[Switch.scala 41:38:@36563.4]
  wire  _T_75406; // @[Switch.scala 41:52:@36565.4]
  wire  output_62_4; // @[Switch.scala 41:38:@36566.4]
  wire  _T_75409; // @[Switch.scala 41:52:@36568.4]
  wire  output_62_5; // @[Switch.scala 41:38:@36569.4]
  wire  _T_75412; // @[Switch.scala 41:52:@36571.4]
  wire  output_62_6; // @[Switch.scala 41:38:@36572.4]
  wire  _T_75415; // @[Switch.scala 41:52:@36574.4]
  wire  output_62_7; // @[Switch.scala 41:38:@36575.4]
  wire  _T_75418; // @[Switch.scala 41:52:@36577.4]
  wire  output_62_8; // @[Switch.scala 41:38:@36578.4]
  wire  _T_75421; // @[Switch.scala 41:52:@36580.4]
  wire  output_62_9; // @[Switch.scala 41:38:@36581.4]
  wire  _T_75424; // @[Switch.scala 41:52:@36583.4]
  wire  output_62_10; // @[Switch.scala 41:38:@36584.4]
  wire  _T_75427; // @[Switch.scala 41:52:@36586.4]
  wire  output_62_11; // @[Switch.scala 41:38:@36587.4]
  wire  _T_75430; // @[Switch.scala 41:52:@36589.4]
  wire  output_62_12; // @[Switch.scala 41:38:@36590.4]
  wire  _T_75433; // @[Switch.scala 41:52:@36592.4]
  wire  output_62_13; // @[Switch.scala 41:38:@36593.4]
  wire  _T_75436; // @[Switch.scala 41:52:@36595.4]
  wire  output_62_14; // @[Switch.scala 41:38:@36596.4]
  wire  _T_75439; // @[Switch.scala 41:52:@36598.4]
  wire  output_62_15; // @[Switch.scala 41:38:@36599.4]
  wire  _T_75442; // @[Switch.scala 41:52:@36601.4]
  wire  output_62_16; // @[Switch.scala 41:38:@36602.4]
  wire  _T_75445; // @[Switch.scala 41:52:@36604.4]
  wire  output_62_17; // @[Switch.scala 41:38:@36605.4]
  wire  _T_75448; // @[Switch.scala 41:52:@36607.4]
  wire  output_62_18; // @[Switch.scala 41:38:@36608.4]
  wire  _T_75451; // @[Switch.scala 41:52:@36610.4]
  wire  output_62_19; // @[Switch.scala 41:38:@36611.4]
  wire  _T_75454; // @[Switch.scala 41:52:@36613.4]
  wire  output_62_20; // @[Switch.scala 41:38:@36614.4]
  wire  _T_75457; // @[Switch.scala 41:52:@36616.4]
  wire  output_62_21; // @[Switch.scala 41:38:@36617.4]
  wire  _T_75460; // @[Switch.scala 41:52:@36619.4]
  wire  output_62_22; // @[Switch.scala 41:38:@36620.4]
  wire  _T_75463; // @[Switch.scala 41:52:@36622.4]
  wire  output_62_23; // @[Switch.scala 41:38:@36623.4]
  wire  _T_75466; // @[Switch.scala 41:52:@36625.4]
  wire  output_62_24; // @[Switch.scala 41:38:@36626.4]
  wire  _T_75469; // @[Switch.scala 41:52:@36628.4]
  wire  output_62_25; // @[Switch.scala 41:38:@36629.4]
  wire  _T_75472; // @[Switch.scala 41:52:@36631.4]
  wire  output_62_26; // @[Switch.scala 41:38:@36632.4]
  wire  _T_75475; // @[Switch.scala 41:52:@36634.4]
  wire  output_62_27; // @[Switch.scala 41:38:@36635.4]
  wire  _T_75478; // @[Switch.scala 41:52:@36637.4]
  wire  output_62_28; // @[Switch.scala 41:38:@36638.4]
  wire  _T_75481; // @[Switch.scala 41:52:@36640.4]
  wire  output_62_29; // @[Switch.scala 41:38:@36641.4]
  wire  _T_75484; // @[Switch.scala 41:52:@36643.4]
  wire  output_62_30; // @[Switch.scala 41:38:@36644.4]
  wire  _T_75487; // @[Switch.scala 41:52:@36646.4]
  wire  output_62_31; // @[Switch.scala 41:38:@36647.4]
  wire  _T_75490; // @[Switch.scala 41:52:@36649.4]
  wire  output_62_32; // @[Switch.scala 41:38:@36650.4]
  wire  _T_75493; // @[Switch.scala 41:52:@36652.4]
  wire  output_62_33; // @[Switch.scala 41:38:@36653.4]
  wire  _T_75496; // @[Switch.scala 41:52:@36655.4]
  wire  output_62_34; // @[Switch.scala 41:38:@36656.4]
  wire  _T_75499; // @[Switch.scala 41:52:@36658.4]
  wire  output_62_35; // @[Switch.scala 41:38:@36659.4]
  wire  _T_75502; // @[Switch.scala 41:52:@36661.4]
  wire  output_62_36; // @[Switch.scala 41:38:@36662.4]
  wire  _T_75505; // @[Switch.scala 41:52:@36664.4]
  wire  output_62_37; // @[Switch.scala 41:38:@36665.4]
  wire  _T_75508; // @[Switch.scala 41:52:@36667.4]
  wire  output_62_38; // @[Switch.scala 41:38:@36668.4]
  wire  _T_75511; // @[Switch.scala 41:52:@36670.4]
  wire  output_62_39; // @[Switch.scala 41:38:@36671.4]
  wire  _T_75514; // @[Switch.scala 41:52:@36673.4]
  wire  output_62_40; // @[Switch.scala 41:38:@36674.4]
  wire  _T_75517; // @[Switch.scala 41:52:@36676.4]
  wire  output_62_41; // @[Switch.scala 41:38:@36677.4]
  wire  _T_75520; // @[Switch.scala 41:52:@36679.4]
  wire  output_62_42; // @[Switch.scala 41:38:@36680.4]
  wire  _T_75523; // @[Switch.scala 41:52:@36682.4]
  wire  output_62_43; // @[Switch.scala 41:38:@36683.4]
  wire  _T_75526; // @[Switch.scala 41:52:@36685.4]
  wire  output_62_44; // @[Switch.scala 41:38:@36686.4]
  wire  _T_75529; // @[Switch.scala 41:52:@36688.4]
  wire  output_62_45; // @[Switch.scala 41:38:@36689.4]
  wire  _T_75532; // @[Switch.scala 41:52:@36691.4]
  wire  output_62_46; // @[Switch.scala 41:38:@36692.4]
  wire  _T_75535; // @[Switch.scala 41:52:@36694.4]
  wire  output_62_47; // @[Switch.scala 41:38:@36695.4]
  wire  _T_75538; // @[Switch.scala 41:52:@36697.4]
  wire  output_62_48; // @[Switch.scala 41:38:@36698.4]
  wire  _T_75541; // @[Switch.scala 41:52:@36700.4]
  wire  output_62_49; // @[Switch.scala 41:38:@36701.4]
  wire  _T_75544; // @[Switch.scala 41:52:@36703.4]
  wire  output_62_50; // @[Switch.scala 41:38:@36704.4]
  wire  _T_75547; // @[Switch.scala 41:52:@36706.4]
  wire  output_62_51; // @[Switch.scala 41:38:@36707.4]
  wire  _T_75550; // @[Switch.scala 41:52:@36709.4]
  wire  output_62_52; // @[Switch.scala 41:38:@36710.4]
  wire  _T_75553; // @[Switch.scala 41:52:@36712.4]
  wire  output_62_53; // @[Switch.scala 41:38:@36713.4]
  wire  _T_75556; // @[Switch.scala 41:52:@36715.4]
  wire  output_62_54; // @[Switch.scala 41:38:@36716.4]
  wire  _T_75559; // @[Switch.scala 41:52:@36718.4]
  wire  output_62_55; // @[Switch.scala 41:38:@36719.4]
  wire  _T_75562; // @[Switch.scala 41:52:@36721.4]
  wire  output_62_56; // @[Switch.scala 41:38:@36722.4]
  wire  _T_75565; // @[Switch.scala 41:52:@36724.4]
  wire  output_62_57; // @[Switch.scala 41:38:@36725.4]
  wire  _T_75568; // @[Switch.scala 41:52:@36727.4]
  wire  output_62_58; // @[Switch.scala 41:38:@36728.4]
  wire  _T_75571; // @[Switch.scala 41:52:@36730.4]
  wire  output_62_59; // @[Switch.scala 41:38:@36731.4]
  wire  _T_75574; // @[Switch.scala 41:52:@36733.4]
  wire  output_62_60; // @[Switch.scala 41:38:@36734.4]
  wire  _T_75577; // @[Switch.scala 41:52:@36736.4]
  wire  output_62_61; // @[Switch.scala 41:38:@36737.4]
  wire  _T_75580; // @[Switch.scala 41:52:@36739.4]
  wire  output_62_62; // @[Switch.scala 41:38:@36740.4]
  wire  _T_75583; // @[Switch.scala 41:52:@36742.4]
  wire  output_62_63; // @[Switch.scala 41:38:@36743.4]
  wire [7:0] _T_75591; // @[Switch.scala 43:31:@36751.4]
  wire [15:0] _T_75599; // @[Switch.scala 43:31:@36759.4]
  wire [7:0] _T_75606; // @[Switch.scala 43:31:@36766.4]
  wire [31:0] _T_75615; // @[Switch.scala 43:31:@36775.4]
  wire [7:0] _T_75622; // @[Switch.scala 43:31:@36782.4]
  wire [15:0] _T_75630; // @[Switch.scala 43:31:@36790.4]
  wire [7:0] _T_75637; // @[Switch.scala 43:31:@36797.4]
  wire [31:0] _T_75646; // @[Switch.scala 43:31:@36806.4]
  wire [63:0] _T_75647; // @[Switch.scala 43:31:@36807.4]
  wire  _T_75651; // @[Switch.scala 41:52:@36810.4]
  wire  output_63_0; // @[Switch.scala 41:38:@36811.4]
  wire  _T_75654; // @[Switch.scala 41:52:@36813.4]
  wire  output_63_1; // @[Switch.scala 41:38:@36814.4]
  wire  _T_75657; // @[Switch.scala 41:52:@36816.4]
  wire  output_63_2; // @[Switch.scala 41:38:@36817.4]
  wire  _T_75660; // @[Switch.scala 41:52:@36819.4]
  wire  output_63_3; // @[Switch.scala 41:38:@36820.4]
  wire  _T_75663; // @[Switch.scala 41:52:@36822.4]
  wire  output_63_4; // @[Switch.scala 41:38:@36823.4]
  wire  _T_75666; // @[Switch.scala 41:52:@36825.4]
  wire  output_63_5; // @[Switch.scala 41:38:@36826.4]
  wire  _T_75669; // @[Switch.scala 41:52:@36828.4]
  wire  output_63_6; // @[Switch.scala 41:38:@36829.4]
  wire  _T_75672; // @[Switch.scala 41:52:@36831.4]
  wire  output_63_7; // @[Switch.scala 41:38:@36832.4]
  wire  _T_75675; // @[Switch.scala 41:52:@36834.4]
  wire  output_63_8; // @[Switch.scala 41:38:@36835.4]
  wire  _T_75678; // @[Switch.scala 41:52:@36837.4]
  wire  output_63_9; // @[Switch.scala 41:38:@36838.4]
  wire  _T_75681; // @[Switch.scala 41:52:@36840.4]
  wire  output_63_10; // @[Switch.scala 41:38:@36841.4]
  wire  _T_75684; // @[Switch.scala 41:52:@36843.4]
  wire  output_63_11; // @[Switch.scala 41:38:@36844.4]
  wire  _T_75687; // @[Switch.scala 41:52:@36846.4]
  wire  output_63_12; // @[Switch.scala 41:38:@36847.4]
  wire  _T_75690; // @[Switch.scala 41:52:@36849.4]
  wire  output_63_13; // @[Switch.scala 41:38:@36850.4]
  wire  _T_75693; // @[Switch.scala 41:52:@36852.4]
  wire  output_63_14; // @[Switch.scala 41:38:@36853.4]
  wire  _T_75696; // @[Switch.scala 41:52:@36855.4]
  wire  output_63_15; // @[Switch.scala 41:38:@36856.4]
  wire  _T_75699; // @[Switch.scala 41:52:@36858.4]
  wire  output_63_16; // @[Switch.scala 41:38:@36859.4]
  wire  _T_75702; // @[Switch.scala 41:52:@36861.4]
  wire  output_63_17; // @[Switch.scala 41:38:@36862.4]
  wire  _T_75705; // @[Switch.scala 41:52:@36864.4]
  wire  output_63_18; // @[Switch.scala 41:38:@36865.4]
  wire  _T_75708; // @[Switch.scala 41:52:@36867.4]
  wire  output_63_19; // @[Switch.scala 41:38:@36868.4]
  wire  _T_75711; // @[Switch.scala 41:52:@36870.4]
  wire  output_63_20; // @[Switch.scala 41:38:@36871.4]
  wire  _T_75714; // @[Switch.scala 41:52:@36873.4]
  wire  output_63_21; // @[Switch.scala 41:38:@36874.4]
  wire  _T_75717; // @[Switch.scala 41:52:@36876.4]
  wire  output_63_22; // @[Switch.scala 41:38:@36877.4]
  wire  _T_75720; // @[Switch.scala 41:52:@36879.4]
  wire  output_63_23; // @[Switch.scala 41:38:@36880.4]
  wire  _T_75723; // @[Switch.scala 41:52:@36882.4]
  wire  output_63_24; // @[Switch.scala 41:38:@36883.4]
  wire  _T_75726; // @[Switch.scala 41:52:@36885.4]
  wire  output_63_25; // @[Switch.scala 41:38:@36886.4]
  wire  _T_75729; // @[Switch.scala 41:52:@36888.4]
  wire  output_63_26; // @[Switch.scala 41:38:@36889.4]
  wire  _T_75732; // @[Switch.scala 41:52:@36891.4]
  wire  output_63_27; // @[Switch.scala 41:38:@36892.4]
  wire  _T_75735; // @[Switch.scala 41:52:@36894.4]
  wire  output_63_28; // @[Switch.scala 41:38:@36895.4]
  wire  _T_75738; // @[Switch.scala 41:52:@36897.4]
  wire  output_63_29; // @[Switch.scala 41:38:@36898.4]
  wire  _T_75741; // @[Switch.scala 41:52:@36900.4]
  wire  output_63_30; // @[Switch.scala 41:38:@36901.4]
  wire  _T_75744; // @[Switch.scala 41:52:@36903.4]
  wire  output_63_31; // @[Switch.scala 41:38:@36904.4]
  wire  _T_75747; // @[Switch.scala 41:52:@36906.4]
  wire  output_63_32; // @[Switch.scala 41:38:@36907.4]
  wire  _T_75750; // @[Switch.scala 41:52:@36909.4]
  wire  output_63_33; // @[Switch.scala 41:38:@36910.4]
  wire  _T_75753; // @[Switch.scala 41:52:@36912.4]
  wire  output_63_34; // @[Switch.scala 41:38:@36913.4]
  wire  _T_75756; // @[Switch.scala 41:52:@36915.4]
  wire  output_63_35; // @[Switch.scala 41:38:@36916.4]
  wire  _T_75759; // @[Switch.scala 41:52:@36918.4]
  wire  output_63_36; // @[Switch.scala 41:38:@36919.4]
  wire  _T_75762; // @[Switch.scala 41:52:@36921.4]
  wire  output_63_37; // @[Switch.scala 41:38:@36922.4]
  wire  _T_75765; // @[Switch.scala 41:52:@36924.4]
  wire  output_63_38; // @[Switch.scala 41:38:@36925.4]
  wire  _T_75768; // @[Switch.scala 41:52:@36927.4]
  wire  output_63_39; // @[Switch.scala 41:38:@36928.4]
  wire  _T_75771; // @[Switch.scala 41:52:@36930.4]
  wire  output_63_40; // @[Switch.scala 41:38:@36931.4]
  wire  _T_75774; // @[Switch.scala 41:52:@36933.4]
  wire  output_63_41; // @[Switch.scala 41:38:@36934.4]
  wire  _T_75777; // @[Switch.scala 41:52:@36936.4]
  wire  output_63_42; // @[Switch.scala 41:38:@36937.4]
  wire  _T_75780; // @[Switch.scala 41:52:@36939.4]
  wire  output_63_43; // @[Switch.scala 41:38:@36940.4]
  wire  _T_75783; // @[Switch.scala 41:52:@36942.4]
  wire  output_63_44; // @[Switch.scala 41:38:@36943.4]
  wire  _T_75786; // @[Switch.scala 41:52:@36945.4]
  wire  output_63_45; // @[Switch.scala 41:38:@36946.4]
  wire  _T_75789; // @[Switch.scala 41:52:@36948.4]
  wire  output_63_46; // @[Switch.scala 41:38:@36949.4]
  wire  _T_75792; // @[Switch.scala 41:52:@36951.4]
  wire  output_63_47; // @[Switch.scala 41:38:@36952.4]
  wire  _T_75795; // @[Switch.scala 41:52:@36954.4]
  wire  output_63_48; // @[Switch.scala 41:38:@36955.4]
  wire  _T_75798; // @[Switch.scala 41:52:@36957.4]
  wire  output_63_49; // @[Switch.scala 41:38:@36958.4]
  wire  _T_75801; // @[Switch.scala 41:52:@36960.4]
  wire  output_63_50; // @[Switch.scala 41:38:@36961.4]
  wire  _T_75804; // @[Switch.scala 41:52:@36963.4]
  wire  output_63_51; // @[Switch.scala 41:38:@36964.4]
  wire  _T_75807; // @[Switch.scala 41:52:@36966.4]
  wire  output_63_52; // @[Switch.scala 41:38:@36967.4]
  wire  _T_75810; // @[Switch.scala 41:52:@36969.4]
  wire  output_63_53; // @[Switch.scala 41:38:@36970.4]
  wire  _T_75813; // @[Switch.scala 41:52:@36972.4]
  wire  output_63_54; // @[Switch.scala 41:38:@36973.4]
  wire  _T_75816; // @[Switch.scala 41:52:@36975.4]
  wire  output_63_55; // @[Switch.scala 41:38:@36976.4]
  wire  _T_75819; // @[Switch.scala 41:52:@36978.4]
  wire  output_63_56; // @[Switch.scala 41:38:@36979.4]
  wire  _T_75822; // @[Switch.scala 41:52:@36981.4]
  wire  output_63_57; // @[Switch.scala 41:38:@36982.4]
  wire  _T_75825; // @[Switch.scala 41:52:@36984.4]
  wire  output_63_58; // @[Switch.scala 41:38:@36985.4]
  wire  _T_75828; // @[Switch.scala 41:52:@36987.4]
  wire  output_63_59; // @[Switch.scala 41:38:@36988.4]
  wire  _T_75831; // @[Switch.scala 41:52:@36990.4]
  wire  output_63_60; // @[Switch.scala 41:38:@36991.4]
  wire  _T_75834; // @[Switch.scala 41:52:@36993.4]
  wire  output_63_61; // @[Switch.scala 41:38:@36994.4]
  wire  _T_75837; // @[Switch.scala 41:52:@36996.4]
  wire  output_63_62; // @[Switch.scala 41:38:@36997.4]
  wire  _T_75840; // @[Switch.scala 41:52:@36999.4]
  wire  output_63_63; // @[Switch.scala 41:38:@37000.4]
  wire [7:0] _T_75848; // @[Switch.scala 43:31:@37008.4]
  wire [15:0] _T_75856; // @[Switch.scala 43:31:@37016.4]
  wire [7:0] _T_75863; // @[Switch.scala 43:31:@37023.4]
  wire [31:0] _T_75872; // @[Switch.scala 43:31:@37032.4]
  wire [7:0] _T_75879; // @[Switch.scala 43:31:@37039.4]
  wire [15:0] _T_75887; // @[Switch.scala 43:31:@37047.4]
  wire [7:0] _T_75894; // @[Switch.scala 43:31:@37054.4]
  wire [31:0] _T_75903; // @[Switch.scala 43:31:@37063.4]
  wire [63:0] _T_75904; // @[Switch.scala 43:31:@37064.4]
  assign _T_17654 = io_inAddr_0 == 6'h0; // @[Switch.scala 30:53:@10.4]
  assign valid_0_0 = io_inValid_0 & _T_17654; // @[Switch.scala 30:36:@11.4]
  assign _T_17657 = io_inAddr_1 == 6'h0; // @[Switch.scala 30:53:@13.4]
  assign valid_0_1 = io_inValid_1 & _T_17657; // @[Switch.scala 30:36:@14.4]
  assign _T_17660 = io_inAddr_2 == 6'h0; // @[Switch.scala 30:53:@16.4]
  assign valid_0_2 = io_inValid_2 & _T_17660; // @[Switch.scala 30:36:@17.4]
  assign _T_17663 = io_inAddr_3 == 6'h0; // @[Switch.scala 30:53:@19.4]
  assign valid_0_3 = io_inValid_3 & _T_17663; // @[Switch.scala 30:36:@20.4]
  assign _T_17666 = io_inAddr_4 == 6'h0; // @[Switch.scala 30:53:@22.4]
  assign valid_0_4 = io_inValid_4 & _T_17666; // @[Switch.scala 30:36:@23.4]
  assign _T_17669 = io_inAddr_5 == 6'h0; // @[Switch.scala 30:53:@25.4]
  assign valid_0_5 = io_inValid_5 & _T_17669; // @[Switch.scala 30:36:@26.4]
  assign _T_17672 = io_inAddr_6 == 6'h0; // @[Switch.scala 30:53:@28.4]
  assign valid_0_6 = io_inValid_6 & _T_17672; // @[Switch.scala 30:36:@29.4]
  assign _T_17675 = io_inAddr_7 == 6'h0; // @[Switch.scala 30:53:@31.4]
  assign valid_0_7 = io_inValid_7 & _T_17675; // @[Switch.scala 30:36:@32.4]
  assign _T_17678 = io_inAddr_8 == 6'h0; // @[Switch.scala 30:53:@34.4]
  assign valid_0_8 = io_inValid_8 & _T_17678; // @[Switch.scala 30:36:@35.4]
  assign _T_17681 = io_inAddr_9 == 6'h0; // @[Switch.scala 30:53:@37.4]
  assign valid_0_9 = io_inValid_9 & _T_17681; // @[Switch.scala 30:36:@38.4]
  assign _T_17684 = io_inAddr_10 == 6'h0; // @[Switch.scala 30:53:@40.4]
  assign valid_0_10 = io_inValid_10 & _T_17684; // @[Switch.scala 30:36:@41.4]
  assign _T_17687 = io_inAddr_11 == 6'h0; // @[Switch.scala 30:53:@43.4]
  assign valid_0_11 = io_inValid_11 & _T_17687; // @[Switch.scala 30:36:@44.4]
  assign _T_17690 = io_inAddr_12 == 6'h0; // @[Switch.scala 30:53:@46.4]
  assign valid_0_12 = io_inValid_12 & _T_17690; // @[Switch.scala 30:36:@47.4]
  assign _T_17693 = io_inAddr_13 == 6'h0; // @[Switch.scala 30:53:@49.4]
  assign valid_0_13 = io_inValid_13 & _T_17693; // @[Switch.scala 30:36:@50.4]
  assign _T_17696 = io_inAddr_14 == 6'h0; // @[Switch.scala 30:53:@52.4]
  assign valid_0_14 = io_inValid_14 & _T_17696; // @[Switch.scala 30:36:@53.4]
  assign _T_17699 = io_inAddr_15 == 6'h0; // @[Switch.scala 30:53:@55.4]
  assign valid_0_15 = io_inValid_15 & _T_17699; // @[Switch.scala 30:36:@56.4]
  assign _T_17702 = io_inAddr_16 == 6'h0; // @[Switch.scala 30:53:@58.4]
  assign valid_0_16 = io_inValid_16 & _T_17702; // @[Switch.scala 30:36:@59.4]
  assign _T_17705 = io_inAddr_17 == 6'h0; // @[Switch.scala 30:53:@61.4]
  assign valid_0_17 = io_inValid_17 & _T_17705; // @[Switch.scala 30:36:@62.4]
  assign _T_17708 = io_inAddr_18 == 6'h0; // @[Switch.scala 30:53:@64.4]
  assign valid_0_18 = io_inValid_18 & _T_17708; // @[Switch.scala 30:36:@65.4]
  assign _T_17711 = io_inAddr_19 == 6'h0; // @[Switch.scala 30:53:@67.4]
  assign valid_0_19 = io_inValid_19 & _T_17711; // @[Switch.scala 30:36:@68.4]
  assign _T_17714 = io_inAddr_20 == 6'h0; // @[Switch.scala 30:53:@70.4]
  assign valid_0_20 = io_inValid_20 & _T_17714; // @[Switch.scala 30:36:@71.4]
  assign _T_17717 = io_inAddr_21 == 6'h0; // @[Switch.scala 30:53:@73.4]
  assign valid_0_21 = io_inValid_21 & _T_17717; // @[Switch.scala 30:36:@74.4]
  assign _T_17720 = io_inAddr_22 == 6'h0; // @[Switch.scala 30:53:@76.4]
  assign valid_0_22 = io_inValid_22 & _T_17720; // @[Switch.scala 30:36:@77.4]
  assign _T_17723 = io_inAddr_23 == 6'h0; // @[Switch.scala 30:53:@79.4]
  assign valid_0_23 = io_inValid_23 & _T_17723; // @[Switch.scala 30:36:@80.4]
  assign _T_17726 = io_inAddr_24 == 6'h0; // @[Switch.scala 30:53:@82.4]
  assign valid_0_24 = io_inValid_24 & _T_17726; // @[Switch.scala 30:36:@83.4]
  assign _T_17729 = io_inAddr_25 == 6'h0; // @[Switch.scala 30:53:@85.4]
  assign valid_0_25 = io_inValid_25 & _T_17729; // @[Switch.scala 30:36:@86.4]
  assign _T_17732 = io_inAddr_26 == 6'h0; // @[Switch.scala 30:53:@88.4]
  assign valid_0_26 = io_inValid_26 & _T_17732; // @[Switch.scala 30:36:@89.4]
  assign _T_17735 = io_inAddr_27 == 6'h0; // @[Switch.scala 30:53:@91.4]
  assign valid_0_27 = io_inValid_27 & _T_17735; // @[Switch.scala 30:36:@92.4]
  assign _T_17738 = io_inAddr_28 == 6'h0; // @[Switch.scala 30:53:@94.4]
  assign valid_0_28 = io_inValid_28 & _T_17738; // @[Switch.scala 30:36:@95.4]
  assign _T_17741 = io_inAddr_29 == 6'h0; // @[Switch.scala 30:53:@97.4]
  assign valid_0_29 = io_inValid_29 & _T_17741; // @[Switch.scala 30:36:@98.4]
  assign _T_17744 = io_inAddr_30 == 6'h0; // @[Switch.scala 30:53:@100.4]
  assign valid_0_30 = io_inValid_30 & _T_17744; // @[Switch.scala 30:36:@101.4]
  assign _T_17747 = io_inAddr_31 == 6'h0; // @[Switch.scala 30:53:@103.4]
  assign valid_0_31 = io_inValid_31 & _T_17747; // @[Switch.scala 30:36:@104.4]
  assign _T_17750 = io_inAddr_32 == 6'h0; // @[Switch.scala 30:53:@106.4]
  assign valid_0_32 = io_inValid_32 & _T_17750; // @[Switch.scala 30:36:@107.4]
  assign _T_17753 = io_inAddr_33 == 6'h0; // @[Switch.scala 30:53:@109.4]
  assign valid_0_33 = io_inValid_33 & _T_17753; // @[Switch.scala 30:36:@110.4]
  assign _T_17756 = io_inAddr_34 == 6'h0; // @[Switch.scala 30:53:@112.4]
  assign valid_0_34 = io_inValid_34 & _T_17756; // @[Switch.scala 30:36:@113.4]
  assign _T_17759 = io_inAddr_35 == 6'h0; // @[Switch.scala 30:53:@115.4]
  assign valid_0_35 = io_inValid_35 & _T_17759; // @[Switch.scala 30:36:@116.4]
  assign _T_17762 = io_inAddr_36 == 6'h0; // @[Switch.scala 30:53:@118.4]
  assign valid_0_36 = io_inValid_36 & _T_17762; // @[Switch.scala 30:36:@119.4]
  assign _T_17765 = io_inAddr_37 == 6'h0; // @[Switch.scala 30:53:@121.4]
  assign valid_0_37 = io_inValid_37 & _T_17765; // @[Switch.scala 30:36:@122.4]
  assign _T_17768 = io_inAddr_38 == 6'h0; // @[Switch.scala 30:53:@124.4]
  assign valid_0_38 = io_inValid_38 & _T_17768; // @[Switch.scala 30:36:@125.4]
  assign _T_17771 = io_inAddr_39 == 6'h0; // @[Switch.scala 30:53:@127.4]
  assign valid_0_39 = io_inValid_39 & _T_17771; // @[Switch.scala 30:36:@128.4]
  assign _T_17774 = io_inAddr_40 == 6'h0; // @[Switch.scala 30:53:@130.4]
  assign valid_0_40 = io_inValid_40 & _T_17774; // @[Switch.scala 30:36:@131.4]
  assign _T_17777 = io_inAddr_41 == 6'h0; // @[Switch.scala 30:53:@133.4]
  assign valid_0_41 = io_inValid_41 & _T_17777; // @[Switch.scala 30:36:@134.4]
  assign _T_17780 = io_inAddr_42 == 6'h0; // @[Switch.scala 30:53:@136.4]
  assign valid_0_42 = io_inValid_42 & _T_17780; // @[Switch.scala 30:36:@137.4]
  assign _T_17783 = io_inAddr_43 == 6'h0; // @[Switch.scala 30:53:@139.4]
  assign valid_0_43 = io_inValid_43 & _T_17783; // @[Switch.scala 30:36:@140.4]
  assign _T_17786 = io_inAddr_44 == 6'h0; // @[Switch.scala 30:53:@142.4]
  assign valid_0_44 = io_inValid_44 & _T_17786; // @[Switch.scala 30:36:@143.4]
  assign _T_17789 = io_inAddr_45 == 6'h0; // @[Switch.scala 30:53:@145.4]
  assign valid_0_45 = io_inValid_45 & _T_17789; // @[Switch.scala 30:36:@146.4]
  assign _T_17792 = io_inAddr_46 == 6'h0; // @[Switch.scala 30:53:@148.4]
  assign valid_0_46 = io_inValid_46 & _T_17792; // @[Switch.scala 30:36:@149.4]
  assign _T_17795 = io_inAddr_47 == 6'h0; // @[Switch.scala 30:53:@151.4]
  assign valid_0_47 = io_inValid_47 & _T_17795; // @[Switch.scala 30:36:@152.4]
  assign _T_17798 = io_inAddr_48 == 6'h0; // @[Switch.scala 30:53:@154.4]
  assign valid_0_48 = io_inValid_48 & _T_17798; // @[Switch.scala 30:36:@155.4]
  assign _T_17801 = io_inAddr_49 == 6'h0; // @[Switch.scala 30:53:@157.4]
  assign valid_0_49 = io_inValid_49 & _T_17801; // @[Switch.scala 30:36:@158.4]
  assign _T_17804 = io_inAddr_50 == 6'h0; // @[Switch.scala 30:53:@160.4]
  assign valid_0_50 = io_inValid_50 & _T_17804; // @[Switch.scala 30:36:@161.4]
  assign _T_17807 = io_inAddr_51 == 6'h0; // @[Switch.scala 30:53:@163.4]
  assign valid_0_51 = io_inValid_51 & _T_17807; // @[Switch.scala 30:36:@164.4]
  assign _T_17810 = io_inAddr_52 == 6'h0; // @[Switch.scala 30:53:@166.4]
  assign valid_0_52 = io_inValid_52 & _T_17810; // @[Switch.scala 30:36:@167.4]
  assign _T_17813 = io_inAddr_53 == 6'h0; // @[Switch.scala 30:53:@169.4]
  assign valid_0_53 = io_inValid_53 & _T_17813; // @[Switch.scala 30:36:@170.4]
  assign _T_17816 = io_inAddr_54 == 6'h0; // @[Switch.scala 30:53:@172.4]
  assign valid_0_54 = io_inValid_54 & _T_17816; // @[Switch.scala 30:36:@173.4]
  assign _T_17819 = io_inAddr_55 == 6'h0; // @[Switch.scala 30:53:@175.4]
  assign valid_0_55 = io_inValid_55 & _T_17819; // @[Switch.scala 30:36:@176.4]
  assign _T_17822 = io_inAddr_56 == 6'h0; // @[Switch.scala 30:53:@178.4]
  assign valid_0_56 = io_inValid_56 & _T_17822; // @[Switch.scala 30:36:@179.4]
  assign _T_17825 = io_inAddr_57 == 6'h0; // @[Switch.scala 30:53:@181.4]
  assign valid_0_57 = io_inValid_57 & _T_17825; // @[Switch.scala 30:36:@182.4]
  assign _T_17828 = io_inAddr_58 == 6'h0; // @[Switch.scala 30:53:@184.4]
  assign valid_0_58 = io_inValid_58 & _T_17828; // @[Switch.scala 30:36:@185.4]
  assign _T_17831 = io_inAddr_59 == 6'h0; // @[Switch.scala 30:53:@187.4]
  assign valid_0_59 = io_inValid_59 & _T_17831; // @[Switch.scala 30:36:@188.4]
  assign _T_17834 = io_inAddr_60 == 6'h0; // @[Switch.scala 30:53:@190.4]
  assign valid_0_60 = io_inValid_60 & _T_17834; // @[Switch.scala 30:36:@191.4]
  assign _T_17837 = io_inAddr_61 == 6'h0; // @[Switch.scala 30:53:@193.4]
  assign valid_0_61 = io_inValid_61 & _T_17837; // @[Switch.scala 30:36:@194.4]
  assign _T_17840 = io_inAddr_62 == 6'h0; // @[Switch.scala 30:53:@196.4]
  assign valid_0_62 = io_inValid_62 & _T_17840; // @[Switch.scala 30:36:@197.4]
  assign _T_17843 = io_inAddr_63 == 6'h0; // @[Switch.scala 30:53:@199.4]
  assign valid_0_63 = io_inValid_63 & _T_17843; // @[Switch.scala 30:36:@200.4]
  assign _T_17909 = valid_0_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@202.4]
  assign _T_17910 = valid_0_61 ? 6'h3d : _T_17909; // @[Mux.scala 31:69:@203.4]
  assign _T_17911 = valid_0_60 ? 6'h3c : _T_17910; // @[Mux.scala 31:69:@204.4]
  assign _T_17912 = valid_0_59 ? 6'h3b : _T_17911; // @[Mux.scala 31:69:@205.4]
  assign _T_17913 = valid_0_58 ? 6'h3a : _T_17912; // @[Mux.scala 31:69:@206.4]
  assign _T_17914 = valid_0_57 ? 6'h39 : _T_17913; // @[Mux.scala 31:69:@207.4]
  assign _T_17915 = valid_0_56 ? 6'h38 : _T_17914; // @[Mux.scala 31:69:@208.4]
  assign _T_17916 = valid_0_55 ? 6'h37 : _T_17915; // @[Mux.scala 31:69:@209.4]
  assign _T_17917 = valid_0_54 ? 6'h36 : _T_17916; // @[Mux.scala 31:69:@210.4]
  assign _T_17918 = valid_0_53 ? 6'h35 : _T_17917; // @[Mux.scala 31:69:@211.4]
  assign _T_17919 = valid_0_52 ? 6'h34 : _T_17918; // @[Mux.scala 31:69:@212.4]
  assign _T_17920 = valid_0_51 ? 6'h33 : _T_17919; // @[Mux.scala 31:69:@213.4]
  assign _T_17921 = valid_0_50 ? 6'h32 : _T_17920; // @[Mux.scala 31:69:@214.4]
  assign _T_17922 = valid_0_49 ? 6'h31 : _T_17921; // @[Mux.scala 31:69:@215.4]
  assign _T_17923 = valid_0_48 ? 6'h30 : _T_17922; // @[Mux.scala 31:69:@216.4]
  assign _T_17924 = valid_0_47 ? 6'h2f : _T_17923; // @[Mux.scala 31:69:@217.4]
  assign _T_17925 = valid_0_46 ? 6'h2e : _T_17924; // @[Mux.scala 31:69:@218.4]
  assign _T_17926 = valid_0_45 ? 6'h2d : _T_17925; // @[Mux.scala 31:69:@219.4]
  assign _T_17927 = valid_0_44 ? 6'h2c : _T_17926; // @[Mux.scala 31:69:@220.4]
  assign _T_17928 = valid_0_43 ? 6'h2b : _T_17927; // @[Mux.scala 31:69:@221.4]
  assign _T_17929 = valid_0_42 ? 6'h2a : _T_17928; // @[Mux.scala 31:69:@222.4]
  assign _T_17930 = valid_0_41 ? 6'h29 : _T_17929; // @[Mux.scala 31:69:@223.4]
  assign _T_17931 = valid_0_40 ? 6'h28 : _T_17930; // @[Mux.scala 31:69:@224.4]
  assign _T_17932 = valid_0_39 ? 6'h27 : _T_17931; // @[Mux.scala 31:69:@225.4]
  assign _T_17933 = valid_0_38 ? 6'h26 : _T_17932; // @[Mux.scala 31:69:@226.4]
  assign _T_17934 = valid_0_37 ? 6'h25 : _T_17933; // @[Mux.scala 31:69:@227.4]
  assign _T_17935 = valid_0_36 ? 6'h24 : _T_17934; // @[Mux.scala 31:69:@228.4]
  assign _T_17936 = valid_0_35 ? 6'h23 : _T_17935; // @[Mux.scala 31:69:@229.4]
  assign _T_17937 = valid_0_34 ? 6'h22 : _T_17936; // @[Mux.scala 31:69:@230.4]
  assign _T_17938 = valid_0_33 ? 6'h21 : _T_17937; // @[Mux.scala 31:69:@231.4]
  assign _T_17939 = valid_0_32 ? 6'h20 : _T_17938; // @[Mux.scala 31:69:@232.4]
  assign _T_17940 = valid_0_31 ? 6'h1f : _T_17939; // @[Mux.scala 31:69:@233.4]
  assign _T_17941 = valid_0_30 ? 6'h1e : _T_17940; // @[Mux.scala 31:69:@234.4]
  assign _T_17942 = valid_0_29 ? 6'h1d : _T_17941; // @[Mux.scala 31:69:@235.4]
  assign _T_17943 = valid_0_28 ? 6'h1c : _T_17942; // @[Mux.scala 31:69:@236.4]
  assign _T_17944 = valid_0_27 ? 6'h1b : _T_17943; // @[Mux.scala 31:69:@237.4]
  assign _T_17945 = valid_0_26 ? 6'h1a : _T_17944; // @[Mux.scala 31:69:@238.4]
  assign _T_17946 = valid_0_25 ? 6'h19 : _T_17945; // @[Mux.scala 31:69:@239.4]
  assign _T_17947 = valid_0_24 ? 6'h18 : _T_17946; // @[Mux.scala 31:69:@240.4]
  assign _T_17948 = valid_0_23 ? 6'h17 : _T_17947; // @[Mux.scala 31:69:@241.4]
  assign _T_17949 = valid_0_22 ? 6'h16 : _T_17948; // @[Mux.scala 31:69:@242.4]
  assign _T_17950 = valid_0_21 ? 6'h15 : _T_17949; // @[Mux.scala 31:69:@243.4]
  assign _T_17951 = valid_0_20 ? 6'h14 : _T_17950; // @[Mux.scala 31:69:@244.4]
  assign _T_17952 = valid_0_19 ? 6'h13 : _T_17951; // @[Mux.scala 31:69:@245.4]
  assign _T_17953 = valid_0_18 ? 6'h12 : _T_17952; // @[Mux.scala 31:69:@246.4]
  assign _T_17954 = valid_0_17 ? 6'h11 : _T_17953; // @[Mux.scala 31:69:@247.4]
  assign _T_17955 = valid_0_16 ? 6'h10 : _T_17954; // @[Mux.scala 31:69:@248.4]
  assign _T_17956 = valid_0_15 ? 6'hf : _T_17955; // @[Mux.scala 31:69:@249.4]
  assign _T_17957 = valid_0_14 ? 6'he : _T_17956; // @[Mux.scala 31:69:@250.4]
  assign _T_17958 = valid_0_13 ? 6'hd : _T_17957; // @[Mux.scala 31:69:@251.4]
  assign _T_17959 = valid_0_12 ? 6'hc : _T_17958; // @[Mux.scala 31:69:@252.4]
  assign _T_17960 = valid_0_11 ? 6'hb : _T_17959; // @[Mux.scala 31:69:@253.4]
  assign _T_17961 = valid_0_10 ? 6'ha : _T_17960; // @[Mux.scala 31:69:@254.4]
  assign _T_17962 = valid_0_9 ? 6'h9 : _T_17961; // @[Mux.scala 31:69:@255.4]
  assign _T_17963 = valid_0_8 ? 6'h8 : _T_17962; // @[Mux.scala 31:69:@256.4]
  assign _T_17964 = valid_0_7 ? 6'h7 : _T_17963; // @[Mux.scala 31:69:@257.4]
  assign _T_17965 = valid_0_6 ? 6'h6 : _T_17964; // @[Mux.scala 31:69:@258.4]
  assign _T_17966 = valid_0_5 ? 6'h5 : _T_17965; // @[Mux.scala 31:69:@259.4]
  assign _T_17967 = valid_0_4 ? 6'h4 : _T_17966; // @[Mux.scala 31:69:@260.4]
  assign _T_17968 = valid_0_3 ? 6'h3 : _T_17967; // @[Mux.scala 31:69:@261.4]
  assign _T_17969 = valid_0_2 ? 6'h2 : _T_17968; // @[Mux.scala 31:69:@262.4]
  assign _T_17970 = valid_0_1 ? 6'h1 : _T_17969; // @[Mux.scala 31:69:@263.4]
  assign select_0 = valid_0_0 ? 6'h0 : _T_17970; // @[Mux.scala 31:69:@264.4]
  assign _GEN_1 = 6'h1 == select_0 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@266.4]
  assign _GEN_2 = 6'h2 == select_0 ? io_inData_2 : _GEN_1; // @[Switch.scala 33:19:@266.4]
  assign _GEN_3 = 6'h3 == select_0 ? io_inData_3 : _GEN_2; // @[Switch.scala 33:19:@266.4]
  assign _GEN_4 = 6'h4 == select_0 ? io_inData_4 : _GEN_3; // @[Switch.scala 33:19:@266.4]
  assign _GEN_5 = 6'h5 == select_0 ? io_inData_5 : _GEN_4; // @[Switch.scala 33:19:@266.4]
  assign _GEN_6 = 6'h6 == select_0 ? io_inData_6 : _GEN_5; // @[Switch.scala 33:19:@266.4]
  assign _GEN_7 = 6'h7 == select_0 ? io_inData_7 : _GEN_6; // @[Switch.scala 33:19:@266.4]
  assign _GEN_8 = 6'h8 == select_0 ? io_inData_8 : _GEN_7; // @[Switch.scala 33:19:@266.4]
  assign _GEN_9 = 6'h9 == select_0 ? io_inData_9 : _GEN_8; // @[Switch.scala 33:19:@266.4]
  assign _GEN_10 = 6'ha == select_0 ? io_inData_10 : _GEN_9; // @[Switch.scala 33:19:@266.4]
  assign _GEN_11 = 6'hb == select_0 ? io_inData_11 : _GEN_10; // @[Switch.scala 33:19:@266.4]
  assign _GEN_12 = 6'hc == select_0 ? io_inData_12 : _GEN_11; // @[Switch.scala 33:19:@266.4]
  assign _GEN_13 = 6'hd == select_0 ? io_inData_13 : _GEN_12; // @[Switch.scala 33:19:@266.4]
  assign _GEN_14 = 6'he == select_0 ? io_inData_14 : _GEN_13; // @[Switch.scala 33:19:@266.4]
  assign _GEN_15 = 6'hf == select_0 ? io_inData_15 : _GEN_14; // @[Switch.scala 33:19:@266.4]
  assign _GEN_16 = 6'h10 == select_0 ? io_inData_16 : _GEN_15; // @[Switch.scala 33:19:@266.4]
  assign _GEN_17 = 6'h11 == select_0 ? io_inData_17 : _GEN_16; // @[Switch.scala 33:19:@266.4]
  assign _GEN_18 = 6'h12 == select_0 ? io_inData_18 : _GEN_17; // @[Switch.scala 33:19:@266.4]
  assign _GEN_19 = 6'h13 == select_0 ? io_inData_19 : _GEN_18; // @[Switch.scala 33:19:@266.4]
  assign _GEN_20 = 6'h14 == select_0 ? io_inData_20 : _GEN_19; // @[Switch.scala 33:19:@266.4]
  assign _GEN_21 = 6'h15 == select_0 ? io_inData_21 : _GEN_20; // @[Switch.scala 33:19:@266.4]
  assign _GEN_22 = 6'h16 == select_0 ? io_inData_22 : _GEN_21; // @[Switch.scala 33:19:@266.4]
  assign _GEN_23 = 6'h17 == select_0 ? io_inData_23 : _GEN_22; // @[Switch.scala 33:19:@266.4]
  assign _GEN_24 = 6'h18 == select_0 ? io_inData_24 : _GEN_23; // @[Switch.scala 33:19:@266.4]
  assign _GEN_25 = 6'h19 == select_0 ? io_inData_25 : _GEN_24; // @[Switch.scala 33:19:@266.4]
  assign _GEN_26 = 6'h1a == select_0 ? io_inData_26 : _GEN_25; // @[Switch.scala 33:19:@266.4]
  assign _GEN_27 = 6'h1b == select_0 ? io_inData_27 : _GEN_26; // @[Switch.scala 33:19:@266.4]
  assign _GEN_28 = 6'h1c == select_0 ? io_inData_28 : _GEN_27; // @[Switch.scala 33:19:@266.4]
  assign _GEN_29 = 6'h1d == select_0 ? io_inData_29 : _GEN_28; // @[Switch.scala 33:19:@266.4]
  assign _GEN_30 = 6'h1e == select_0 ? io_inData_30 : _GEN_29; // @[Switch.scala 33:19:@266.4]
  assign _GEN_31 = 6'h1f == select_0 ? io_inData_31 : _GEN_30; // @[Switch.scala 33:19:@266.4]
  assign _GEN_32 = 6'h20 == select_0 ? io_inData_32 : _GEN_31; // @[Switch.scala 33:19:@266.4]
  assign _GEN_33 = 6'h21 == select_0 ? io_inData_33 : _GEN_32; // @[Switch.scala 33:19:@266.4]
  assign _GEN_34 = 6'h22 == select_0 ? io_inData_34 : _GEN_33; // @[Switch.scala 33:19:@266.4]
  assign _GEN_35 = 6'h23 == select_0 ? io_inData_35 : _GEN_34; // @[Switch.scala 33:19:@266.4]
  assign _GEN_36 = 6'h24 == select_0 ? io_inData_36 : _GEN_35; // @[Switch.scala 33:19:@266.4]
  assign _GEN_37 = 6'h25 == select_0 ? io_inData_37 : _GEN_36; // @[Switch.scala 33:19:@266.4]
  assign _GEN_38 = 6'h26 == select_0 ? io_inData_38 : _GEN_37; // @[Switch.scala 33:19:@266.4]
  assign _GEN_39 = 6'h27 == select_0 ? io_inData_39 : _GEN_38; // @[Switch.scala 33:19:@266.4]
  assign _GEN_40 = 6'h28 == select_0 ? io_inData_40 : _GEN_39; // @[Switch.scala 33:19:@266.4]
  assign _GEN_41 = 6'h29 == select_0 ? io_inData_41 : _GEN_40; // @[Switch.scala 33:19:@266.4]
  assign _GEN_42 = 6'h2a == select_0 ? io_inData_42 : _GEN_41; // @[Switch.scala 33:19:@266.4]
  assign _GEN_43 = 6'h2b == select_0 ? io_inData_43 : _GEN_42; // @[Switch.scala 33:19:@266.4]
  assign _GEN_44 = 6'h2c == select_0 ? io_inData_44 : _GEN_43; // @[Switch.scala 33:19:@266.4]
  assign _GEN_45 = 6'h2d == select_0 ? io_inData_45 : _GEN_44; // @[Switch.scala 33:19:@266.4]
  assign _GEN_46 = 6'h2e == select_0 ? io_inData_46 : _GEN_45; // @[Switch.scala 33:19:@266.4]
  assign _GEN_47 = 6'h2f == select_0 ? io_inData_47 : _GEN_46; // @[Switch.scala 33:19:@266.4]
  assign _GEN_48 = 6'h30 == select_0 ? io_inData_48 : _GEN_47; // @[Switch.scala 33:19:@266.4]
  assign _GEN_49 = 6'h31 == select_0 ? io_inData_49 : _GEN_48; // @[Switch.scala 33:19:@266.4]
  assign _GEN_50 = 6'h32 == select_0 ? io_inData_50 : _GEN_49; // @[Switch.scala 33:19:@266.4]
  assign _GEN_51 = 6'h33 == select_0 ? io_inData_51 : _GEN_50; // @[Switch.scala 33:19:@266.4]
  assign _GEN_52 = 6'h34 == select_0 ? io_inData_52 : _GEN_51; // @[Switch.scala 33:19:@266.4]
  assign _GEN_53 = 6'h35 == select_0 ? io_inData_53 : _GEN_52; // @[Switch.scala 33:19:@266.4]
  assign _GEN_54 = 6'h36 == select_0 ? io_inData_54 : _GEN_53; // @[Switch.scala 33:19:@266.4]
  assign _GEN_55 = 6'h37 == select_0 ? io_inData_55 : _GEN_54; // @[Switch.scala 33:19:@266.4]
  assign _GEN_56 = 6'h38 == select_0 ? io_inData_56 : _GEN_55; // @[Switch.scala 33:19:@266.4]
  assign _GEN_57 = 6'h39 == select_0 ? io_inData_57 : _GEN_56; // @[Switch.scala 33:19:@266.4]
  assign _GEN_58 = 6'h3a == select_0 ? io_inData_58 : _GEN_57; // @[Switch.scala 33:19:@266.4]
  assign _GEN_59 = 6'h3b == select_0 ? io_inData_59 : _GEN_58; // @[Switch.scala 33:19:@266.4]
  assign _GEN_60 = 6'h3c == select_0 ? io_inData_60 : _GEN_59; // @[Switch.scala 33:19:@266.4]
  assign _GEN_61 = 6'h3d == select_0 ? io_inData_61 : _GEN_60; // @[Switch.scala 33:19:@266.4]
  assign _GEN_62 = 6'h3e == select_0 ? io_inData_62 : _GEN_61; // @[Switch.scala 33:19:@266.4]
  assign _T_17979 = {valid_0_7,valid_0_6,valid_0_5,valid_0_4,valid_0_3,valid_0_2,valid_0_1,valid_0_0}; // @[Switch.scala 34:32:@273.4]
  assign _T_17987 = {valid_0_15,valid_0_14,valid_0_13,valid_0_12,valid_0_11,valid_0_10,valid_0_9,valid_0_8,_T_17979}; // @[Switch.scala 34:32:@281.4]
  assign _T_17994 = {valid_0_23,valid_0_22,valid_0_21,valid_0_20,valid_0_19,valid_0_18,valid_0_17,valid_0_16}; // @[Switch.scala 34:32:@288.4]
  assign _T_18003 = {valid_0_31,valid_0_30,valid_0_29,valid_0_28,valid_0_27,valid_0_26,valid_0_25,valid_0_24,_T_17994,_T_17987}; // @[Switch.scala 34:32:@297.4]
  assign _T_18010 = {valid_0_39,valid_0_38,valid_0_37,valid_0_36,valid_0_35,valid_0_34,valid_0_33,valid_0_32}; // @[Switch.scala 34:32:@304.4]
  assign _T_18018 = {valid_0_47,valid_0_46,valid_0_45,valid_0_44,valid_0_43,valid_0_42,valid_0_41,valid_0_40,_T_18010}; // @[Switch.scala 34:32:@312.4]
  assign _T_18025 = {valid_0_55,valid_0_54,valid_0_53,valid_0_52,valid_0_51,valid_0_50,valid_0_49,valid_0_48}; // @[Switch.scala 34:32:@319.4]
  assign _T_18034 = {valid_0_63,valid_0_62,valid_0_61,valid_0_60,valid_0_59,valid_0_58,valid_0_57,valid_0_56,_T_18025,_T_18018}; // @[Switch.scala 34:32:@328.4]
  assign _T_18035 = {_T_18034,_T_18003}; // @[Switch.scala 34:32:@329.4]
  assign _T_18039 = io_inAddr_0 == 6'h1; // @[Switch.scala 30:53:@332.4]
  assign valid_1_0 = io_inValid_0 & _T_18039; // @[Switch.scala 30:36:@333.4]
  assign _T_18042 = io_inAddr_1 == 6'h1; // @[Switch.scala 30:53:@335.4]
  assign valid_1_1 = io_inValid_1 & _T_18042; // @[Switch.scala 30:36:@336.4]
  assign _T_18045 = io_inAddr_2 == 6'h1; // @[Switch.scala 30:53:@338.4]
  assign valid_1_2 = io_inValid_2 & _T_18045; // @[Switch.scala 30:36:@339.4]
  assign _T_18048 = io_inAddr_3 == 6'h1; // @[Switch.scala 30:53:@341.4]
  assign valid_1_3 = io_inValid_3 & _T_18048; // @[Switch.scala 30:36:@342.4]
  assign _T_18051 = io_inAddr_4 == 6'h1; // @[Switch.scala 30:53:@344.4]
  assign valid_1_4 = io_inValid_4 & _T_18051; // @[Switch.scala 30:36:@345.4]
  assign _T_18054 = io_inAddr_5 == 6'h1; // @[Switch.scala 30:53:@347.4]
  assign valid_1_5 = io_inValid_5 & _T_18054; // @[Switch.scala 30:36:@348.4]
  assign _T_18057 = io_inAddr_6 == 6'h1; // @[Switch.scala 30:53:@350.4]
  assign valid_1_6 = io_inValid_6 & _T_18057; // @[Switch.scala 30:36:@351.4]
  assign _T_18060 = io_inAddr_7 == 6'h1; // @[Switch.scala 30:53:@353.4]
  assign valid_1_7 = io_inValid_7 & _T_18060; // @[Switch.scala 30:36:@354.4]
  assign _T_18063 = io_inAddr_8 == 6'h1; // @[Switch.scala 30:53:@356.4]
  assign valid_1_8 = io_inValid_8 & _T_18063; // @[Switch.scala 30:36:@357.4]
  assign _T_18066 = io_inAddr_9 == 6'h1; // @[Switch.scala 30:53:@359.4]
  assign valid_1_9 = io_inValid_9 & _T_18066; // @[Switch.scala 30:36:@360.4]
  assign _T_18069 = io_inAddr_10 == 6'h1; // @[Switch.scala 30:53:@362.4]
  assign valid_1_10 = io_inValid_10 & _T_18069; // @[Switch.scala 30:36:@363.4]
  assign _T_18072 = io_inAddr_11 == 6'h1; // @[Switch.scala 30:53:@365.4]
  assign valid_1_11 = io_inValid_11 & _T_18072; // @[Switch.scala 30:36:@366.4]
  assign _T_18075 = io_inAddr_12 == 6'h1; // @[Switch.scala 30:53:@368.4]
  assign valid_1_12 = io_inValid_12 & _T_18075; // @[Switch.scala 30:36:@369.4]
  assign _T_18078 = io_inAddr_13 == 6'h1; // @[Switch.scala 30:53:@371.4]
  assign valid_1_13 = io_inValid_13 & _T_18078; // @[Switch.scala 30:36:@372.4]
  assign _T_18081 = io_inAddr_14 == 6'h1; // @[Switch.scala 30:53:@374.4]
  assign valid_1_14 = io_inValid_14 & _T_18081; // @[Switch.scala 30:36:@375.4]
  assign _T_18084 = io_inAddr_15 == 6'h1; // @[Switch.scala 30:53:@377.4]
  assign valid_1_15 = io_inValid_15 & _T_18084; // @[Switch.scala 30:36:@378.4]
  assign _T_18087 = io_inAddr_16 == 6'h1; // @[Switch.scala 30:53:@380.4]
  assign valid_1_16 = io_inValid_16 & _T_18087; // @[Switch.scala 30:36:@381.4]
  assign _T_18090 = io_inAddr_17 == 6'h1; // @[Switch.scala 30:53:@383.4]
  assign valid_1_17 = io_inValid_17 & _T_18090; // @[Switch.scala 30:36:@384.4]
  assign _T_18093 = io_inAddr_18 == 6'h1; // @[Switch.scala 30:53:@386.4]
  assign valid_1_18 = io_inValid_18 & _T_18093; // @[Switch.scala 30:36:@387.4]
  assign _T_18096 = io_inAddr_19 == 6'h1; // @[Switch.scala 30:53:@389.4]
  assign valid_1_19 = io_inValid_19 & _T_18096; // @[Switch.scala 30:36:@390.4]
  assign _T_18099 = io_inAddr_20 == 6'h1; // @[Switch.scala 30:53:@392.4]
  assign valid_1_20 = io_inValid_20 & _T_18099; // @[Switch.scala 30:36:@393.4]
  assign _T_18102 = io_inAddr_21 == 6'h1; // @[Switch.scala 30:53:@395.4]
  assign valid_1_21 = io_inValid_21 & _T_18102; // @[Switch.scala 30:36:@396.4]
  assign _T_18105 = io_inAddr_22 == 6'h1; // @[Switch.scala 30:53:@398.4]
  assign valid_1_22 = io_inValid_22 & _T_18105; // @[Switch.scala 30:36:@399.4]
  assign _T_18108 = io_inAddr_23 == 6'h1; // @[Switch.scala 30:53:@401.4]
  assign valid_1_23 = io_inValid_23 & _T_18108; // @[Switch.scala 30:36:@402.4]
  assign _T_18111 = io_inAddr_24 == 6'h1; // @[Switch.scala 30:53:@404.4]
  assign valid_1_24 = io_inValid_24 & _T_18111; // @[Switch.scala 30:36:@405.4]
  assign _T_18114 = io_inAddr_25 == 6'h1; // @[Switch.scala 30:53:@407.4]
  assign valid_1_25 = io_inValid_25 & _T_18114; // @[Switch.scala 30:36:@408.4]
  assign _T_18117 = io_inAddr_26 == 6'h1; // @[Switch.scala 30:53:@410.4]
  assign valid_1_26 = io_inValid_26 & _T_18117; // @[Switch.scala 30:36:@411.4]
  assign _T_18120 = io_inAddr_27 == 6'h1; // @[Switch.scala 30:53:@413.4]
  assign valid_1_27 = io_inValid_27 & _T_18120; // @[Switch.scala 30:36:@414.4]
  assign _T_18123 = io_inAddr_28 == 6'h1; // @[Switch.scala 30:53:@416.4]
  assign valid_1_28 = io_inValid_28 & _T_18123; // @[Switch.scala 30:36:@417.4]
  assign _T_18126 = io_inAddr_29 == 6'h1; // @[Switch.scala 30:53:@419.4]
  assign valid_1_29 = io_inValid_29 & _T_18126; // @[Switch.scala 30:36:@420.4]
  assign _T_18129 = io_inAddr_30 == 6'h1; // @[Switch.scala 30:53:@422.4]
  assign valid_1_30 = io_inValid_30 & _T_18129; // @[Switch.scala 30:36:@423.4]
  assign _T_18132 = io_inAddr_31 == 6'h1; // @[Switch.scala 30:53:@425.4]
  assign valid_1_31 = io_inValid_31 & _T_18132; // @[Switch.scala 30:36:@426.4]
  assign _T_18135 = io_inAddr_32 == 6'h1; // @[Switch.scala 30:53:@428.4]
  assign valid_1_32 = io_inValid_32 & _T_18135; // @[Switch.scala 30:36:@429.4]
  assign _T_18138 = io_inAddr_33 == 6'h1; // @[Switch.scala 30:53:@431.4]
  assign valid_1_33 = io_inValid_33 & _T_18138; // @[Switch.scala 30:36:@432.4]
  assign _T_18141 = io_inAddr_34 == 6'h1; // @[Switch.scala 30:53:@434.4]
  assign valid_1_34 = io_inValid_34 & _T_18141; // @[Switch.scala 30:36:@435.4]
  assign _T_18144 = io_inAddr_35 == 6'h1; // @[Switch.scala 30:53:@437.4]
  assign valid_1_35 = io_inValid_35 & _T_18144; // @[Switch.scala 30:36:@438.4]
  assign _T_18147 = io_inAddr_36 == 6'h1; // @[Switch.scala 30:53:@440.4]
  assign valid_1_36 = io_inValid_36 & _T_18147; // @[Switch.scala 30:36:@441.4]
  assign _T_18150 = io_inAddr_37 == 6'h1; // @[Switch.scala 30:53:@443.4]
  assign valid_1_37 = io_inValid_37 & _T_18150; // @[Switch.scala 30:36:@444.4]
  assign _T_18153 = io_inAddr_38 == 6'h1; // @[Switch.scala 30:53:@446.4]
  assign valid_1_38 = io_inValid_38 & _T_18153; // @[Switch.scala 30:36:@447.4]
  assign _T_18156 = io_inAddr_39 == 6'h1; // @[Switch.scala 30:53:@449.4]
  assign valid_1_39 = io_inValid_39 & _T_18156; // @[Switch.scala 30:36:@450.4]
  assign _T_18159 = io_inAddr_40 == 6'h1; // @[Switch.scala 30:53:@452.4]
  assign valid_1_40 = io_inValid_40 & _T_18159; // @[Switch.scala 30:36:@453.4]
  assign _T_18162 = io_inAddr_41 == 6'h1; // @[Switch.scala 30:53:@455.4]
  assign valid_1_41 = io_inValid_41 & _T_18162; // @[Switch.scala 30:36:@456.4]
  assign _T_18165 = io_inAddr_42 == 6'h1; // @[Switch.scala 30:53:@458.4]
  assign valid_1_42 = io_inValid_42 & _T_18165; // @[Switch.scala 30:36:@459.4]
  assign _T_18168 = io_inAddr_43 == 6'h1; // @[Switch.scala 30:53:@461.4]
  assign valid_1_43 = io_inValid_43 & _T_18168; // @[Switch.scala 30:36:@462.4]
  assign _T_18171 = io_inAddr_44 == 6'h1; // @[Switch.scala 30:53:@464.4]
  assign valid_1_44 = io_inValid_44 & _T_18171; // @[Switch.scala 30:36:@465.4]
  assign _T_18174 = io_inAddr_45 == 6'h1; // @[Switch.scala 30:53:@467.4]
  assign valid_1_45 = io_inValid_45 & _T_18174; // @[Switch.scala 30:36:@468.4]
  assign _T_18177 = io_inAddr_46 == 6'h1; // @[Switch.scala 30:53:@470.4]
  assign valid_1_46 = io_inValid_46 & _T_18177; // @[Switch.scala 30:36:@471.4]
  assign _T_18180 = io_inAddr_47 == 6'h1; // @[Switch.scala 30:53:@473.4]
  assign valid_1_47 = io_inValid_47 & _T_18180; // @[Switch.scala 30:36:@474.4]
  assign _T_18183 = io_inAddr_48 == 6'h1; // @[Switch.scala 30:53:@476.4]
  assign valid_1_48 = io_inValid_48 & _T_18183; // @[Switch.scala 30:36:@477.4]
  assign _T_18186 = io_inAddr_49 == 6'h1; // @[Switch.scala 30:53:@479.4]
  assign valid_1_49 = io_inValid_49 & _T_18186; // @[Switch.scala 30:36:@480.4]
  assign _T_18189 = io_inAddr_50 == 6'h1; // @[Switch.scala 30:53:@482.4]
  assign valid_1_50 = io_inValid_50 & _T_18189; // @[Switch.scala 30:36:@483.4]
  assign _T_18192 = io_inAddr_51 == 6'h1; // @[Switch.scala 30:53:@485.4]
  assign valid_1_51 = io_inValid_51 & _T_18192; // @[Switch.scala 30:36:@486.4]
  assign _T_18195 = io_inAddr_52 == 6'h1; // @[Switch.scala 30:53:@488.4]
  assign valid_1_52 = io_inValid_52 & _T_18195; // @[Switch.scala 30:36:@489.4]
  assign _T_18198 = io_inAddr_53 == 6'h1; // @[Switch.scala 30:53:@491.4]
  assign valid_1_53 = io_inValid_53 & _T_18198; // @[Switch.scala 30:36:@492.4]
  assign _T_18201 = io_inAddr_54 == 6'h1; // @[Switch.scala 30:53:@494.4]
  assign valid_1_54 = io_inValid_54 & _T_18201; // @[Switch.scala 30:36:@495.4]
  assign _T_18204 = io_inAddr_55 == 6'h1; // @[Switch.scala 30:53:@497.4]
  assign valid_1_55 = io_inValid_55 & _T_18204; // @[Switch.scala 30:36:@498.4]
  assign _T_18207 = io_inAddr_56 == 6'h1; // @[Switch.scala 30:53:@500.4]
  assign valid_1_56 = io_inValid_56 & _T_18207; // @[Switch.scala 30:36:@501.4]
  assign _T_18210 = io_inAddr_57 == 6'h1; // @[Switch.scala 30:53:@503.4]
  assign valid_1_57 = io_inValid_57 & _T_18210; // @[Switch.scala 30:36:@504.4]
  assign _T_18213 = io_inAddr_58 == 6'h1; // @[Switch.scala 30:53:@506.4]
  assign valid_1_58 = io_inValid_58 & _T_18213; // @[Switch.scala 30:36:@507.4]
  assign _T_18216 = io_inAddr_59 == 6'h1; // @[Switch.scala 30:53:@509.4]
  assign valid_1_59 = io_inValid_59 & _T_18216; // @[Switch.scala 30:36:@510.4]
  assign _T_18219 = io_inAddr_60 == 6'h1; // @[Switch.scala 30:53:@512.4]
  assign valid_1_60 = io_inValid_60 & _T_18219; // @[Switch.scala 30:36:@513.4]
  assign _T_18222 = io_inAddr_61 == 6'h1; // @[Switch.scala 30:53:@515.4]
  assign valid_1_61 = io_inValid_61 & _T_18222; // @[Switch.scala 30:36:@516.4]
  assign _T_18225 = io_inAddr_62 == 6'h1; // @[Switch.scala 30:53:@518.4]
  assign valid_1_62 = io_inValid_62 & _T_18225; // @[Switch.scala 30:36:@519.4]
  assign _T_18228 = io_inAddr_63 == 6'h1; // @[Switch.scala 30:53:@521.4]
  assign valid_1_63 = io_inValid_63 & _T_18228; // @[Switch.scala 30:36:@522.4]
  assign _T_18294 = valid_1_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@524.4]
  assign _T_18295 = valid_1_61 ? 6'h3d : _T_18294; // @[Mux.scala 31:69:@525.4]
  assign _T_18296 = valid_1_60 ? 6'h3c : _T_18295; // @[Mux.scala 31:69:@526.4]
  assign _T_18297 = valid_1_59 ? 6'h3b : _T_18296; // @[Mux.scala 31:69:@527.4]
  assign _T_18298 = valid_1_58 ? 6'h3a : _T_18297; // @[Mux.scala 31:69:@528.4]
  assign _T_18299 = valid_1_57 ? 6'h39 : _T_18298; // @[Mux.scala 31:69:@529.4]
  assign _T_18300 = valid_1_56 ? 6'h38 : _T_18299; // @[Mux.scala 31:69:@530.4]
  assign _T_18301 = valid_1_55 ? 6'h37 : _T_18300; // @[Mux.scala 31:69:@531.4]
  assign _T_18302 = valid_1_54 ? 6'h36 : _T_18301; // @[Mux.scala 31:69:@532.4]
  assign _T_18303 = valid_1_53 ? 6'h35 : _T_18302; // @[Mux.scala 31:69:@533.4]
  assign _T_18304 = valid_1_52 ? 6'h34 : _T_18303; // @[Mux.scala 31:69:@534.4]
  assign _T_18305 = valid_1_51 ? 6'h33 : _T_18304; // @[Mux.scala 31:69:@535.4]
  assign _T_18306 = valid_1_50 ? 6'h32 : _T_18305; // @[Mux.scala 31:69:@536.4]
  assign _T_18307 = valid_1_49 ? 6'h31 : _T_18306; // @[Mux.scala 31:69:@537.4]
  assign _T_18308 = valid_1_48 ? 6'h30 : _T_18307; // @[Mux.scala 31:69:@538.4]
  assign _T_18309 = valid_1_47 ? 6'h2f : _T_18308; // @[Mux.scala 31:69:@539.4]
  assign _T_18310 = valid_1_46 ? 6'h2e : _T_18309; // @[Mux.scala 31:69:@540.4]
  assign _T_18311 = valid_1_45 ? 6'h2d : _T_18310; // @[Mux.scala 31:69:@541.4]
  assign _T_18312 = valid_1_44 ? 6'h2c : _T_18311; // @[Mux.scala 31:69:@542.4]
  assign _T_18313 = valid_1_43 ? 6'h2b : _T_18312; // @[Mux.scala 31:69:@543.4]
  assign _T_18314 = valid_1_42 ? 6'h2a : _T_18313; // @[Mux.scala 31:69:@544.4]
  assign _T_18315 = valid_1_41 ? 6'h29 : _T_18314; // @[Mux.scala 31:69:@545.4]
  assign _T_18316 = valid_1_40 ? 6'h28 : _T_18315; // @[Mux.scala 31:69:@546.4]
  assign _T_18317 = valid_1_39 ? 6'h27 : _T_18316; // @[Mux.scala 31:69:@547.4]
  assign _T_18318 = valid_1_38 ? 6'h26 : _T_18317; // @[Mux.scala 31:69:@548.4]
  assign _T_18319 = valid_1_37 ? 6'h25 : _T_18318; // @[Mux.scala 31:69:@549.4]
  assign _T_18320 = valid_1_36 ? 6'h24 : _T_18319; // @[Mux.scala 31:69:@550.4]
  assign _T_18321 = valid_1_35 ? 6'h23 : _T_18320; // @[Mux.scala 31:69:@551.4]
  assign _T_18322 = valid_1_34 ? 6'h22 : _T_18321; // @[Mux.scala 31:69:@552.4]
  assign _T_18323 = valid_1_33 ? 6'h21 : _T_18322; // @[Mux.scala 31:69:@553.4]
  assign _T_18324 = valid_1_32 ? 6'h20 : _T_18323; // @[Mux.scala 31:69:@554.4]
  assign _T_18325 = valid_1_31 ? 6'h1f : _T_18324; // @[Mux.scala 31:69:@555.4]
  assign _T_18326 = valid_1_30 ? 6'h1e : _T_18325; // @[Mux.scala 31:69:@556.4]
  assign _T_18327 = valid_1_29 ? 6'h1d : _T_18326; // @[Mux.scala 31:69:@557.4]
  assign _T_18328 = valid_1_28 ? 6'h1c : _T_18327; // @[Mux.scala 31:69:@558.4]
  assign _T_18329 = valid_1_27 ? 6'h1b : _T_18328; // @[Mux.scala 31:69:@559.4]
  assign _T_18330 = valid_1_26 ? 6'h1a : _T_18329; // @[Mux.scala 31:69:@560.4]
  assign _T_18331 = valid_1_25 ? 6'h19 : _T_18330; // @[Mux.scala 31:69:@561.4]
  assign _T_18332 = valid_1_24 ? 6'h18 : _T_18331; // @[Mux.scala 31:69:@562.4]
  assign _T_18333 = valid_1_23 ? 6'h17 : _T_18332; // @[Mux.scala 31:69:@563.4]
  assign _T_18334 = valid_1_22 ? 6'h16 : _T_18333; // @[Mux.scala 31:69:@564.4]
  assign _T_18335 = valid_1_21 ? 6'h15 : _T_18334; // @[Mux.scala 31:69:@565.4]
  assign _T_18336 = valid_1_20 ? 6'h14 : _T_18335; // @[Mux.scala 31:69:@566.4]
  assign _T_18337 = valid_1_19 ? 6'h13 : _T_18336; // @[Mux.scala 31:69:@567.4]
  assign _T_18338 = valid_1_18 ? 6'h12 : _T_18337; // @[Mux.scala 31:69:@568.4]
  assign _T_18339 = valid_1_17 ? 6'h11 : _T_18338; // @[Mux.scala 31:69:@569.4]
  assign _T_18340 = valid_1_16 ? 6'h10 : _T_18339; // @[Mux.scala 31:69:@570.4]
  assign _T_18341 = valid_1_15 ? 6'hf : _T_18340; // @[Mux.scala 31:69:@571.4]
  assign _T_18342 = valid_1_14 ? 6'he : _T_18341; // @[Mux.scala 31:69:@572.4]
  assign _T_18343 = valid_1_13 ? 6'hd : _T_18342; // @[Mux.scala 31:69:@573.4]
  assign _T_18344 = valid_1_12 ? 6'hc : _T_18343; // @[Mux.scala 31:69:@574.4]
  assign _T_18345 = valid_1_11 ? 6'hb : _T_18344; // @[Mux.scala 31:69:@575.4]
  assign _T_18346 = valid_1_10 ? 6'ha : _T_18345; // @[Mux.scala 31:69:@576.4]
  assign _T_18347 = valid_1_9 ? 6'h9 : _T_18346; // @[Mux.scala 31:69:@577.4]
  assign _T_18348 = valid_1_8 ? 6'h8 : _T_18347; // @[Mux.scala 31:69:@578.4]
  assign _T_18349 = valid_1_7 ? 6'h7 : _T_18348; // @[Mux.scala 31:69:@579.4]
  assign _T_18350 = valid_1_6 ? 6'h6 : _T_18349; // @[Mux.scala 31:69:@580.4]
  assign _T_18351 = valid_1_5 ? 6'h5 : _T_18350; // @[Mux.scala 31:69:@581.4]
  assign _T_18352 = valid_1_4 ? 6'h4 : _T_18351; // @[Mux.scala 31:69:@582.4]
  assign _T_18353 = valid_1_3 ? 6'h3 : _T_18352; // @[Mux.scala 31:69:@583.4]
  assign _T_18354 = valid_1_2 ? 6'h2 : _T_18353; // @[Mux.scala 31:69:@584.4]
  assign _T_18355 = valid_1_1 ? 6'h1 : _T_18354; // @[Mux.scala 31:69:@585.4]
  assign select_1 = valid_1_0 ? 6'h0 : _T_18355; // @[Mux.scala 31:69:@586.4]
  assign _GEN_65 = 6'h1 == select_1 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@588.4]
  assign _GEN_66 = 6'h2 == select_1 ? io_inData_2 : _GEN_65; // @[Switch.scala 33:19:@588.4]
  assign _GEN_67 = 6'h3 == select_1 ? io_inData_3 : _GEN_66; // @[Switch.scala 33:19:@588.4]
  assign _GEN_68 = 6'h4 == select_1 ? io_inData_4 : _GEN_67; // @[Switch.scala 33:19:@588.4]
  assign _GEN_69 = 6'h5 == select_1 ? io_inData_5 : _GEN_68; // @[Switch.scala 33:19:@588.4]
  assign _GEN_70 = 6'h6 == select_1 ? io_inData_6 : _GEN_69; // @[Switch.scala 33:19:@588.4]
  assign _GEN_71 = 6'h7 == select_1 ? io_inData_7 : _GEN_70; // @[Switch.scala 33:19:@588.4]
  assign _GEN_72 = 6'h8 == select_1 ? io_inData_8 : _GEN_71; // @[Switch.scala 33:19:@588.4]
  assign _GEN_73 = 6'h9 == select_1 ? io_inData_9 : _GEN_72; // @[Switch.scala 33:19:@588.4]
  assign _GEN_74 = 6'ha == select_1 ? io_inData_10 : _GEN_73; // @[Switch.scala 33:19:@588.4]
  assign _GEN_75 = 6'hb == select_1 ? io_inData_11 : _GEN_74; // @[Switch.scala 33:19:@588.4]
  assign _GEN_76 = 6'hc == select_1 ? io_inData_12 : _GEN_75; // @[Switch.scala 33:19:@588.4]
  assign _GEN_77 = 6'hd == select_1 ? io_inData_13 : _GEN_76; // @[Switch.scala 33:19:@588.4]
  assign _GEN_78 = 6'he == select_1 ? io_inData_14 : _GEN_77; // @[Switch.scala 33:19:@588.4]
  assign _GEN_79 = 6'hf == select_1 ? io_inData_15 : _GEN_78; // @[Switch.scala 33:19:@588.4]
  assign _GEN_80 = 6'h10 == select_1 ? io_inData_16 : _GEN_79; // @[Switch.scala 33:19:@588.4]
  assign _GEN_81 = 6'h11 == select_1 ? io_inData_17 : _GEN_80; // @[Switch.scala 33:19:@588.4]
  assign _GEN_82 = 6'h12 == select_1 ? io_inData_18 : _GEN_81; // @[Switch.scala 33:19:@588.4]
  assign _GEN_83 = 6'h13 == select_1 ? io_inData_19 : _GEN_82; // @[Switch.scala 33:19:@588.4]
  assign _GEN_84 = 6'h14 == select_1 ? io_inData_20 : _GEN_83; // @[Switch.scala 33:19:@588.4]
  assign _GEN_85 = 6'h15 == select_1 ? io_inData_21 : _GEN_84; // @[Switch.scala 33:19:@588.4]
  assign _GEN_86 = 6'h16 == select_1 ? io_inData_22 : _GEN_85; // @[Switch.scala 33:19:@588.4]
  assign _GEN_87 = 6'h17 == select_1 ? io_inData_23 : _GEN_86; // @[Switch.scala 33:19:@588.4]
  assign _GEN_88 = 6'h18 == select_1 ? io_inData_24 : _GEN_87; // @[Switch.scala 33:19:@588.4]
  assign _GEN_89 = 6'h19 == select_1 ? io_inData_25 : _GEN_88; // @[Switch.scala 33:19:@588.4]
  assign _GEN_90 = 6'h1a == select_1 ? io_inData_26 : _GEN_89; // @[Switch.scala 33:19:@588.4]
  assign _GEN_91 = 6'h1b == select_1 ? io_inData_27 : _GEN_90; // @[Switch.scala 33:19:@588.4]
  assign _GEN_92 = 6'h1c == select_1 ? io_inData_28 : _GEN_91; // @[Switch.scala 33:19:@588.4]
  assign _GEN_93 = 6'h1d == select_1 ? io_inData_29 : _GEN_92; // @[Switch.scala 33:19:@588.4]
  assign _GEN_94 = 6'h1e == select_1 ? io_inData_30 : _GEN_93; // @[Switch.scala 33:19:@588.4]
  assign _GEN_95 = 6'h1f == select_1 ? io_inData_31 : _GEN_94; // @[Switch.scala 33:19:@588.4]
  assign _GEN_96 = 6'h20 == select_1 ? io_inData_32 : _GEN_95; // @[Switch.scala 33:19:@588.4]
  assign _GEN_97 = 6'h21 == select_1 ? io_inData_33 : _GEN_96; // @[Switch.scala 33:19:@588.4]
  assign _GEN_98 = 6'h22 == select_1 ? io_inData_34 : _GEN_97; // @[Switch.scala 33:19:@588.4]
  assign _GEN_99 = 6'h23 == select_1 ? io_inData_35 : _GEN_98; // @[Switch.scala 33:19:@588.4]
  assign _GEN_100 = 6'h24 == select_1 ? io_inData_36 : _GEN_99; // @[Switch.scala 33:19:@588.4]
  assign _GEN_101 = 6'h25 == select_1 ? io_inData_37 : _GEN_100; // @[Switch.scala 33:19:@588.4]
  assign _GEN_102 = 6'h26 == select_1 ? io_inData_38 : _GEN_101; // @[Switch.scala 33:19:@588.4]
  assign _GEN_103 = 6'h27 == select_1 ? io_inData_39 : _GEN_102; // @[Switch.scala 33:19:@588.4]
  assign _GEN_104 = 6'h28 == select_1 ? io_inData_40 : _GEN_103; // @[Switch.scala 33:19:@588.4]
  assign _GEN_105 = 6'h29 == select_1 ? io_inData_41 : _GEN_104; // @[Switch.scala 33:19:@588.4]
  assign _GEN_106 = 6'h2a == select_1 ? io_inData_42 : _GEN_105; // @[Switch.scala 33:19:@588.4]
  assign _GEN_107 = 6'h2b == select_1 ? io_inData_43 : _GEN_106; // @[Switch.scala 33:19:@588.4]
  assign _GEN_108 = 6'h2c == select_1 ? io_inData_44 : _GEN_107; // @[Switch.scala 33:19:@588.4]
  assign _GEN_109 = 6'h2d == select_1 ? io_inData_45 : _GEN_108; // @[Switch.scala 33:19:@588.4]
  assign _GEN_110 = 6'h2e == select_1 ? io_inData_46 : _GEN_109; // @[Switch.scala 33:19:@588.4]
  assign _GEN_111 = 6'h2f == select_1 ? io_inData_47 : _GEN_110; // @[Switch.scala 33:19:@588.4]
  assign _GEN_112 = 6'h30 == select_1 ? io_inData_48 : _GEN_111; // @[Switch.scala 33:19:@588.4]
  assign _GEN_113 = 6'h31 == select_1 ? io_inData_49 : _GEN_112; // @[Switch.scala 33:19:@588.4]
  assign _GEN_114 = 6'h32 == select_1 ? io_inData_50 : _GEN_113; // @[Switch.scala 33:19:@588.4]
  assign _GEN_115 = 6'h33 == select_1 ? io_inData_51 : _GEN_114; // @[Switch.scala 33:19:@588.4]
  assign _GEN_116 = 6'h34 == select_1 ? io_inData_52 : _GEN_115; // @[Switch.scala 33:19:@588.4]
  assign _GEN_117 = 6'h35 == select_1 ? io_inData_53 : _GEN_116; // @[Switch.scala 33:19:@588.4]
  assign _GEN_118 = 6'h36 == select_1 ? io_inData_54 : _GEN_117; // @[Switch.scala 33:19:@588.4]
  assign _GEN_119 = 6'h37 == select_1 ? io_inData_55 : _GEN_118; // @[Switch.scala 33:19:@588.4]
  assign _GEN_120 = 6'h38 == select_1 ? io_inData_56 : _GEN_119; // @[Switch.scala 33:19:@588.4]
  assign _GEN_121 = 6'h39 == select_1 ? io_inData_57 : _GEN_120; // @[Switch.scala 33:19:@588.4]
  assign _GEN_122 = 6'h3a == select_1 ? io_inData_58 : _GEN_121; // @[Switch.scala 33:19:@588.4]
  assign _GEN_123 = 6'h3b == select_1 ? io_inData_59 : _GEN_122; // @[Switch.scala 33:19:@588.4]
  assign _GEN_124 = 6'h3c == select_1 ? io_inData_60 : _GEN_123; // @[Switch.scala 33:19:@588.4]
  assign _GEN_125 = 6'h3d == select_1 ? io_inData_61 : _GEN_124; // @[Switch.scala 33:19:@588.4]
  assign _GEN_126 = 6'h3e == select_1 ? io_inData_62 : _GEN_125; // @[Switch.scala 33:19:@588.4]
  assign _T_18364 = {valid_1_7,valid_1_6,valid_1_5,valid_1_4,valid_1_3,valid_1_2,valid_1_1,valid_1_0}; // @[Switch.scala 34:32:@595.4]
  assign _T_18372 = {valid_1_15,valid_1_14,valid_1_13,valid_1_12,valid_1_11,valid_1_10,valid_1_9,valid_1_8,_T_18364}; // @[Switch.scala 34:32:@603.4]
  assign _T_18379 = {valid_1_23,valid_1_22,valid_1_21,valid_1_20,valid_1_19,valid_1_18,valid_1_17,valid_1_16}; // @[Switch.scala 34:32:@610.4]
  assign _T_18388 = {valid_1_31,valid_1_30,valid_1_29,valid_1_28,valid_1_27,valid_1_26,valid_1_25,valid_1_24,_T_18379,_T_18372}; // @[Switch.scala 34:32:@619.4]
  assign _T_18395 = {valid_1_39,valid_1_38,valid_1_37,valid_1_36,valid_1_35,valid_1_34,valid_1_33,valid_1_32}; // @[Switch.scala 34:32:@626.4]
  assign _T_18403 = {valid_1_47,valid_1_46,valid_1_45,valid_1_44,valid_1_43,valid_1_42,valid_1_41,valid_1_40,_T_18395}; // @[Switch.scala 34:32:@634.4]
  assign _T_18410 = {valid_1_55,valid_1_54,valid_1_53,valid_1_52,valid_1_51,valid_1_50,valid_1_49,valid_1_48}; // @[Switch.scala 34:32:@641.4]
  assign _T_18419 = {valid_1_63,valid_1_62,valid_1_61,valid_1_60,valid_1_59,valid_1_58,valid_1_57,valid_1_56,_T_18410,_T_18403}; // @[Switch.scala 34:32:@650.4]
  assign _T_18420 = {_T_18419,_T_18388}; // @[Switch.scala 34:32:@651.4]
  assign _T_18424 = io_inAddr_0 == 6'h2; // @[Switch.scala 30:53:@654.4]
  assign valid_2_0 = io_inValid_0 & _T_18424; // @[Switch.scala 30:36:@655.4]
  assign _T_18427 = io_inAddr_1 == 6'h2; // @[Switch.scala 30:53:@657.4]
  assign valid_2_1 = io_inValid_1 & _T_18427; // @[Switch.scala 30:36:@658.4]
  assign _T_18430 = io_inAddr_2 == 6'h2; // @[Switch.scala 30:53:@660.4]
  assign valid_2_2 = io_inValid_2 & _T_18430; // @[Switch.scala 30:36:@661.4]
  assign _T_18433 = io_inAddr_3 == 6'h2; // @[Switch.scala 30:53:@663.4]
  assign valid_2_3 = io_inValid_3 & _T_18433; // @[Switch.scala 30:36:@664.4]
  assign _T_18436 = io_inAddr_4 == 6'h2; // @[Switch.scala 30:53:@666.4]
  assign valid_2_4 = io_inValid_4 & _T_18436; // @[Switch.scala 30:36:@667.4]
  assign _T_18439 = io_inAddr_5 == 6'h2; // @[Switch.scala 30:53:@669.4]
  assign valid_2_5 = io_inValid_5 & _T_18439; // @[Switch.scala 30:36:@670.4]
  assign _T_18442 = io_inAddr_6 == 6'h2; // @[Switch.scala 30:53:@672.4]
  assign valid_2_6 = io_inValid_6 & _T_18442; // @[Switch.scala 30:36:@673.4]
  assign _T_18445 = io_inAddr_7 == 6'h2; // @[Switch.scala 30:53:@675.4]
  assign valid_2_7 = io_inValid_7 & _T_18445; // @[Switch.scala 30:36:@676.4]
  assign _T_18448 = io_inAddr_8 == 6'h2; // @[Switch.scala 30:53:@678.4]
  assign valid_2_8 = io_inValid_8 & _T_18448; // @[Switch.scala 30:36:@679.4]
  assign _T_18451 = io_inAddr_9 == 6'h2; // @[Switch.scala 30:53:@681.4]
  assign valid_2_9 = io_inValid_9 & _T_18451; // @[Switch.scala 30:36:@682.4]
  assign _T_18454 = io_inAddr_10 == 6'h2; // @[Switch.scala 30:53:@684.4]
  assign valid_2_10 = io_inValid_10 & _T_18454; // @[Switch.scala 30:36:@685.4]
  assign _T_18457 = io_inAddr_11 == 6'h2; // @[Switch.scala 30:53:@687.4]
  assign valid_2_11 = io_inValid_11 & _T_18457; // @[Switch.scala 30:36:@688.4]
  assign _T_18460 = io_inAddr_12 == 6'h2; // @[Switch.scala 30:53:@690.4]
  assign valid_2_12 = io_inValid_12 & _T_18460; // @[Switch.scala 30:36:@691.4]
  assign _T_18463 = io_inAddr_13 == 6'h2; // @[Switch.scala 30:53:@693.4]
  assign valid_2_13 = io_inValid_13 & _T_18463; // @[Switch.scala 30:36:@694.4]
  assign _T_18466 = io_inAddr_14 == 6'h2; // @[Switch.scala 30:53:@696.4]
  assign valid_2_14 = io_inValid_14 & _T_18466; // @[Switch.scala 30:36:@697.4]
  assign _T_18469 = io_inAddr_15 == 6'h2; // @[Switch.scala 30:53:@699.4]
  assign valid_2_15 = io_inValid_15 & _T_18469; // @[Switch.scala 30:36:@700.4]
  assign _T_18472 = io_inAddr_16 == 6'h2; // @[Switch.scala 30:53:@702.4]
  assign valid_2_16 = io_inValid_16 & _T_18472; // @[Switch.scala 30:36:@703.4]
  assign _T_18475 = io_inAddr_17 == 6'h2; // @[Switch.scala 30:53:@705.4]
  assign valid_2_17 = io_inValid_17 & _T_18475; // @[Switch.scala 30:36:@706.4]
  assign _T_18478 = io_inAddr_18 == 6'h2; // @[Switch.scala 30:53:@708.4]
  assign valid_2_18 = io_inValid_18 & _T_18478; // @[Switch.scala 30:36:@709.4]
  assign _T_18481 = io_inAddr_19 == 6'h2; // @[Switch.scala 30:53:@711.4]
  assign valid_2_19 = io_inValid_19 & _T_18481; // @[Switch.scala 30:36:@712.4]
  assign _T_18484 = io_inAddr_20 == 6'h2; // @[Switch.scala 30:53:@714.4]
  assign valid_2_20 = io_inValid_20 & _T_18484; // @[Switch.scala 30:36:@715.4]
  assign _T_18487 = io_inAddr_21 == 6'h2; // @[Switch.scala 30:53:@717.4]
  assign valid_2_21 = io_inValid_21 & _T_18487; // @[Switch.scala 30:36:@718.4]
  assign _T_18490 = io_inAddr_22 == 6'h2; // @[Switch.scala 30:53:@720.4]
  assign valid_2_22 = io_inValid_22 & _T_18490; // @[Switch.scala 30:36:@721.4]
  assign _T_18493 = io_inAddr_23 == 6'h2; // @[Switch.scala 30:53:@723.4]
  assign valid_2_23 = io_inValid_23 & _T_18493; // @[Switch.scala 30:36:@724.4]
  assign _T_18496 = io_inAddr_24 == 6'h2; // @[Switch.scala 30:53:@726.4]
  assign valid_2_24 = io_inValid_24 & _T_18496; // @[Switch.scala 30:36:@727.4]
  assign _T_18499 = io_inAddr_25 == 6'h2; // @[Switch.scala 30:53:@729.4]
  assign valid_2_25 = io_inValid_25 & _T_18499; // @[Switch.scala 30:36:@730.4]
  assign _T_18502 = io_inAddr_26 == 6'h2; // @[Switch.scala 30:53:@732.4]
  assign valid_2_26 = io_inValid_26 & _T_18502; // @[Switch.scala 30:36:@733.4]
  assign _T_18505 = io_inAddr_27 == 6'h2; // @[Switch.scala 30:53:@735.4]
  assign valid_2_27 = io_inValid_27 & _T_18505; // @[Switch.scala 30:36:@736.4]
  assign _T_18508 = io_inAddr_28 == 6'h2; // @[Switch.scala 30:53:@738.4]
  assign valid_2_28 = io_inValid_28 & _T_18508; // @[Switch.scala 30:36:@739.4]
  assign _T_18511 = io_inAddr_29 == 6'h2; // @[Switch.scala 30:53:@741.4]
  assign valid_2_29 = io_inValid_29 & _T_18511; // @[Switch.scala 30:36:@742.4]
  assign _T_18514 = io_inAddr_30 == 6'h2; // @[Switch.scala 30:53:@744.4]
  assign valid_2_30 = io_inValid_30 & _T_18514; // @[Switch.scala 30:36:@745.4]
  assign _T_18517 = io_inAddr_31 == 6'h2; // @[Switch.scala 30:53:@747.4]
  assign valid_2_31 = io_inValid_31 & _T_18517; // @[Switch.scala 30:36:@748.4]
  assign _T_18520 = io_inAddr_32 == 6'h2; // @[Switch.scala 30:53:@750.4]
  assign valid_2_32 = io_inValid_32 & _T_18520; // @[Switch.scala 30:36:@751.4]
  assign _T_18523 = io_inAddr_33 == 6'h2; // @[Switch.scala 30:53:@753.4]
  assign valid_2_33 = io_inValid_33 & _T_18523; // @[Switch.scala 30:36:@754.4]
  assign _T_18526 = io_inAddr_34 == 6'h2; // @[Switch.scala 30:53:@756.4]
  assign valid_2_34 = io_inValid_34 & _T_18526; // @[Switch.scala 30:36:@757.4]
  assign _T_18529 = io_inAddr_35 == 6'h2; // @[Switch.scala 30:53:@759.4]
  assign valid_2_35 = io_inValid_35 & _T_18529; // @[Switch.scala 30:36:@760.4]
  assign _T_18532 = io_inAddr_36 == 6'h2; // @[Switch.scala 30:53:@762.4]
  assign valid_2_36 = io_inValid_36 & _T_18532; // @[Switch.scala 30:36:@763.4]
  assign _T_18535 = io_inAddr_37 == 6'h2; // @[Switch.scala 30:53:@765.4]
  assign valid_2_37 = io_inValid_37 & _T_18535; // @[Switch.scala 30:36:@766.4]
  assign _T_18538 = io_inAddr_38 == 6'h2; // @[Switch.scala 30:53:@768.4]
  assign valid_2_38 = io_inValid_38 & _T_18538; // @[Switch.scala 30:36:@769.4]
  assign _T_18541 = io_inAddr_39 == 6'h2; // @[Switch.scala 30:53:@771.4]
  assign valid_2_39 = io_inValid_39 & _T_18541; // @[Switch.scala 30:36:@772.4]
  assign _T_18544 = io_inAddr_40 == 6'h2; // @[Switch.scala 30:53:@774.4]
  assign valid_2_40 = io_inValid_40 & _T_18544; // @[Switch.scala 30:36:@775.4]
  assign _T_18547 = io_inAddr_41 == 6'h2; // @[Switch.scala 30:53:@777.4]
  assign valid_2_41 = io_inValid_41 & _T_18547; // @[Switch.scala 30:36:@778.4]
  assign _T_18550 = io_inAddr_42 == 6'h2; // @[Switch.scala 30:53:@780.4]
  assign valid_2_42 = io_inValid_42 & _T_18550; // @[Switch.scala 30:36:@781.4]
  assign _T_18553 = io_inAddr_43 == 6'h2; // @[Switch.scala 30:53:@783.4]
  assign valid_2_43 = io_inValid_43 & _T_18553; // @[Switch.scala 30:36:@784.4]
  assign _T_18556 = io_inAddr_44 == 6'h2; // @[Switch.scala 30:53:@786.4]
  assign valid_2_44 = io_inValid_44 & _T_18556; // @[Switch.scala 30:36:@787.4]
  assign _T_18559 = io_inAddr_45 == 6'h2; // @[Switch.scala 30:53:@789.4]
  assign valid_2_45 = io_inValid_45 & _T_18559; // @[Switch.scala 30:36:@790.4]
  assign _T_18562 = io_inAddr_46 == 6'h2; // @[Switch.scala 30:53:@792.4]
  assign valid_2_46 = io_inValid_46 & _T_18562; // @[Switch.scala 30:36:@793.4]
  assign _T_18565 = io_inAddr_47 == 6'h2; // @[Switch.scala 30:53:@795.4]
  assign valid_2_47 = io_inValid_47 & _T_18565; // @[Switch.scala 30:36:@796.4]
  assign _T_18568 = io_inAddr_48 == 6'h2; // @[Switch.scala 30:53:@798.4]
  assign valid_2_48 = io_inValid_48 & _T_18568; // @[Switch.scala 30:36:@799.4]
  assign _T_18571 = io_inAddr_49 == 6'h2; // @[Switch.scala 30:53:@801.4]
  assign valid_2_49 = io_inValid_49 & _T_18571; // @[Switch.scala 30:36:@802.4]
  assign _T_18574 = io_inAddr_50 == 6'h2; // @[Switch.scala 30:53:@804.4]
  assign valid_2_50 = io_inValid_50 & _T_18574; // @[Switch.scala 30:36:@805.4]
  assign _T_18577 = io_inAddr_51 == 6'h2; // @[Switch.scala 30:53:@807.4]
  assign valid_2_51 = io_inValid_51 & _T_18577; // @[Switch.scala 30:36:@808.4]
  assign _T_18580 = io_inAddr_52 == 6'h2; // @[Switch.scala 30:53:@810.4]
  assign valid_2_52 = io_inValid_52 & _T_18580; // @[Switch.scala 30:36:@811.4]
  assign _T_18583 = io_inAddr_53 == 6'h2; // @[Switch.scala 30:53:@813.4]
  assign valid_2_53 = io_inValid_53 & _T_18583; // @[Switch.scala 30:36:@814.4]
  assign _T_18586 = io_inAddr_54 == 6'h2; // @[Switch.scala 30:53:@816.4]
  assign valid_2_54 = io_inValid_54 & _T_18586; // @[Switch.scala 30:36:@817.4]
  assign _T_18589 = io_inAddr_55 == 6'h2; // @[Switch.scala 30:53:@819.4]
  assign valid_2_55 = io_inValid_55 & _T_18589; // @[Switch.scala 30:36:@820.4]
  assign _T_18592 = io_inAddr_56 == 6'h2; // @[Switch.scala 30:53:@822.4]
  assign valid_2_56 = io_inValid_56 & _T_18592; // @[Switch.scala 30:36:@823.4]
  assign _T_18595 = io_inAddr_57 == 6'h2; // @[Switch.scala 30:53:@825.4]
  assign valid_2_57 = io_inValid_57 & _T_18595; // @[Switch.scala 30:36:@826.4]
  assign _T_18598 = io_inAddr_58 == 6'h2; // @[Switch.scala 30:53:@828.4]
  assign valid_2_58 = io_inValid_58 & _T_18598; // @[Switch.scala 30:36:@829.4]
  assign _T_18601 = io_inAddr_59 == 6'h2; // @[Switch.scala 30:53:@831.4]
  assign valid_2_59 = io_inValid_59 & _T_18601; // @[Switch.scala 30:36:@832.4]
  assign _T_18604 = io_inAddr_60 == 6'h2; // @[Switch.scala 30:53:@834.4]
  assign valid_2_60 = io_inValid_60 & _T_18604; // @[Switch.scala 30:36:@835.4]
  assign _T_18607 = io_inAddr_61 == 6'h2; // @[Switch.scala 30:53:@837.4]
  assign valid_2_61 = io_inValid_61 & _T_18607; // @[Switch.scala 30:36:@838.4]
  assign _T_18610 = io_inAddr_62 == 6'h2; // @[Switch.scala 30:53:@840.4]
  assign valid_2_62 = io_inValid_62 & _T_18610; // @[Switch.scala 30:36:@841.4]
  assign _T_18613 = io_inAddr_63 == 6'h2; // @[Switch.scala 30:53:@843.4]
  assign valid_2_63 = io_inValid_63 & _T_18613; // @[Switch.scala 30:36:@844.4]
  assign _T_18679 = valid_2_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@846.4]
  assign _T_18680 = valid_2_61 ? 6'h3d : _T_18679; // @[Mux.scala 31:69:@847.4]
  assign _T_18681 = valid_2_60 ? 6'h3c : _T_18680; // @[Mux.scala 31:69:@848.4]
  assign _T_18682 = valid_2_59 ? 6'h3b : _T_18681; // @[Mux.scala 31:69:@849.4]
  assign _T_18683 = valid_2_58 ? 6'h3a : _T_18682; // @[Mux.scala 31:69:@850.4]
  assign _T_18684 = valid_2_57 ? 6'h39 : _T_18683; // @[Mux.scala 31:69:@851.4]
  assign _T_18685 = valid_2_56 ? 6'h38 : _T_18684; // @[Mux.scala 31:69:@852.4]
  assign _T_18686 = valid_2_55 ? 6'h37 : _T_18685; // @[Mux.scala 31:69:@853.4]
  assign _T_18687 = valid_2_54 ? 6'h36 : _T_18686; // @[Mux.scala 31:69:@854.4]
  assign _T_18688 = valid_2_53 ? 6'h35 : _T_18687; // @[Mux.scala 31:69:@855.4]
  assign _T_18689 = valid_2_52 ? 6'h34 : _T_18688; // @[Mux.scala 31:69:@856.4]
  assign _T_18690 = valid_2_51 ? 6'h33 : _T_18689; // @[Mux.scala 31:69:@857.4]
  assign _T_18691 = valid_2_50 ? 6'h32 : _T_18690; // @[Mux.scala 31:69:@858.4]
  assign _T_18692 = valid_2_49 ? 6'h31 : _T_18691; // @[Mux.scala 31:69:@859.4]
  assign _T_18693 = valid_2_48 ? 6'h30 : _T_18692; // @[Mux.scala 31:69:@860.4]
  assign _T_18694 = valid_2_47 ? 6'h2f : _T_18693; // @[Mux.scala 31:69:@861.4]
  assign _T_18695 = valid_2_46 ? 6'h2e : _T_18694; // @[Mux.scala 31:69:@862.4]
  assign _T_18696 = valid_2_45 ? 6'h2d : _T_18695; // @[Mux.scala 31:69:@863.4]
  assign _T_18697 = valid_2_44 ? 6'h2c : _T_18696; // @[Mux.scala 31:69:@864.4]
  assign _T_18698 = valid_2_43 ? 6'h2b : _T_18697; // @[Mux.scala 31:69:@865.4]
  assign _T_18699 = valid_2_42 ? 6'h2a : _T_18698; // @[Mux.scala 31:69:@866.4]
  assign _T_18700 = valid_2_41 ? 6'h29 : _T_18699; // @[Mux.scala 31:69:@867.4]
  assign _T_18701 = valid_2_40 ? 6'h28 : _T_18700; // @[Mux.scala 31:69:@868.4]
  assign _T_18702 = valid_2_39 ? 6'h27 : _T_18701; // @[Mux.scala 31:69:@869.4]
  assign _T_18703 = valid_2_38 ? 6'h26 : _T_18702; // @[Mux.scala 31:69:@870.4]
  assign _T_18704 = valid_2_37 ? 6'h25 : _T_18703; // @[Mux.scala 31:69:@871.4]
  assign _T_18705 = valid_2_36 ? 6'h24 : _T_18704; // @[Mux.scala 31:69:@872.4]
  assign _T_18706 = valid_2_35 ? 6'h23 : _T_18705; // @[Mux.scala 31:69:@873.4]
  assign _T_18707 = valid_2_34 ? 6'h22 : _T_18706; // @[Mux.scala 31:69:@874.4]
  assign _T_18708 = valid_2_33 ? 6'h21 : _T_18707; // @[Mux.scala 31:69:@875.4]
  assign _T_18709 = valid_2_32 ? 6'h20 : _T_18708; // @[Mux.scala 31:69:@876.4]
  assign _T_18710 = valid_2_31 ? 6'h1f : _T_18709; // @[Mux.scala 31:69:@877.4]
  assign _T_18711 = valid_2_30 ? 6'h1e : _T_18710; // @[Mux.scala 31:69:@878.4]
  assign _T_18712 = valid_2_29 ? 6'h1d : _T_18711; // @[Mux.scala 31:69:@879.4]
  assign _T_18713 = valid_2_28 ? 6'h1c : _T_18712; // @[Mux.scala 31:69:@880.4]
  assign _T_18714 = valid_2_27 ? 6'h1b : _T_18713; // @[Mux.scala 31:69:@881.4]
  assign _T_18715 = valid_2_26 ? 6'h1a : _T_18714; // @[Mux.scala 31:69:@882.4]
  assign _T_18716 = valid_2_25 ? 6'h19 : _T_18715; // @[Mux.scala 31:69:@883.4]
  assign _T_18717 = valid_2_24 ? 6'h18 : _T_18716; // @[Mux.scala 31:69:@884.4]
  assign _T_18718 = valid_2_23 ? 6'h17 : _T_18717; // @[Mux.scala 31:69:@885.4]
  assign _T_18719 = valid_2_22 ? 6'h16 : _T_18718; // @[Mux.scala 31:69:@886.4]
  assign _T_18720 = valid_2_21 ? 6'h15 : _T_18719; // @[Mux.scala 31:69:@887.4]
  assign _T_18721 = valid_2_20 ? 6'h14 : _T_18720; // @[Mux.scala 31:69:@888.4]
  assign _T_18722 = valid_2_19 ? 6'h13 : _T_18721; // @[Mux.scala 31:69:@889.4]
  assign _T_18723 = valid_2_18 ? 6'h12 : _T_18722; // @[Mux.scala 31:69:@890.4]
  assign _T_18724 = valid_2_17 ? 6'h11 : _T_18723; // @[Mux.scala 31:69:@891.4]
  assign _T_18725 = valid_2_16 ? 6'h10 : _T_18724; // @[Mux.scala 31:69:@892.4]
  assign _T_18726 = valid_2_15 ? 6'hf : _T_18725; // @[Mux.scala 31:69:@893.4]
  assign _T_18727 = valid_2_14 ? 6'he : _T_18726; // @[Mux.scala 31:69:@894.4]
  assign _T_18728 = valid_2_13 ? 6'hd : _T_18727; // @[Mux.scala 31:69:@895.4]
  assign _T_18729 = valid_2_12 ? 6'hc : _T_18728; // @[Mux.scala 31:69:@896.4]
  assign _T_18730 = valid_2_11 ? 6'hb : _T_18729; // @[Mux.scala 31:69:@897.4]
  assign _T_18731 = valid_2_10 ? 6'ha : _T_18730; // @[Mux.scala 31:69:@898.4]
  assign _T_18732 = valid_2_9 ? 6'h9 : _T_18731; // @[Mux.scala 31:69:@899.4]
  assign _T_18733 = valid_2_8 ? 6'h8 : _T_18732; // @[Mux.scala 31:69:@900.4]
  assign _T_18734 = valid_2_7 ? 6'h7 : _T_18733; // @[Mux.scala 31:69:@901.4]
  assign _T_18735 = valid_2_6 ? 6'h6 : _T_18734; // @[Mux.scala 31:69:@902.4]
  assign _T_18736 = valid_2_5 ? 6'h5 : _T_18735; // @[Mux.scala 31:69:@903.4]
  assign _T_18737 = valid_2_4 ? 6'h4 : _T_18736; // @[Mux.scala 31:69:@904.4]
  assign _T_18738 = valid_2_3 ? 6'h3 : _T_18737; // @[Mux.scala 31:69:@905.4]
  assign _T_18739 = valid_2_2 ? 6'h2 : _T_18738; // @[Mux.scala 31:69:@906.4]
  assign _T_18740 = valid_2_1 ? 6'h1 : _T_18739; // @[Mux.scala 31:69:@907.4]
  assign select_2 = valid_2_0 ? 6'h0 : _T_18740; // @[Mux.scala 31:69:@908.4]
  assign _GEN_129 = 6'h1 == select_2 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@910.4]
  assign _GEN_130 = 6'h2 == select_2 ? io_inData_2 : _GEN_129; // @[Switch.scala 33:19:@910.4]
  assign _GEN_131 = 6'h3 == select_2 ? io_inData_3 : _GEN_130; // @[Switch.scala 33:19:@910.4]
  assign _GEN_132 = 6'h4 == select_2 ? io_inData_4 : _GEN_131; // @[Switch.scala 33:19:@910.4]
  assign _GEN_133 = 6'h5 == select_2 ? io_inData_5 : _GEN_132; // @[Switch.scala 33:19:@910.4]
  assign _GEN_134 = 6'h6 == select_2 ? io_inData_6 : _GEN_133; // @[Switch.scala 33:19:@910.4]
  assign _GEN_135 = 6'h7 == select_2 ? io_inData_7 : _GEN_134; // @[Switch.scala 33:19:@910.4]
  assign _GEN_136 = 6'h8 == select_2 ? io_inData_8 : _GEN_135; // @[Switch.scala 33:19:@910.4]
  assign _GEN_137 = 6'h9 == select_2 ? io_inData_9 : _GEN_136; // @[Switch.scala 33:19:@910.4]
  assign _GEN_138 = 6'ha == select_2 ? io_inData_10 : _GEN_137; // @[Switch.scala 33:19:@910.4]
  assign _GEN_139 = 6'hb == select_2 ? io_inData_11 : _GEN_138; // @[Switch.scala 33:19:@910.4]
  assign _GEN_140 = 6'hc == select_2 ? io_inData_12 : _GEN_139; // @[Switch.scala 33:19:@910.4]
  assign _GEN_141 = 6'hd == select_2 ? io_inData_13 : _GEN_140; // @[Switch.scala 33:19:@910.4]
  assign _GEN_142 = 6'he == select_2 ? io_inData_14 : _GEN_141; // @[Switch.scala 33:19:@910.4]
  assign _GEN_143 = 6'hf == select_2 ? io_inData_15 : _GEN_142; // @[Switch.scala 33:19:@910.4]
  assign _GEN_144 = 6'h10 == select_2 ? io_inData_16 : _GEN_143; // @[Switch.scala 33:19:@910.4]
  assign _GEN_145 = 6'h11 == select_2 ? io_inData_17 : _GEN_144; // @[Switch.scala 33:19:@910.4]
  assign _GEN_146 = 6'h12 == select_2 ? io_inData_18 : _GEN_145; // @[Switch.scala 33:19:@910.4]
  assign _GEN_147 = 6'h13 == select_2 ? io_inData_19 : _GEN_146; // @[Switch.scala 33:19:@910.4]
  assign _GEN_148 = 6'h14 == select_2 ? io_inData_20 : _GEN_147; // @[Switch.scala 33:19:@910.4]
  assign _GEN_149 = 6'h15 == select_2 ? io_inData_21 : _GEN_148; // @[Switch.scala 33:19:@910.4]
  assign _GEN_150 = 6'h16 == select_2 ? io_inData_22 : _GEN_149; // @[Switch.scala 33:19:@910.4]
  assign _GEN_151 = 6'h17 == select_2 ? io_inData_23 : _GEN_150; // @[Switch.scala 33:19:@910.4]
  assign _GEN_152 = 6'h18 == select_2 ? io_inData_24 : _GEN_151; // @[Switch.scala 33:19:@910.4]
  assign _GEN_153 = 6'h19 == select_2 ? io_inData_25 : _GEN_152; // @[Switch.scala 33:19:@910.4]
  assign _GEN_154 = 6'h1a == select_2 ? io_inData_26 : _GEN_153; // @[Switch.scala 33:19:@910.4]
  assign _GEN_155 = 6'h1b == select_2 ? io_inData_27 : _GEN_154; // @[Switch.scala 33:19:@910.4]
  assign _GEN_156 = 6'h1c == select_2 ? io_inData_28 : _GEN_155; // @[Switch.scala 33:19:@910.4]
  assign _GEN_157 = 6'h1d == select_2 ? io_inData_29 : _GEN_156; // @[Switch.scala 33:19:@910.4]
  assign _GEN_158 = 6'h1e == select_2 ? io_inData_30 : _GEN_157; // @[Switch.scala 33:19:@910.4]
  assign _GEN_159 = 6'h1f == select_2 ? io_inData_31 : _GEN_158; // @[Switch.scala 33:19:@910.4]
  assign _GEN_160 = 6'h20 == select_2 ? io_inData_32 : _GEN_159; // @[Switch.scala 33:19:@910.4]
  assign _GEN_161 = 6'h21 == select_2 ? io_inData_33 : _GEN_160; // @[Switch.scala 33:19:@910.4]
  assign _GEN_162 = 6'h22 == select_2 ? io_inData_34 : _GEN_161; // @[Switch.scala 33:19:@910.4]
  assign _GEN_163 = 6'h23 == select_2 ? io_inData_35 : _GEN_162; // @[Switch.scala 33:19:@910.4]
  assign _GEN_164 = 6'h24 == select_2 ? io_inData_36 : _GEN_163; // @[Switch.scala 33:19:@910.4]
  assign _GEN_165 = 6'h25 == select_2 ? io_inData_37 : _GEN_164; // @[Switch.scala 33:19:@910.4]
  assign _GEN_166 = 6'h26 == select_2 ? io_inData_38 : _GEN_165; // @[Switch.scala 33:19:@910.4]
  assign _GEN_167 = 6'h27 == select_2 ? io_inData_39 : _GEN_166; // @[Switch.scala 33:19:@910.4]
  assign _GEN_168 = 6'h28 == select_2 ? io_inData_40 : _GEN_167; // @[Switch.scala 33:19:@910.4]
  assign _GEN_169 = 6'h29 == select_2 ? io_inData_41 : _GEN_168; // @[Switch.scala 33:19:@910.4]
  assign _GEN_170 = 6'h2a == select_2 ? io_inData_42 : _GEN_169; // @[Switch.scala 33:19:@910.4]
  assign _GEN_171 = 6'h2b == select_2 ? io_inData_43 : _GEN_170; // @[Switch.scala 33:19:@910.4]
  assign _GEN_172 = 6'h2c == select_2 ? io_inData_44 : _GEN_171; // @[Switch.scala 33:19:@910.4]
  assign _GEN_173 = 6'h2d == select_2 ? io_inData_45 : _GEN_172; // @[Switch.scala 33:19:@910.4]
  assign _GEN_174 = 6'h2e == select_2 ? io_inData_46 : _GEN_173; // @[Switch.scala 33:19:@910.4]
  assign _GEN_175 = 6'h2f == select_2 ? io_inData_47 : _GEN_174; // @[Switch.scala 33:19:@910.4]
  assign _GEN_176 = 6'h30 == select_2 ? io_inData_48 : _GEN_175; // @[Switch.scala 33:19:@910.4]
  assign _GEN_177 = 6'h31 == select_2 ? io_inData_49 : _GEN_176; // @[Switch.scala 33:19:@910.4]
  assign _GEN_178 = 6'h32 == select_2 ? io_inData_50 : _GEN_177; // @[Switch.scala 33:19:@910.4]
  assign _GEN_179 = 6'h33 == select_2 ? io_inData_51 : _GEN_178; // @[Switch.scala 33:19:@910.4]
  assign _GEN_180 = 6'h34 == select_2 ? io_inData_52 : _GEN_179; // @[Switch.scala 33:19:@910.4]
  assign _GEN_181 = 6'h35 == select_2 ? io_inData_53 : _GEN_180; // @[Switch.scala 33:19:@910.4]
  assign _GEN_182 = 6'h36 == select_2 ? io_inData_54 : _GEN_181; // @[Switch.scala 33:19:@910.4]
  assign _GEN_183 = 6'h37 == select_2 ? io_inData_55 : _GEN_182; // @[Switch.scala 33:19:@910.4]
  assign _GEN_184 = 6'h38 == select_2 ? io_inData_56 : _GEN_183; // @[Switch.scala 33:19:@910.4]
  assign _GEN_185 = 6'h39 == select_2 ? io_inData_57 : _GEN_184; // @[Switch.scala 33:19:@910.4]
  assign _GEN_186 = 6'h3a == select_2 ? io_inData_58 : _GEN_185; // @[Switch.scala 33:19:@910.4]
  assign _GEN_187 = 6'h3b == select_2 ? io_inData_59 : _GEN_186; // @[Switch.scala 33:19:@910.4]
  assign _GEN_188 = 6'h3c == select_2 ? io_inData_60 : _GEN_187; // @[Switch.scala 33:19:@910.4]
  assign _GEN_189 = 6'h3d == select_2 ? io_inData_61 : _GEN_188; // @[Switch.scala 33:19:@910.4]
  assign _GEN_190 = 6'h3e == select_2 ? io_inData_62 : _GEN_189; // @[Switch.scala 33:19:@910.4]
  assign _T_18749 = {valid_2_7,valid_2_6,valid_2_5,valid_2_4,valid_2_3,valid_2_2,valid_2_1,valid_2_0}; // @[Switch.scala 34:32:@917.4]
  assign _T_18757 = {valid_2_15,valid_2_14,valid_2_13,valid_2_12,valid_2_11,valid_2_10,valid_2_9,valid_2_8,_T_18749}; // @[Switch.scala 34:32:@925.4]
  assign _T_18764 = {valid_2_23,valid_2_22,valid_2_21,valid_2_20,valid_2_19,valid_2_18,valid_2_17,valid_2_16}; // @[Switch.scala 34:32:@932.4]
  assign _T_18773 = {valid_2_31,valid_2_30,valid_2_29,valid_2_28,valid_2_27,valid_2_26,valid_2_25,valid_2_24,_T_18764,_T_18757}; // @[Switch.scala 34:32:@941.4]
  assign _T_18780 = {valid_2_39,valid_2_38,valid_2_37,valid_2_36,valid_2_35,valid_2_34,valid_2_33,valid_2_32}; // @[Switch.scala 34:32:@948.4]
  assign _T_18788 = {valid_2_47,valid_2_46,valid_2_45,valid_2_44,valid_2_43,valid_2_42,valid_2_41,valid_2_40,_T_18780}; // @[Switch.scala 34:32:@956.4]
  assign _T_18795 = {valid_2_55,valid_2_54,valid_2_53,valid_2_52,valid_2_51,valid_2_50,valid_2_49,valid_2_48}; // @[Switch.scala 34:32:@963.4]
  assign _T_18804 = {valid_2_63,valid_2_62,valid_2_61,valid_2_60,valid_2_59,valid_2_58,valid_2_57,valid_2_56,_T_18795,_T_18788}; // @[Switch.scala 34:32:@972.4]
  assign _T_18805 = {_T_18804,_T_18773}; // @[Switch.scala 34:32:@973.4]
  assign _T_18809 = io_inAddr_0 == 6'h3; // @[Switch.scala 30:53:@976.4]
  assign valid_3_0 = io_inValid_0 & _T_18809; // @[Switch.scala 30:36:@977.4]
  assign _T_18812 = io_inAddr_1 == 6'h3; // @[Switch.scala 30:53:@979.4]
  assign valid_3_1 = io_inValid_1 & _T_18812; // @[Switch.scala 30:36:@980.4]
  assign _T_18815 = io_inAddr_2 == 6'h3; // @[Switch.scala 30:53:@982.4]
  assign valid_3_2 = io_inValid_2 & _T_18815; // @[Switch.scala 30:36:@983.4]
  assign _T_18818 = io_inAddr_3 == 6'h3; // @[Switch.scala 30:53:@985.4]
  assign valid_3_3 = io_inValid_3 & _T_18818; // @[Switch.scala 30:36:@986.4]
  assign _T_18821 = io_inAddr_4 == 6'h3; // @[Switch.scala 30:53:@988.4]
  assign valid_3_4 = io_inValid_4 & _T_18821; // @[Switch.scala 30:36:@989.4]
  assign _T_18824 = io_inAddr_5 == 6'h3; // @[Switch.scala 30:53:@991.4]
  assign valid_3_5 = io_inValid_5 & _T_18824; // @[Switch.scala 30:36:@992.4]
  assign _T_18827 = io_inAddr_6 == 6'h3; // @[Switch.scala 30:53:@994.4]
  assign valid_3_6 = io_inValid_6 & _T_18827; // @[Switch.scala 30:36:@995.4]
  assign _T_18830 = io_inAddr_7 == 6'h3; // @[Switch.scala 30:53:@997.4]
  assign valid_3_7 = io_inValid_7 & _T_18830; // @[Switch.scala 30:36:@998.4]
  assign _T_18833 = io_inAddr_8 == 6'h3; // @[Switch.scala 30:53:@1000.4]
  assign valid_3_8 = io_inValid_8 & _T_18833; // @[Switch.scala 30:36:@1001.4]
  assign _T_18836 = io_inAddr_9 == 6'h3; // @[Switch.scala 30:53:@1003.4]
  assign valid_3_9 = io_inValid_9 & _T_18836; // @[Switch.scala 30:36:@1004.4]
  assign _T_18839 = io_inAddr_10 == 6'h3; // @[Switch.scala 30:53:@1006.4]
  assign valid_3_10 = io_inValid_10 & _T_18839; // @[Switch.scala 30:36:@1007.4]
  assign _T_18842 = io_inAddr_11 == 6'h3; // @[Switch.scala 30:53:@1009.4]
  assign valid_3_11 = io_inValid_11 & _T_18842; // @[Switch.scala 30:36:@1010.4]
  assign _T_18845 = io_inAddr_12 == 6'h3; // @[Switch.scala 30:53:@1012.4]
  assign valid_3_12 = io_inValid_12 & _T_18845; // @[Switch.scala 30:36:@1013.4]
  assign _T_18848 = io_inAddr_13 == 6'h3; // @[Switch.scala 30:53:@1015.4]
  assign valid_3_13 = io_inValid_13 & _T_18848; // @[Switch.scala 30:36:@1016.4]
  assign _T_18851 = io_inAddr_14 == 6'h3; // @[Switch.scala 30:53:@1018.4]
  assign valid_3_14 = io_inValid_14 & _T_18851; // @[Switch.scala 30:36:@1019.4]
  assign _T_18854 = io_inAddr_15 == 6'h3; // @[Switch.scala 30:53:@1021.4]
  assign valid_3_15 = io_inValid_15 & _T_18854; // @[Switch.scala 30:36:@1022.4]
  assign _T_18857 = io_inAddr_16 == 6'h3; // @[Switch.scala 30:53:@1024.4]
  assign valid_3_16 = io_inValid_16 & _T_18857; // @[Switch.scala 30:36:@1025.4]
  assign _T_18860 = io_inAddr_17 == 6'h3; // @[Switch.scala 30:53:@1027.4]
  assign valid_3_17 = io_inValid_17 & _T_18860; // @[Switch.scala 30:36:@1028.4]
  assign _T_18863 = io_inAddr_18 == 6'h3; // @[Switch.scala 30:53:@1030.4]
  assign valid_3_18 = io_inValid_18 & _T_18863; // @[Switch.scala 30:36:@1031.4]
  assign _T_18866 = io_inAddr_19 == 6'h3; // @[Switch.scala 30:53:@1033.4]
  assign valid_3_19 = io_inValid_19 & _T_18866; // @[Switch.scala 30:36:@1034.4]
  assign _T_18869 = io_inAddr_20 == 6'h3; // @[Switch.scala 30:53:@1036.4]
  assign valid_3_20 = io_inValid_20 & _T_18869; // @[Switch.scala 30:36:@1037.4]
  assign _T_18872 = io_inAddr_21 == 6'h3; // @[Switch.scala 30:53:@1039.4]
  assign valid_3_21 = io_inValid_21 & _T_18872; // @[Switch.scala 30:36:@1040.4]
  assign _T_18875 = io_inAddr_22 == 6'h3; // @[Switch.scala 30:53:@1042.4]
  assign valid_3_22 = io_inValid_22 & _T_18875; // @[Switch.scala 30:36:@1043.4]
  assign _T_18878 = io_inAddr_23 == 6'h3; // @[Switch.scala 30:53:@1045.4]
  assign valid_3_23 = io_inValid_23 & _T_18878; // @[Switch.scala 30:36:@1046.4]
  assign _T_18881 = io_inAddr_24 == 6'h3; // @[Switch.scala 30:53:@1048.4]
  assign valid_3_24 = io_inValid_24 & _T_18881; // @[Switch.scala 30:36:@1049.4]
  assign _T_18884 = io_inAddr_25 == 6'h3; // @[Switch.scala 30:53:@1051.4]
  assign valid_3_25 = io_inValid_25 & _T_18884; // @[Switch.scala 30:36:@1052.4]
  assign _T_18887 = io_inAddr_26 == 6'h3; // @[Switch.scala 30:53:@1054.4]
  assign valid_3_26 = io_inValid_26 & _T_18887; // @[Switch.scala 30:36:@1055.4]
  assign _T_18890 = io_inAddr_27 == 6'h3; // @[Switch.scala 30:53:@1057.4]
  assign valid_3_27 = io_inValid_27 & _T_18890; // @[Switch.scala 30:36:@1058.4]
  assign _T_18893 = io_inAddr_28 == 6'h3; // @[Switch.scala 30:53:@1060.4]
  assign valid_3_28 = io_inValid_28 & _T_18893; // @[Switch.scala 30:36:@1061.4]
  assign _T_18896 = io_inAddr_29 == 6'h3; // @[Switch.scala 30:53:@1063.4]
  assign valid_3_29 = io_inValid_29 & _T_18896; // @[Switch.scala 30:36:@1064.4]
  assign _T_18899 = io_inAddr_30 == 6'h3; // @[Switch.scala 30:53:@1066.4]
  assign valid_3_30 = io_inValid_30 & _T_18899; // @[Switch.scala 30:36:@1067.4]
  assign _T_18902 = io_inAddr_31 == 6'h3; // @[Switch.scala 30:53:@1069.4]
  assign valid_3_31 = io_inValid_31 & _T_18902; // @[Switch.scala 30:36:@1070.4]
  assign _T_18905 = io_inAddr_32 == 6'h3; // @[Switch.scala 30:53:@1072.4]
  assign valid_3_32 = io_inValid_32 & _T_18905; // @[Switch.scala 30:36:@1073.4]
  assign _T_18908 = io_inAddr_33 == 6'h3; // @[Switch.scala 30:53:@1075.4]
  assign valid_3_33 = io_inValid_33 & _T_18908; // @[Switch.scala 30:36:@1076.4]
  assign _T_18911 = io_inAddr_34 == 6'h3; // @[Switch.scala 30:53:@1078.4]
  assign valid_3_34 = io_inValid_34 & _T_18911; // @[Switch.scala 30:36:@1079.4]
  assign _T_18914 = io_inAddr_35 == 6'h3; // @[Switch.scala 30:53:@1081.4]
  assign valid_3_35 = io_inValid_35 & _T_18914; // @[Switch.scala 30:36:@1082.4]
  assign _T_18917 = io_inAddr_36 == 6'h3; // @[Switch.scala 30:53:@1084.4]
  assign valid_3_36 = io_inValid_36 & _T_18917; // @[Switch.scala 30:36:@1085.4]
  assign _T_18920 = io_inAddr_37 == 6'h3; // @[Switch.scala 30:53:@1087.4]
  assign valid_3_37 = io_inValid_37 & _T_18920; // @[Switch.scala 30:36:@1088.4]
  assign _T_18923 = io_inAddr_38 == 6'h3; // @[Switch.scala 30:53:@1090.4]
  assign valid_3_38 = io_inValid_38 & _T_18923; // @[Switch.scala 30:36:@1091.4]
  assign _T_18926 = io_inAddr_39 == 6'h3; // @[Switch.scala 30:53:@1093.4]
  assign valid_3_39 = io_inValid_39 & _T_18926; // @[Switch.scala 30:36:@1094.4]
  assign _T_18929 = io_inAddr_40 == 6'h3; // @[Switch.scala 30:53:@1096.4]
  assign valid_3_40 = io_inValid_40 & _T_18929; // @[Switch.scala 30:36:@1097.4]
  assign _T_18932 = io_inAddr_41 == 6'h3; // @[Switch.scala 30:53:@1099.4]
  assign valid_3_41 = io_inValid_41 & _T_18932; // @[Switch.scala 30:36:@1100.4]
  assign _T_18935 = io_inAddr_42 == 6'h3; // @[Switch.scala 30:53:@1102.4]
  assign valid_3_42 = io_inValid_42 & _T_18935; // @[Switch.scala 30:36:@1103.4]
  assign _T_18938 = io_inAddr_43 == 6'h3; // @[Switch.scala 30:53:@1105.4]
  assign valid_3_43 = io_inValid_43 & _T_18938; // @[Switch.scala 30:36:@1106.4]
  assign _T_18941 = io_inAddr_44 == 6'h3; // @[Switch.scala 30:53:@1108.4]
  assign valid_3_44 = io_inValid_44 & _T_18941; // @[Switch.scala 30:36:@1109.4]
  assign _T_18944 = io_inAddr_45 == 6'h3; // @[Switch.scala 30:53:@1111.4]
  assign valid_3_45 = io_inValid_45 & _T_18944; // @[Switch.scala 30:36:@1112.4]
  assign _T_18947 = io_inAddr_46 == 6'h3; // @[Switch.scala 30:53:@1114.4]
  assign valid_3_46 = io_inValid_46 & _T_18947; // @[Switch.scala 30:36:@1115.4]
  assign _T_18950 = io_inAddr_47 == 6'h3; // @[Switch.scala 30:53:@1117.4]
  assign valid_3_47 = io_inValid_47 & _T_18950; // @[Switch.scala 30:36:@1118.4]
  assign _T_18953 = io_inAddr_48 == 6'h3; // @[Switch.scala 30:53:@1120.4]
  assign valid_3_48 = io_inValid_48 & _T_18953; // @[Switch.scala 30:36:@1121.4]
  assign _T_18956 = io_inAddr_49 == 6'h3; // @[Switch.scala 30:53:@1123.4]
  assign valid_3_49 = io_inValid_49 & _T_18956; // @[Switch.scala 30:36:@1124.4]
  assign _T_18959 = io_inAddr_50 == 6'h3; // @[Switch.scala 30:53:@1126.4]
  assign valid_3_50 = io_inValid_50 & _T_18959; // @[Switch.scala 30:36:@1127.4]
  assign _T_18962 = io_inAddr_51 == 6'h3; // @[Switch.scala 30:53:@1129.4]
  assign valid_3_51 = io_inValid_51 & _T_18962; // @[Switch.scala 30:36:@1130.4]
  assign _T_18965 = io_inAddr_52 == 6'h3; // @[Switch.scala 30:53:@1132.4]
  assign valid_3_52 = io_inValid_52 & _T_18965; // @[Switch.scala 30:36:@1133.4]
  assign _T_18968 = io_inAddr_53 == 6'h3; // @[Switch.scala 30:53:@1135.4]
  assign valid_3_53 = io_inValid_53 & _T_18968; // @[Switch.scala 30:36:@1136.4]
  assign _T_18971 = io_inAddr_54 == 6'h3; // @[Switch.scala 30:53:@1138.4]
  assign valid_3_54 = io_inValid_54 & _T_18971; // @[Switch.scala 30:36:@1139.4]
  assign _T_18974 = io_inAddr_55 == 6'h3; // @[Switch.scala 30:53:@1141.4]
  assign valid_3_55 = io_inValid_55 & _T_18974; // @[Switch.scala 30:36:@1142.4]
  assign _T_18977 = io_inAddr_56 == 6'h3; // @[Switch.scala 30:53:@1144.4]
  assign valid_3_56 = io_inValid_56 & _T_18977; // @[Switch.scala 30:36:@1145.4]
  assign _T_18980 = io_inAddr_57 == 6'h3; // @[Switch.scala 30:53:@1147.4]
  assign valid_3_57 = io_inValid_57 & _T_18980; // @[Switch.scala 30:36:@1148.4]
  assign _T_18983 = io_inAddr_58 == 6'h3; // @[Switch.scala 30:53:@1150.4]
  assign valid_3_58 = io_inValid_58 & _T_18983; // @[Switch.scala 30:36:@1151.4]
  assign _T_18986 = io_inAddr_59 == 6'h3; // @[Switch.scala 30:53:@1153.4]
  assign valid_3_59 = io_inValid_59 & _T_18986; // @[Switch.scala 30:36:@1154.4]
  assign _T_18989 = io_inAddr_60 == 6'h3; // @[Switch.scala 30:53:@1156.4]
  assign valid_3_60 = io_inValid_60 & _T_18989; // @[Switch.scala 30:36:@1157.4]
  assign _T_18992 = io_inAddr_61 == 6'h3; // @[Switch.scala 30:53:@1159.4]
  assign valid_3_61 = io_inValid_61 & _T_18992; // @[Switch.scala 30:36:@1160.4]
  assign _T_18995 = io_inAddr_62 == 6'h3; // @[Switch.scala 30:53:@1162.4]
  assign valid_3_62 = io_inValid_62 & _T_18995; // @[Switch.scala 30:36:@1163.4]
  assign _T_18998 = io_inAddr_63 == 6'h3; // @[Switch.scala 30:53:@1165.4]
  assign valid_3_63 = io_inValid_63 & _T_18998; // @[Switch.scala 30:36:@1166.4]
  assign _T_19064 = valid_3_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@1168.4]
  assign _T_19065 = valid_3_61 ? 6'h3d : _T_19064; // @[Mux.scala 31:69:@1169.4]
  assign _T_19066 = valid_3_60 ? 6'h3c : _T_19065; // @[Mux.scala 31:69:@1170.4]
  assign _T_19067 = valid_3_59 ? 6'h3b : _T_19066; // @[Mux.scala 31:69:@1171.4]
  assign _T_19068 = valid_3_58 ? 6'h3a : _T_19067; // @[Mux.scala 31:69:@1172.4]
  assign _T_19069 = valid_3_57 ? 6'h39 : _T_19068; // @[Mux.scala 31:69:@1173.4]
  assign _T_19070 = valid_3_56 ? 6'h38 : _T_19069; // @[Mux.scala 31:69:@1174.4]
  assign _T_19071 = valid_3_55 ? 6'h37 : _T_19070; // @[Mux.scala 31:69:@1175.4]
  assign _T_19072 = valid_3_54 ? 6'h36 : _T_19071; // @[Mux.scala 31:69:@1176.4]
  assign _T_19073 = valid_3_53 ? 6'h35 : _T_19072; // @[Mux.scala 31:69:@1177.4]
  assign _T_19074 = valid_3_52 ? 6'h34 : _T_19073; // @[Mux.scala 31:69:@1178.4]
  assign _T_19075 = valid_3_51 ? 6'h33 : _T_19074; // @[Mux.scala 31:69:@1179.4]
  assign _T_19076 = valid_3_50 ? 6'h32 : _T_19075; // @[Mux.scala 31:69:@1180.4]
  assign _T_19077 = valid_3_49 ? 6'h31 : _T_19076; // @[Mux.scala 31:69:@1181.4]
  assign _T_19078 = valid_3_48 ? 6'h30 : _T_19077; // @[Mux.scala 31:69:@1182.4]
  assign _T_19079 = valid_3_47 ? 6'h2f : _T_19078; // @[Mux.scala 31:69:@1183.4]
  assign _T_19080 = valid_3_46 ? 6'h2e : _T_19079; // @[Mux.scala 31:69:@1184.4]
  assign _T_19081 = valid_3_45 ? 6'h2d : _T_19080; // @[Mux.scala 31:69:@1185.4]
  assign _T_19082 = valid_3_44 ? 6'h2c : _T_19081; // @[Mux.scala 31:69:@1186.4]
  assign _T_19083 = valid_3_43 ? 6'h2b : _T_19082; // @[Mux.scala 31:69:@1187.4]
  assign _T_19084 = valid_3_42 ? 6'h2a : _T_19083; // @[Mux.scala 31:69:@1188.4]
  assign _T_19085 = valid_3_41 ? 6'h29 : _T_19084; // @[Mux.scala 31:69:@1189.4]
  assign _T_19086 = valid_3_40 ? 6'h28 : _T_19085; // @[Mux.scala 31:69:@1190.4]
  assign _T_19087 = valid_3_39 ? 6'h27 : _T_19086; // @[Mux.scala 31:69:@1191.4]
  assign _T_19088 = valid_3_38 ? 6'h26 : _T_19087; // @[Mux.scala 31:69:@1192.4]
  assign _T_19089 = valid_3_37 ? 6'h25 : _T_19088; // @[Mux.scala 31:69:@1193.4]
  assign _T_19090 = valid_3_36 ? 6'h24 : _T_19089; // @[Mux.scala 31:69:@1194.4]
  assign _T_19091 = valid_3_35 ? 6'h23 : _T_19090; // @[Mux.scala 31:69:@1195.4]
  assign _T_19092 = valid_3_34 ? 6'h22 : _T_19091; // @[Mux.scala 31:69:@1196.4]
  assign _T_19093 = valid_3_33 ? 6'h21 : _T_19092; // @[Mux.scala 31:69:@1197.4]
  assign _T_19094 = valid_3_32 ? 6'h20 : _T_19093; // @[Mux.scala 31:69:@1198.4]
  assign _T_19095 = valid_3_31 ? 6'h1f : _T_19094; // @[Mux.scala 31:69:@1199.4]
  assign _T_19096 = valid_3_30 ? 6'h1e : _T_19095; // @[Mux.scala 31:69:@1200.4]
  assign _T_19097 = valid_3_29 ? 6'h1d : _T_19096; // @[Mux.scala 31:69:@1201.4]
  assign _T_19098 = valid_3_28 ? 6'h1c : _T_19097; // @[Mux.scala 31:69:@1202.4]
  assign _T_19099 = valid_3_27 ? 6'h1b : _T_19098; // @[Mux.scala 31:69:@1203.4]
  assign _T_19100 = valid_3_26 ? 6'h1a : _T_19099; // @[Mux.scala 31:69:@1204.4]
  assign _T_19101 = valid_3_25 ? 6'h19 : _T_19100; // @[Mux.scala 31:69:@1205.4]
  assign _T_19102 = valid_3_24 ? 6'h18 : _T_19101; // @[Mux.scala 31:69:@1206.4]
  assign _T_19103 = valid_3_23 ? 6'h17 : _T_19102; // @[Mux.scala 31:69:@1207.4]
  assign _T_19104 = valid_3_22 ? 6'h16 : _T_19103; // @[Mux.scala 31:69:@1208.4]
  assign _T_19105 = valid_3_21 ? 6'h15 : _T_19104; // @[Mux.scala 31:69:@1209.4]
  assign _T_19106 = valid_3_20 ? 6'h14 : _T_19105; // @[Mux.scala 31:69:@1210.4]
  assign _T_19107 = valid_3_19 ? 6'h13 : _T_19106; // @[Mux.scala 31:69:@1211.4]
  assign _T_19108 = valid_3_18 ? 6'h12 : _T_19107; // @[Mux.scala 31:69:@1212.4]
  assign _T_19109 = valid_3_17 ? 6'h11 : _T_19108; // @[Mux.scala 31:69:@1213.4]
  assign _T_19110 = valid_3_16 ? 6'h10 : _T_19109; // @[Mux.scala 31:69:@1214.4]
  assign _T_19111 = valid_3_15 ? 6'hf : _T_19110; // @[Mux.scala 31:69:@1215.4]
  assign _T_19112 = valid_3_14 ? 6'he : _T_19111; // @[Mux.scala 31:69:@1216.4]
  assign _T_19113 = valid_3_13 ? 6'hd : _T_19112; // @[Mux.scala 31:69:@1217.4]
  assign _T_19114 = valid_3_12 ? 6'hc : _T_19113; // @[Mux.scala 31:69:@1218.4]
  assign _T_19115 = valid_3_11 ? 6'hb : _T_19114; // @[Mux.scala 31:69:@1219.4]
  assign _T_19116 = valid_3_10 ? 6'ha : _T_19115; // @[Mux.scala 31:69:@1220.4]
  assign _T_19117 = valid_3_9 ? 6'h9 : _T_19116; // @[Mux.scala 31:69:@1221.4]
  assign _T_19118 = valid_3_8 ? 6'h8 : _T_19117; // @[Mux.scala 31:69:@1222.4]
  assign _T_19119 = valid_3_7 ? 6'h7 : _T_19118; // @[Mux.scala 31:69:@1223.4]
  assign _T_19120 = valid_3_6 ? 6'h6 : _T_19119; // @[Mux.scala 31:69:@1224.4]
  assign _T_19121 = valid_3_5 ? 6'h5 : _T_19120; // @[Mux.scala 31:69:@1225.4]
  assign _T_19122 = valid_3_4 ? 6'h4 : _T_19121; // @[Mux.scala 31:69:@1226.4]
  assign _T_19123 = valid_3_3 ? 6'h3 : _T_19122; // @[Mux.scala 31:69:@1227.4]
  assign _T_19124 = valid_3_2 ? 6'h2 : _T_19123; // @[Mux.scala 31:69:@1228.4]
  assign _T_19125 = valid_3_1 ? 6'h1 : _T_19124; // @[Mux.scala 31:69:@1229.4]
  assign select_3 = valid_3_0 ? 6'h0 : _T_19125; // @[Mux.scala 31:69:@1230.4]
  assign _GEN_193 = 6'h1 == select_3 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_194 = 6'h2 == select_3 ? io_inData_2 : _GEN_193; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_195 = 6'h3 == select_3 ? io_inData_3 : _GEN_194; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_196 = 6'h4 == select_3 ? io_inData_4 : _GEN_195; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_197 = 6'h5 == select_3 ? io_inData_5 : _GEN_196; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_198 = 6'h6 == select_3 ? io_inData_6 : _GEN_197; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_199 = 6'h7 == select_3 ? io_inData_7 : _GEN_198; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_200 = 6'h8 == select_3 ? io_inData_8 : _GEN_199; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_201 = 6'h9 == select_3 ? io_inData_9 : _GEN_200; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_202 = 6'ha == select_3 ? io_inData_10 : _GEN_201; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_203 = 6'hb == select_3 ? io_inData_11 : _GEN_202; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_204 = 6'hc == select_3 ? io_inData_12 : _GEN_203; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_205 = 6'hd == select_3 ? io_inData_13 : _GEN_204; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_206 = 6'he == select_3 ? io_inData_14 : _GEN_205; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_207 = 6'hf == select_3 ? io_inData_15 : _GEN_206; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_208 = 6'h10 == select_3 ? io_inData_16 : _GEN_207; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_209 = 6'h11 == select_3 ? io_inData_17 : _GEN_208; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_210 = 6'h12 == select_3 ? io_inData_18 : _GEN_209; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_211 = 6'h13 == select_3 ? io_inData_19 : _GEN_210; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_212 = 6'h14 == select_3 ? io_inData_20 : _GEN_211; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_213 = 6'h15 == select_3 ? io_inData_21 : _GEN_212; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_214 = 6'h16 == select_3 ? io_inData_22 : _GEN_213; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_215 = 6'h17 == select_3 ? io_inData_23 : _GEN_214; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_216 = 6'h18 == select_3 ? io_inData_24 : _GEN_215; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_217 = 6'h19 == select_3 ? io_inData_25 : _GEN_216; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_218 = 6'h1a == select_3 ? io_inData_26 : _GEN_217; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_219 = 6'h1b == select_3 ? io_inData_27 : _GEN_218; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_220 = 6'h1c == select_3 ? io_inData_28 : _GEN_219; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_221 = 6'h1d == select_3 ? io_inData_29 : _GEN_220; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_222 = 6'h1e == select_3 ? io_inData_30 : _GEN_221; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_223 = 6'h1f == select_3 ? io_inData_31 : _GEN_222; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_224 = 6'h20 == select_3 ? io_inData_32 : _GEN_223; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_225 = 6'h21 == select_3 ? io_inData_33 : _GEN_224; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_226 = 6'h22 == select_3 ? io_inData_34 : _GEN_225; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_227 = 6'h23 == select_3 ? io_inData_35 : _GEN_226; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_228 = 6'h24 == select_3 ? io_inData_36 : _GEN_227; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_229 = 6'h25 == select_3 ? io_inData_37 : _GEN_228; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_230 = 6'h26 == select_3 ? io_inData_38 : _GEN_229; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_231 = 6'h27 == select_3 ? io_inData_39 : _GEN_230; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_232 = 6'h28 == select_3 ? io_inData_40 : _GEN_231; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_233 = 6'h29 == select_3 ? io_inData_41 : _GEN_232; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_234 = 6'h2a == select_3 ? io_inData_42 : _GEN_233; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_235 = 6'h2b == select_3 ? io_inData_43 : _GEN_234; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_236 = 6'h2c == select_3 ? io_inData_44 : _GEN_235; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_237 = 6'h2d == select_3 ? io_inData_45 : _GEN_236; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_238 = 6'h2e == select_3 ? io_inData_46 : _GEN_237; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_239 = 6'h2f == select_3 ? io_inData_47 : _GEN_238; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_240 = 6'h30 == select_3 ? io_inData_48 : _GEN_239; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_241 = 6'h31 == select_3 ? io_inData_49 : _GEN_240; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_242 = 6'h32 == select_3 ? io_inData_50 : _GEN_241; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_243 = 6'h33 == select_3 ? io_inData_51 : _GEN_242; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_244 = 6'h34 == select_3 ? io_inData_52 : _GEN_243; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_245 = 6'h35 == select_3 ? io_inData_53 : _GEN_244; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_246 = 6'h36 == select_3 ? io_inData_54 : _GEN_245; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_247 = 6'h37 == select_3 ? io_inData_55 : _GEN_246; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_248 = 6'h38 == select_3 ? io_inData_56 : _GEN_247; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_249 = 6'h39 == select_3 ? io_inData_57 : _GEN_248; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_250 = 6'h3a == select_3 ? io_inData_58 : _GEN_249; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_251 = 6'h3b == select_3 ? io_inData_59 : _GEN_250; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_252 = 6'h3c == select_3 ? io_inData_60 : _GEN_251; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_253 = 6'h3d == select_3 ? io_inData_61 : _GEN_252; // @[Switch.scala 33:19:@1232.4]
  assign _GEN_254 = 6'h3e == select_3 ? io_inData_62 : _GEN_253; // @[Switch.scala 33:19:@1232.4]
  assign _T_19134 = {valid_3_7,valid_3_6,valid_3_5,valid_3_4,valid_3_3,valid_3_2,valid_3_1,valid_3_0}; // @[Switch.scala 34:32:@1239.4]
  assign _T_19142 = {valid_3_15,valid_3_14,valid_3_13,valid_3_12,valid_3_11,valid_3_10,valid_3_9,valid_3_8,_T_19134}; // @[Switch.scala 34:32:@1247.4]
  assign _T_19149 = {valid_3_23,valid_3_22,valid_3_21,valid_3_20,valid_3_19,valid_3_18,valid_3_17,valid_3_16}; // @[Switch.scala 34:32:@1254.4]
  assign _T_19158 = {valid_3_31,valid_3_30,valid_3_29,valid_3_28,valid_3_27,valid_3_26,valid_3_25,valid_3_24,_T_19149,_T_19142}; // @[Switch.scala 34:32:@1263.4]
  assign _T_19165 = {valid_3_39,valid_3_38,valid_3_37,valid_3_36,valid_3_35,valid_3_34,valid_3_33,valid_3_32}; // @[Switch.scala 34:32:@1270.4]
  assign _T_19173 = {valid_3_47,valid_3_46,valid_3_45,valid_3_44,valid_3_43,valid_3_42,valid_3_41,valid_3_40,_T_19165}; // @[Switch.scala 34:32:@1278.4]
  assign _T_19180 = {valid_3_55,valid_3_54,valid_3_53,valid_3_52,valid_3_51,valid_3_50,valid_3_49,valid_3_48}; // @[Switch.scala 34:32:@1285.4]
  assign _T_19189 = {valid_3_63,valid_3_62,valid_3_61,valid_3_60,valid_3_59,valid_3_58,valid_3_57,valid_3_56,_T_19180,_T_19173}; // @[Switch.scala 34:32:@1294.4]
  assign _T_19190 = {_T_19189,_T_19158}; // @[Switch.scala 34:32:@1295.4]
  assign _T_19194 = io_inAddr_0 == 6'h4; // @[Switch.scala 30:53:@1298.4]
  assign valid_4_0 = io_inValid_0 & _T_19194; // @[Switch.scala 30:36:@1299.4]
  assign _T_19197 = io_inAddr_1 == 6'h4; // @[Switch.scala 30:53:@1301.4]
  assign valid_4_1 = io_inValid_1 & _T_19197; // @[Switch.scala 30:36:@1302.4]
  assign _T_19200 = io_inAddr_2 == 6'h4; // @[Switch.scala 30:53:@1304.4]
  assign valid_4_2 = io_inValid_2 & _T_19200; // @[Switch.scala 30:36:@1305.4]
  assign _T_19203 = io_inAddr_3 == 6'h4; // @[Switch.scala 30:53:@1307.4]
  assign valid_4_3 = io_inValid_3 & _T_19203; // @[Switch.scala 30:36:@1308.4]
  assign _T_19206 = io_inAddr_4 == 6'h4; // @[Switch.scala 30:53:@1310.4]
  assign valid_4_4 = io_inValid_4 & _T_19206; // @[Switch.scala 30:36:@1311.4]
  assign _T_19209 = io_inAddr_5 == 6'h4; // @[Switch.scala 30:53:@1313.4]
  assign valid_4_5 = io_inValid_5 & _T_19209; // @[Switch.scala 30:36:@1314.4]
  assign _T_19212 = io_inAddr_6 == 6'h4; // @[Switch.scala 30:53:@1316.4]
  assign valid_4_6 = io_inValid_6 & _T_19212; // @[Switch.scala 30:36:@1317.4]
  assign _T_19215 = io_inAddr_7 == 6'h4; // @[Switch.scala 30:53:@1319.4]
  assign valid_4_7 = io_inValid_7 & _T_19215; // @[Switch.scala 30:36:@1320.4]
  assign _T_19218 = io_inAddr_8 == 6'h4; // @[Switch.scala 30:53:@1322.4]
  assign valid_4_8 = io_inValid_8 & _T_19218; // @[Switch.scala 30:36:@1323.4]
  assign _T_19221 = io_inAddr_9 == 6'h4; // @[Switch.scala 30:53:@1325.4]
  assign valid_4_9 = io_inValid_9 & _T_19221; // @[Switch.scala 30:36:@1326.4]
  assign _T_19224 = io_inAddr_10 == 6'h4; // @[Switch.scala 30:53:@1328.4]
  assign valid_4_10 = io_inValid_10 & _T_19224; // @[Switch.scala 30:36:@1329.4]
  assign _T_19227 = io_inAddr_11 == 6'h4; // @[Switch.scala 30:53:@1331.4]
  assign valid_4_11 = io_inValid_11 & _T_19227; // @[Switch.scala 30:36:@1332.4]
  assign _T_19230 = io_inAddr_12 == 6'h4; // @[Switch.scala 30:53:@1334.4]
  assign valid_4_12 = io_inValid_12 & _T_19230; // @[Switch.scala 30:36:@1335.4]
  assign _T_19233 = io_inAddr_13 == 6'h4; // @[Switch.scala 30:53:@1337.4]
  assign valid_4_13 = io_inValid_13 & _T_19233; // @[Switch.scala 30:36:@1338.4]
  assign _T_19236 = io_inAddr_14 == 6'h4; // @[Switch.scala 30:53:@1340.4]
  assign valid_4_14 = io_inValid_14 & _T_19236; // @[Switch.scala 30:36:@1341.4]
  assign _T_19239 = io_inAddr_15 == 6'h4; // @[Switch.scala 30:53:@1343.4]
  assign valid_4_15 = io_inValid_15 & _T_19239; // @[Switch.scala 30:36:@1344.4]
  assign _T_19242 = io_inAddr_16 == 6'h4; // @[Switch.scala 30:53:@1346.4]
  assign valid_4_16 = io_inValid_16 & _T_19242; // @[Switch.scala 30:36:@1347.4]
  assign _T_19245 = io_inAddr_17 == 6'h4; // @[Switch.scala 30:53:@1349.4]
  assign valid_4_17 = io_inValid_17 & _T_19245; // @[Switch.scala 30:36:@1350.4]
  assign _T_19248 = io_inAddr_18 == 6'h4; // @[Switch.scala 30:53:@1352.4]
  assign valid_4_18 = io_inValid_18 & _T_19248; // @[Switch.scala 30:36:@1353.4]
  assign _T_19251 = io_inAddr_19 == 6'h4; // @[Switch.scala 30:53:@1355.4]
  assign valid_4_19 = io_inValid_19 & _T_19251; // @[Switch.scala 30:36:@1356.4]
  assign _T_19254 = io_inAddr_20 == 6'h4; // @[Switch.scala 30:53:@1358.4]
  assign valid_4_20 = io_inValid_20 & _T_19254; // @[Switch.scala 30:36:@1359.4]
  assign _T_19257 = io_inAddr_21 == 6'h4; // @[Switch.scala 30:53:@1361.4]
  assign valid_4_21 = io_inValid_21 & _T_19257; // @[Switch.scala 30:36:@1362.4]
  assign _T_19260 = io_inAddr_22 == 6'h4; // @[Switch.scala 30:53:@1364.4]
  assign valid_4_22 = io_inValid_22 & _T_19260; // @[Switch.scala 30:36:@1365.4]
  assign _T_19263 = io_inAddr_23 == 6'h4; // @[Switch.scala 30:53:@1367.4]
  assign valid_4_23 = io_inValid_23 & _T_19263; // @[Switch.scala 30:36:@1368.4]
  assign _T_19266 = io_inAddr_24 == 6'h4; // @[Switch.scala 30:53:@1370.4]
  assign valid_4_24 = io_inValid_24 & _T_19266; // @[Switch.scala 30:36:@1371.4]
  assign _T_19269 = io_inAddr_25 == 6'h4; // @[Switch.scala 30:53:@1373.4]
  assign valid_4_25 = io_inValid_25 & _T_19269; // @[Switch.scala 30:36:@1374.4]
  assign _T_19272 = io_inAddr_26 == 6'h4; // @[Switch.scala 30:53:@1376.4]
  assign valid_4_26 = io_inValid_26 & _T_19272; // @[Switch.scala 30:36:@1377.4]
  assign _T_19275 = io_inAddr_27 == 6'h4; // @[Switch.scala 30:53:@1379.4]
  assign valid_4_27 = io_inValid_27 & _T_19275; // @[Switch.scala 30:36:@1380.4]
  assign _T_19278 = io_inAddr_28 == 6'h4; // @[Switch.scala 30:53:@1382.4]
  assign valid_4_28 = io_inValid_28 & _T_19278; // @[Switch.scala 30:36:@1383.4]
  assign _T_19281 = io_inAddr_29 == 6'h4; // @[Switch.scala 30:53:@1385.4]
  assign valid_4_29 = io_inValid_29 & _T_19281; // @[Switch.scala 30:36:@1386.4]
  assign _T_19284 = io_inAddr_30 == 6'h4; // @[Switch.scala 30:53:@1388.4]
  assign valid_4_30 = io_inValid_30 & _T_19284; // @[Switch.scala 30:36:@1389.4]
  assign _T_19287 = io_inAddr_31 == 6'h4; // @[Switch.scala 30:53:@1391.4]
  assign valid_4_31 = io_inValid_31 & _T_19287; // @[Switch.scala 30:36:@1392.4]
  assign _T_19290 = io_inAddr_32 == 6'h4; // @[Switch.scala 30:53:@1394.4]
  assign valid_4_32 = io_inValid_32 & _T_19290; // @[Switch.scala 30:36:@1395.4]
  assign _T_19293 = io_inAddr_33 == 6'h4; // @[Switch.scala 30:53:@1397.4]
  assign valid_4_33 = io_inValid_33 & _T_19293; // @[Switch.scala 30:36:@1398.4]
  assign _T_19296 = io_inAddr_34 == 6'h4; // @[Switch.scala 30:53:@1400.4]
  assign valid_4_34 = io_inValid_34 & _T_19296; // @[Switch.scala 30:36:@1401.4]
  assign _T_19299 = io_inAddr_35 == 6'h4; // @[Switch.scala 30:53:@1403.4]
  assign valid_4_35 = io_inValid_35 & _T_19299; // @[Switch.scala 30:36:@1404.4]
  assign _T_19302 = io_inAddr_36 == 6'h4; // @[Switch.scala 30:53:@1406.4]
  assign valid_4_36 = io_inValid_36 & _T_19302; // @[Switch.scala 30:36:@1407.4]
  assign _T_19305 = io_inAddr_37 == 6'h4; // @[Switch.scala 30:53:@1409.4]
  assign valid_4_37 = io_inValid_37 & _T_19305; // @[Switch.scala 30:36:@1410.4]
  assign _T_19308 = io_inAddr_38 == 6'h4; // @[Switch.scala 30:53:@1412.4]
  assign valid_4_38 = io_inValid_38 & _T_19308; // @[Switch.scala 30:36:@1413.4]
  assign _T_19311 = io_inAddr_39 == 6'h4; // @[Switch.scala 30:53:@1415.4]
  assign valid_4_39 = io_inValid_39 & _T_19311; // @[Switch.scala 30:36:@1416.4]
  assign _T_19314 = io_inAddr_40 == 6'h4; // @[Switch.scala 30:53:@1418.4]
  assign valid_4_40 = io_inValid_40 & _T_19314; // @[Switch.scala 30:36:@1419.4]
  assign _T_19317 = io_inAddr_41 == 6'h4; // @[Switch.scala 30:53:@1421.4]
  assign valid_4_41 = io_inValid_41 & _T_19317; // @[Switch.scala 30:36:@1422.4]
  assign _T_19320 = io_inAddr_42 == 6'h4; // @[Switch.scala 30:53:@1424.4]
  assign valid_4_42 = io_inValid_42 & _T_19320; // @[Switch.scala 30:36:@1425.4]
  assign _T_19323 = io_inAddr_43 == 6'h4; // @[Switch.scala 30:53:@1427.4]
  assign valid_4_43 = io_inValid_43 & _T_19323; // @[Switch.scala 30:36:@1428.4]
  assign _T_19326 = io_inAddr_44 == 6'h4; // @[Switch.scala 30:53:@1430.4]
  assign valid_4_44 = io_inValid_44 & _T_19326; // @[Switch.scala 30:36:@1431.4]
  assign _T_19329 = io_inAddr_45 == 6'h4; // @[Switch.scala 30:53:@1433.4]
  assign valid_4_45 = io_inValid_45 & _T_19329; // @[Switch.scala 30:36:@1434.4]
  assign _T_19332 = io_inAddr_46 == 6'h4; // @[Switch.scala 30:53:@1436.4]
  assign valid_4_46 = io_inValid_46 & _T_19332; // @[Switch.scala 30:36:@1437.4]
  assign _T_19335 = io_inAddr_47 == 6'h4; // @[Switch.scala 30:53:@1439.4]
  assign valid_4_47 = io_inValid_47 & _T_19335; // @[Switch.scala 30:36:@1440.4]
  assign _T_19338 = io_inAddr_48 == 6'h4; // @[Switch.scala 30:53:@1442.4]
  assign valid_4_48 = io_inValid_48 & _T_19338; // @[Switch.scala 30:36:@1443.4]
  assign _T_19341 = io_inAddr_49 == 6'h4; // @[Switch.scala 30:53:@1445.4]
  assign valid_4_49 = io_inValid_49 & _T_19341; // @[Switch.scala 30:36:@1446.4]
  assign _T_19344 = io_inAddr_50 == 6'h4; // @[Switch.scala 30:53:@1448.4]
  assign valid_4_50 = io_inValid_50 & _T_19344; // @[Switch.scala 30:36:@1449.4]
  assign _T_19347 = io_inAddr_51 == 6'h4; // @[Switch.scala 30:53:@1451.4]
  assign valid_4_51 = io_inValid_51 & _T_19347; // @[Switch.scala 30:36:@1452.4]
  assign _T_19350 = io_inAddr_52 == 6'h4; // @[Switch.scala 30:53:@1454.4]
  assign valid_4_52 = io_inValid_52 & _T_19350; // @[Switch.scala 30:36:@1455.4]
  assign _T_19353 = io_inAddr_53 == 6'h4; // @[Switch.scala 30:53:@1457.4]
  assign valid_4_53 = io_inValid_53 & _T_19353; // @[Switch.scala 30:36:@1458.4]
  assign _T_19356 = io_inAddr_54 == 6'h4; // @[Switch.scala 30:53:@1460.4]
  assign valid_4_54 = io_inValid_54 & _T_19356; // @[Switch.scala 30:36:@1461.4]
  assign _T_19359 = io_inAddr_55 == 6'h4; // @[Switch.scala 30:53:@1463.4]
  assign valid_4_55 = io_inValid_55 & _T_19359; // @[Switch.scala 30:36:@1464.4]
  assign _T_19362 = io_inAddr_56 == 6'h4; // @[Switch.scala 30:53:@1466.4]
  assign valid_4_56 = io_inValid_56 & _T_19362; // @[Switch.scala 30:36:@1467.4]
  assign _T_19365 = io_inAddr_57 == 6'h4; // @[Switch.scala 30:53:@1469.4]
  assign valid_4_57 = io_inValid_57 & _T_19365; // @[Switch.scala 30:36:@1470.4]
  assign _T_19368 = io_inAddr_58 == 6'h4; // @[Switch.scala 30:53:@1472.4]
  assign valid_4_58 = io_inValid_58 & _T_19368; // @[Switch.scala 30:36:@1473.4]
  assign _T_19371 = io_inAddr_59 == 6'h4; // @[Switch.scala 30:53:@1475.4]
  assign valid_4_59 = io_inValid_59 & _T_19371; // @[Switch.scala 30:36:@1476.4]
  assign _T_19374 = io_inAddr_60 == 6'h4; // @[Switch.scala 30:53:@1478.4]
  assign valid_4_60 = io_inValid_60 & _T_19374; // @[Switch.scala 30:36:@1479.4]
  assign _T_19377 = io_inAddr_61 == 6'h4; // @[Switch.scala 30:53:@1481.4]
  assign valid_4_61 = io_inValid_61 & _T_19377; // @[Switch.scala 30:36:@1482.4]
  assign _T_19380 = io_inAddr_62 == 6'h4; // @[Switch.scala 30:53:@1484.4]
  assign valid_4_62 = io_inValid_62 & _T_19380; // @[Switch.scala 30:36:@1485.4]
  assign _T_19383 = io_inAddr_63 == 6'h4; // @[Switch.scala 30:53:@1487.4]
  assign valid_4_63 = io_inValid_63 & _T_19383; // @[Switch.scala 30:36:@1488.4]
  assign _T_19449 = valid_4_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@1490.4]
  assign _T_19450 = valid_4_61 ? 6'h3d : _T_19449; // @[Mux.scala 31:69:@1491.4]
  assign _T_19451 = valid_4_60 ? 6'h3c : _T_19450; // @[Mux.scala 31:69:@1492.4]
  assign _T_19452 = valid_4_59 ? 6'h3b : _T_19451; // @[Mux.scala 31:69:@1493.4]
  assign _T_19453 = valid_4_58 ? 6'h3a : _T_19452; // @[Mux.scala 31:69:@1494.4]
  assign _T_19454 = valid_4_57 ? 6'h39 : _T_19453; // @[Mux.scala 31:69:@1495.4]
  assign _T_19455 = valid_4_56 ? 6'h38 : _T_19454; // @[Mux.scala 31:69:@1496.4]
  assign _T_19456 = valid_4_55 ? 6'h37 : _T_19455; // @[Mux.scala 31:69:@1497.4]
  assign _T_19457 = valid_4_54 ? 6'h36 : _T_19456; // @[Mux.scala 31:69:@1498.4]
  assign _T_19458 = valid_4_53 ? 6'h35 : _T_19457; // @[Mux.scala 31:69:@1499.4]
  assign _T_19459 = valid_4_52 ? 6'h34 : _T_19458; // @[Mux.scala 31:69:@1500.4]
  assign _T_19460 = valid_4_51 ? 6'h33 : _T_19459; // @[Mux.scala 31:69:@1501.4]
  assign _T_19461 = valid_4_50 ? 6'h32 : _T_19460; // @[Mux.scala 31:69:@1502.4]
  assign _T_19462 = valid_4_49 ? 6'h31 : _T_19461; // @[Mux.scala 31:69:@1503.4]
  assign _T_19463 = valid_4_48 ? 6'h30 : _T_19462; // @[Mux.scala 31:69:@1504.4]
  assign _T_19464 = valid_4_47 ? 6'h2f : _T_19463; // @[Mux.scala 31:69:@1505.4]
  assign _T_19465 = valid_4_46 ? 6'h2e : _T_19464; // @[Mux.scala 31:69:@1506.4]
  assign _T_19466 = valid_4_45 ? 6'h2d : _T_19465; // @[Mux.scala 31:69:@1507.4]
  assign _T_19467 = valid_4_44 ? 6'h2c : _T_19466; // @[Mux.scala 31:69:@1508.4]
  assign _T_19468 = valid_4_43 ? 6'h2b : _T_19467; // @[Mux.scala 31:69:@1509.4]
  assign _T_19469 = valid_4_42 ? 6'h2a : _T_19468; // @[Mux.scala 31:69:@1510.4]
  assign _T_19470 = valid_4_41 ? 6'h29 : _T_19469; // @[Mux.scala 31:69:@1511.4]
  assign _T_19471 = valid_4_40 ? 6'h28 : _T_19470; // @[Mux.scala 31:69:@1512.4]
  assign _T_19472 = valid_4_39 ? 6'h27 : _T_19471; // @[Mux.scala 31:69:@1513.4]
  assign _T_19473 = valid_4_38 ? 6'h26 : _T_19472; // @[Mux.scala 31:69:@1514.4]
  assign _T_19474 = valid_4_37 ? 6'h25 : _T_19473; // @[Mux.scala 31:69:@1515.4]
  assign _T_19475 = valid_4_36 ? 6'h24 : _T_19474; // @[Mux.scala 31:69:@1516.4]
  assign _T_19476 = valid_4_35 ? 6'h23 : _T_19475; // @[Mux.scala 31:69:@1517.4]
  assign _T_19477 = valid_4_34 ? 6'h22 : _T_19476; // @[Mux.scala 31:69:@1518.4]
  assign _T_19478 = valid_4_33 ? 6'h21 : _T_19477; // @[Mux.scala 31:69:@1519.4]
  assign _T_19479 = valid_4_32 ? 6'h20 : _T_19478; // @[Mux.scala 31:69:@1520.4]
  assign _T_19480 = valid_4_31 ? 6'h1f : _T_19479; // @[Mux.scala 31:69:@1521.4]
  assign _T_19481 = valid_4_30 ? 6'h1e : _T_19480; // @[Mux.scala 31:69:@1522.4]
  assign _T_19482 = valid_4_29 ? 6'h1d : _T_19481; // @[Mux.scala 31:69:@1523.4]
  assign _T_19483 = valid_4_28 ? 6'h1c : _T_19482; // @[Mux.scala 31:69:@1524.4]
  assign _T_19484 = valid_4_27 ? 6'h1b : _T_19483; // @[Mux.scala 31:69:@1525.4]
  assign _T_19485 = valid_4_26 ? 6'h1a : _T_19484; // @[Mux.scala 31:69:@1526.4]
  assign _T_19486 = valid_4_25 ? 6'h19 : _T_19485; // @[Mux.scala 31:69:@1527.4]
  assign _T_19487 = valid_4_24 ? 6'h18 : _T_19486; // @[Mux.scala 31:69:@1528.4]
  assign _T_19488 = valid_4_23 ? 6'h17 : _T_19487; // @[Mux.scala 31:69:@1529.4]
  assign _T_19489 = valid_4_22 ? 6'h16 : _T_19488; // @[Mux.scala 31:69:@1530.4]
  assign _T_19490 = valid_4_21 ? 6'h15 : _T_19489; // @[Mux.scala 31:69:@1531.4]
  assign _T_19491 = valid_4_20 ? 6'h14 : _T_19490; // @[Mux.scala 31:69:@1532.4]
  assign _T_19492 = valid_4_19 ? 6'h13 : _T_19491; // @[Mux.scala 31:69:@1533.4]
  assign _T_19493 = valid_4_18 ? 6'h12 : _T_19492; // @[Mux.scala 31:69:@1534.4]
  assign _T_19494 = valid_4_17 ? 6'h11 : _T_19493; // @[Mux.scala 31:69:@1535.4]
  assign _T_19495 = valid_4_16 ? 6'h10 : _T_19494; // @[Mux.scala 31:69:@1536.4]
  assign _T_19496 = valid_4_15 ? 6'hf : _T_19495; // @[Mux.scala 31:69:@1537.4]
  assign _T_19497 = valid_4_14 ? 6'he : _T_19496; // @[Mux.scala 31:69:@1538.4]
  assign _T_19498 = valid_4_13 ? 6'hd : _T_19497; // @[Mux.scala 31:69:@1539.4]
  assign _T_19499 = valid_4_12 ? 6'hc : _T_19498; // @[Mux.scala 31:69:@1540.4]
  assign _T_19500 = valid_4_11 ? 6'hb : _T_19499; // @[Mux.scala 31:69:@1541.4]
  assign _T_19501 = valid_4_10 ? 6'ha : _T_19500; // @[Mux.scala 31:69:@1542.4]
  assign _T_19502 = valid_4_9 ? 6'h9 : _T_19501; // @[Mux.scala 31:69:@1543.4]
  assign _T_19503 = valid_4_8 ? 6'h8 : _T_19502; // @[Mux.scala 31:69:@1544.4]
  assign _T_19504 = valid_4_7 ? 6'h7 : _T_19503; // @[Mux.scala 31:69:@1545.4]
  assign _T_19505 = valid_4_6 ? 6'h6 : _T_19504; // @[Mux.scala 31:69:@1546.4]
  assign _T_19506 = valid_4_5 ? 6'h5 : _T_19505; // @[Mux.scala 31:69:@1547.4]
  assign _T_19507 = valid_4_4 ? 6'h4 : _T_19506; // @[Mux.scala 31:69:@1548.4]
  assign _T_19508 = valid_4_3 ? 6'h3 : _T_19507; // @[Mux.scala 31:69:@1549.4]
  assign _T_19509 = valid_4_2 ? 6'h2 : _T_19508; // @[Mux.scala 31:69:@1550.4]
  assign _T_19510 = valid_4_1 ? 6'h1 : _T_19509; // @[Mux.scala 31:69:@1551.4]
  assign select_4 = valid_4_0 ? 6'h0 : _T_19510; // @[Mux.scala 31:69:@1552.4]
  assign _GEN_257 = 6'h1 == select_4 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_258 = 6'h2 == select_4 ? io_inData_2 : _GEN_257; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_259 = 6'h3 == select_4 ? io_inData_3 : _GEN_258; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_260 = 6'h4 == select_4 ? io_inData_4 : _GEN_259; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_261 = 6'h5 == select_4 ? io_inData_5 : _GEN_260; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_262 = 6'h6 == select_4 ? io_inData_6 : _GEN_261; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_263 = 6'h7 == select_4 ? io_inData_7 : _GEN_262; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_264 = 6'h8 == select_4 ? io_inData_8 : _GEN_263; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_265 = 6'h9 == select_4 ? io_inData_9 : _GEN_264; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_266 = 6'ha == select_4 ? io_inData_10 : _GEN_265; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_267 = 6'hb == select_4 ? io_inData_11 : _GEN_266; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_268 = 6'hc == select_4 ? io_inData_12 : _GEN_267; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_269 = 6'hd == select_4 ? io_inData_13 : _GEN_268; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_270 = 6'he == select_4 ? io_inData_14 : _GEN_269; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_271 = 6'hf == select_4 ? io_inData_15 : _GEN_270; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_272 = 6'h10 == select_4 ? io_inData_16 : _GEN_271; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_273 = 6'h11 == select_4 ? io_inData_17 : _GEN_272; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_274 = 6'h12 == select_4 ? io_inData_18 : _GEN_273; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_275 = 6'h13 == select_4 ? io_inData_19 : _GEN_274; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_276 = 6'h14 == select_4 ? io_inData_20 : _GEN_275; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_277 = 6'h15 == select_4 ? io_inData_21 : _GEN_276; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_278 = 6'h16 == select_4 ? io_inData_22 : _GEN_277; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_279 = 6'h17 == select_4 ? io_inData_23 : _GEN_278; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_280 = 6'h18 == select_4 ? io_inData_24 : _GEN_279; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_281 = 6'h19 == select_4 ? io_inData_25 : _GEN_280; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_282 = 6'h1a == select_4 ? io_inData_26 : _GEN_281; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_283 = 6'h1b == select_4 ? io_inData_27 : _GEN_282; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_284 = 6'h1c == select_4 ? io_inData_28 : _GEN_283; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_285 = 6'h1d == select_4 ? io_inData_29 : _GEN_284; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_286 = 6'h1e == select_4 ? io_inData_30 : _GEN_285; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_287 = 6'h1f == select_4 ? io_inData_31 : _GEN_286; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_288 = 6'h20 == select_4 ? io_inData_32 : _GEN_287; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_289 = 6'h21 == select_4 ? io_inData_33 : _GEN_288; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_290 = 6'h22 == select_4 ? io_inData_34 : _GEN_289; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_291 = 6'h23 == select_4 ? io_inData_35 : _GEN_290; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_292 = 6'h24 == select_4 ? io_inData_36 : _GEN_291; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_293 = 6'h25 == select_4 ? io_inData_37 : _GEN_292; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_294 = 6'h26 == select_4 ? io_inData_38 : _GEN_293; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_295 = 6'h27 == select_4 ? io_inData_39 : _GEN_294; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_296 = 6'h28 == select_4 ? io_inData_40 : _GEN_295; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_297 = 6'h29 == select_4 ? io_inData_41 : _GEN_296; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_298 = 6'h2a == select_4 ? io_inData_42 : _GEN_297; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_299 = 6'h2b == select_4 ? io_inData_43 : _GEN_298; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_300 = 6'h2c == select_4 ? io_inData_44 : _GEN_299; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_301 = 6'h2d == select_4 ? io_inData_45 : _GEN_300; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_302 = 6'h2e == select_4 ? io_inData_46 : _GEN_301; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_303 = 6'h2f == select_4 ? io_inData_47 : _GEN_302; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_304 = 6'h30 == select_4 ? io_inData_48 : _GEN_303; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_305 = 6'h31 == select_4 ? io_inData_49 : _GEN_304; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_306 = 6'h32 == select_4 ? io_inData_50 : _GEN_305; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_307 = 6'h33 == select_4 ? io_inData_51 : _GEN_306; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_308 = 6'h34 == select_4 ? io_inData_52 : _GEN_307; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_309 = 6'h35 == select_4 ? io_inData_53 : _GEN_308; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_310 = 6'h36 == select_4 ? io_inData_54 : _GEN_309; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_311 = 6'h37 == select_4 ? io_inData_55 : _GEN_310; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_312 = 6'h38 == select_4 ? io_inData_56 : _GEN_311; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_313 = 6'h39 == select_4 ? io_inData_57 : _GEN_312; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_314 = 6'h3a == select_4 ? io_inData_58 : _GEN_313; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_315 = 6'h3b == select_4 ? io_inData_59 : _GEN_314; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_316 = 6'h3c == select_4 ? io_inData_60 : _GEN_315; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_317 = 6'h3d == select_4 ? io_inData_61 : _GEN_316; // @[Switch.scala 33:19:@1554.4]
  assign _GEN_318 = 6'h3e == select_4 ? io_inData_62 : _GEN_317; // @[Switch.scala 33:19:@1554.4]
  assign _T_19519 = {valid_4_7,valid_4_6,valid_4_5,valid_4_4,valid_4_3,valid_4_2,valid_4_1,valid_4_0}; // @[Switch.scala 34:32:@1561.4]
  assign _T_19527 = {valid_4_15,valid_4_14,valid_4_13,valid_4_12,valid_4_11,valid_4_10,valid_4_9,valid_4_8,_T_19519}; // @[Switch.scala 34:32:@1569.4]
  assign _T_19534 = {valid_4_23,valid_4_22,valid_4_21,valid_4_20,valid_4_19,valid_4_18,valid_4_17,valid_4_16}; // @[Switch.scala 34:32:@1576.4]
  assign _T_19543 = {valid_4_31,valid_4_30,valid_4_29,valid_4_28,valid_4_27,valid_4_26,valid_4_25,valid_4_24,_T_19534,_T_19527}; // @[Switch.scala 34:32:@1585.4]
  assign _T_19550 = {valid_4_39,valid_4_38,valid_4_37,valid_4_36,valid_4_35,valid_4_34,valid_4_33,valid_4_32}; // @[Switch.scala 34:32:@1592.4]
  assign _T_19558 = {valid_4_47,valid_4_46,valid_4_45,valid_4_44,valid_4_43,valid_4_42,valid_4_41,valid_4_40,_T_19550}; // @[Switch.scala 34:32:@1600.4]
  assign _T_19565 = {valid_4_55,valid_4_54,valid_4_53,valid_4_52,valid_4_51,valid_4_50,valid_4_49,valid_4_48}; // @[Switch.scala 34:32:@1607.4]
  assign _T_19574 = {valid_4_63,valid_4_62,valid_4_61,valid_4_60,valid_4_59,valid_4_58,valid_4_57,valid_4_56,_T_19565,_T_19558}; // @[Switch.scala 34:32:@1616.4]
  assign _T_19575 = {_T_19574,_T_19543}; // @[Switch.scala 34:32:@1617.4]
  assign _T_19579 = io_inAddr_0 == 6'h5; // @[Switch.scala 30:53:@1620.4]
  assign valid_5_0 = io_inValid_0 & _T_19579; // @[Switch.scala 30:36:@1621.4]
  assign _T_19582 = io_inAddr_1 == 6'h5; // @[Switch.scala 30:53:@1623.4]
  assign valid_5_1 = io_inValid_1 & _T_19582; // @[Switch.scala 30:36:@1624.4]
  assign _T_19585 = io_inAddr_2 == 6'h5; // @[Switch.scala 30:53:@1626.4]
  assign valid_5_2 = io_inValid_2 & _T_19585; // @[Switch.scala 30:36:@1627.4]
  assign _T_19588 = io_inAddr_3 == 6'h5; // @[Switch.scala 30:53:@1629.4]
  assign valid_5_3 = io_inValid_3 & _T_19588; // @[Switch.scala 30:36:@1630.4]
  assign _T_19591 = io_inAddr_4 == 6'h5; // @[Switch.scala 30:53:@1632.4]
  assign valid_5_4 = io_inValid_4 & _T_19591; // @[Switch.scala 30:36:@1633.4]
  assign _T_19594 = io_inAddr_5 == 6'h5; // @[Switch.scala 30:53:@1635.4]
  assign valid_5_5 = io_inValid_5 & _T_19594; // @[Switch.scala 30:36:@1636.4]
  assign _T_19597 = io_inAddr_6 == 6'h5; // @[Switch.scala 30:53:@1638.4]
  assign valid_5_6 = io_inValid_6 & _T_19597; // @[Switch.scala 30:36:@1639.4]
  assign _T_19600 = io_inAddr_7 == 6'h5; // @[Switch.scala 30:53:@1641.4]
  assign valid_5_7 = io_inValid_7 & _T_19600; // @[Switch.scala 30:36:@1642.4]
  assign _T_19603 = io_inAddr_8 == 6'h5; // @[Switch.scala 30:53:@1644.4]
  assign valid_5_8 = io_inValid_8 & _T_19603; // @[Switch.scala 30:36:@1645.4]
  assign _T_19606 = io_inAddr_9 == 6'h5; // @[Switch.scala 30:53:@1647.4]
  assign valid_5_9 = io_inValid_9 & _T_19606; // @[Switch.scala 30:36:@1648.4]
  assign _T_19609 = io_inAddr_10 == 6'h5; // @[Switch.scala 30:53:@1650.4]
  assign valid_5_10 = io_inValid_10 & _T_19609; // @[Switch.scala 30:36:@1651.4]
  assign _T_19612 = io_inAddr_11 == 6'h5; // @[Switch.scala 30:53:@1653.4]
  assign valid_5_11 = io_inValid_11 & _T_19612; // @[Switch.scala 30:36:@1654.4]
  assign _T_19615 = io_inAddr_12 == 6'h5; // @[Switch.scala 30:53:@1656.4]
  assign valid_5_12 = io_inValid_12 & _T_19615; // @[Switch.scala 30:36:@1657.4]
  assign _T_19618 = io_inAddr_13 == 6'h5; // @[Switch.scala 30:53:@1659.4]
  assign valid_5_13 = io_inValid_13 & _T_19618; // @[Switch.scala 30:36:@1660.4]
  assign _T_19621 = io_inAddr_14 == 6'h5; // @[Switch.scala 30:53:@1662.4]
  assign valid_5_14 = io_inValid_14 & _T_19621; // @[Switch.scala 30:36:@1663.4]
  assign _T_19624 = io_inAddr_15 == 6'h5; // @[Switch.scala 30:53:@1665.4]
  assign valid_5_15 = io_inValid_15 & _T_19624; // @[Switch.scala 30:36:@1666.4]
  assign _T_19627 = io_inAddr_16 == 6'h5; // @[Switch.scala 30:53:@1668.4]
  assign valid_5_16 = io_inValid_16 & _T_19627; // @[Switch.scala 30:36:@1669.4]
  assign _T_19630 = io_inAddr_17 == 6'h5; // @[Switch.scala 30:53:@1671.4]
  assign valid_5_17 = io_inValid_17 & _T_19630; // @[Switch.scala 30:36:@1672.4]
  assign _T_19633 = io_inAddr_18 == 6'h5; // @[Switch.scala 30:53:@1674.4]
  assign valid_5_18 = io_inValid_18 & _T_19633; // @[Switch.scala 30:36:@1675.4]
  assign _T_19636 = io_inAddr_19 == 6'h5; // @[Switch.scala 30:53:@1677.4]
  assign valid_5_19 = io_inValid_19 & _T_19636; // @[Switch.scala 30:36:@1678.4]
  assign _T_19639 = io_inAddr_20 == 6'h5; // @[Switch.scala 30:53:@1680.4]
  assign valid_5_20 = io_inValid_20 & _T_19639; // @[Switch.scala 30:36:@1681.4]
  assign _T_19642 = io_inAddr_21 == 6'h5; // @[Switch.scala 30:53:@1683.4]
  assign valid_5_21 = io_inValid_21 & _T_19642; // @[Switch.scala 30:36:@1684.4]
  assign _T_19645 = io_inAddr_22 == 6'h5; // @[Switch.scala 30:53:@1686.4]
  assign valid_5_22 = io_inValid_22 & _T_19645; // @[Switch.scala 30:36:@1687.4]
  assign _T_19648 = io_inAddr_23 == 6'h5; // @[Switch.scala 30:53:@1689.4]
  assign valid_5_23 = io_inValid_23 & _T_19648; // @[Switch.scala 30:36:@1690.4]
  assign _T_19651 = io_inAddr_24 == 6'h5; // @[Switch.scala 30:53:@1692.4]
  assign valid_5_24 = io_inValid_24 & _T_19651; // @[Switch.scala 30:36:@1693.4]
  assign _T_19654 = io_inAddr_25 == 6'h5; // @[Switch.scala 30:53:@1695.4]
  assign valid_5_25 = io_inValid_25 & _T_19654; // @[Switch.scala 30:36:@1696.4]
  assign _T_19657 = io_inAddr_26 == 6'h5; // @[Switch.scala 30:53:@1698.4]
  assign valid_5_26 = io_inValid_26 & _T_19657; // @[Switch.scala 30:36:@1699.4]
  assign _T_19660 = io_inAddr_27 == 6'h5; // @[Switch.scala 30:53:@1701.4]
  assign valid_5_27 = io_inValid_27 & _T_19660; // @[Switch.scala 30:36:@1702.4]
  assign _T_19663 = io_inAddr_28 == 6'h5; // @[Switch.scala 30:53:@1704.4]
  assign valid_5_28 = io_inValid_28 & _T_19663; // @[Switch.scala 30:36:@1705.4]
  assign _T_19666 = io_inAddr_29 == 6'h5; // @[Switch.scala 30:53:@1707.4]
  assign valid_5_29 = io_inValid_29 & _T_19666; // @[Switch.scala 30:36:@1708.4]
  assign _T_19669 = io_inAddr_30 == 6'h5; // @[Switch.scala 30:53:@1710.4]
  assign valid_5_30 = io_inValid_30 & _T_19669; // @[Switch.scala 30:36:@1711.4]
  assign _T_19672 = io_inAddr_31 == 6'h5; // @[Switch.scala 30:53:@1713.4]
  assign valid_5_31 = io_inValid_31 & _T_19672; // @[Switch.scala 30:36:@1714.4]
  assign _T_19675 = io_inAddr_32 == 6'h5; // @[Switch.scala 30:53:@1716.4]
  assign valid_5_32 = io_inValid_32 & _T_19675; // @[Switch.scala 30:36:@1717.4]
  assign _T_19678 = io_inAddr_33 == 6'h5; // @[Switch.scala 30:53:@1719.4]
  assign valid_5_33 = io_inValid_33 & _T_19678; // @[Switch.scala 30:36:@1720.4]
  assign _T_19681 = io_inAddr_34 == 6'h5; // @[Switch.scala 30:53:@1722.4]
  assign valid_5_34 = io_inValid_34 & _T_19681; // @[Switch.scala 30:36:@1723.4]
  assign _T_19684 = io_inAddr_35 == 6'h5; // @[Switch.scala 30:53:@1725.4]
  assign valid_5_35 = io_inValid_35 & _T_19684; // @[Switch.scala 30:36:@1726.4]
  assign _T_19687 = io_inAddr_36 == 6'h5; // @[Switch.scala 30:53:@1728.4]
  assign valid_5_36 = io_inValid_36 & _T_19687; // @[Switch.scala 30:36:@1729.4]
  assign _T_19690 = io_inAddr_37 == 6'h5; // @[Switch.scala 30:53:@1731.4]
  assign valid_5_37 = io_inValid_37 & _T_19690; // @[Switch.scala 30:36:@1732.4]
  assign _T_19693 = io_inAddr_38 == 6'h5; // @[Switch.scala 30:53:@1734.4]
  assign valid_5_38 = io_inValid_38 & _T_19693; // @[Switch.scala 30:36:@1735.4]
  assign _T_19696 = io_inAddr_39 == 6'h5; // @[Switch.scala 30:53:@1737.4]
  assign valid_5_39 = io_inValid_39 & _T_19696; // @[Switch.scala 30:36:@1738.4]
  assign _T_19699 = io_inAddr_40 == 6'h5; // @[Switch.scala 30:53:@1740.4]
  assign valid_5_40 = io_inValid_40 & _T_19699; // @[Switch.scala 30:36:@1741.4]
  assign _T_19702 = io_inAddr_41 == 6'h5; // @[Switch.scala 30:53:@1743.4]
  assign valid_5_41 = io_inValid_41 & _T_19702; // @[Switch.scala 30:36:@1744.4]
  assign _T_19705 = io_inAddr_42 == 6'h5; // @[Switch.scala 30:53:@1746.4]
  assign valid_5_42 = io_inValid_42 & _T_19705; // @[Switch.scala 30:36:@1747.4]
  assign _T_19708 = io_inAddr_43 == 6'h5; // @[Switch.scala 30:53:@1749.4]
  assign valid_5_43 = io_inValid_43 & _T_19708; // @[Switch.scala 30:36:@1750.4]
  assign _T_19711 = io_inAddr_44 == 6'h5; // @[Switch.scala 30:53:@1752.4]
  assign valid_5_44 = io_inValid_44 & _T_19711; // @[Switch.scala 30:36:@1753.4]
  assign _T_19714 = io_inAddr_45 == 6'h5; // @[Switch.scala 30:53:@1755.4]
  assign valid_5_45 = io_inValid_45 & _T_19714; // @[Switch.scala 30:36:@1756.4]
  assign _T_19717 = io_inAddr_46 == 6'h5; // @[Switch.scala 30:53:@1758.4]
  assign valid_5_46 = io_inValid_46 & _T_19717; // @[Switch.scala 30:36:@1759.4]
  assign _T_19720 = io_inAddr_47 == 6'h5; // @[Switch.scala 30:53:@1761.4]
  assign valid_5_47 = io_inValid_47 & _T_19720; // @[Switch.scala 30:36:@1762.4]
  assign _T_19723 = io_inAddr_48 == 6'h5; // @[Switch.scala 30:53:@1764.4]
  assign valid_5_48 = io_inValid_48 & _T_19723; // @[Switch.scala 30:36:@1765.4]
  assign _T_19726 = io_inAddr_49 == 6'h5; // @[Switch.scala 30:53:@1767.4]
  assign valid_5_49 = io_inValid_49 & _T_19726; // @[Switch.scala 30:36:@1768.4]
  assign _T_19729 = io_inAddr_50 == 6'h5; // @[Switch.scala 30:53:@1770.4]
  assign valid_5_50 = io_inValid_50 & _T_19729; // @[Switch.scala 30:36:@1771.4]
  assign _T_19732 = io_inAddr_51 == 6'h5; // @[Switch.scala 30:53:@1773.4]
  assign valid_5_51 = io_inValid_51 & _T_19732; // @[Switch.scala 30:36:@1774.4]
  assign _T_19735 = io_inAddr_52 == 6'h5; // @[Switch.scala 30:53:@1776.4]
  assign valid_5_52 = io_inValid_52 & _T_19735; // @[Switch.scala 30:36:@1777.4]
  assign _T_19738 = io_inAddr_53 == 6'h5; // @[Switch.scala 30:53:@1779.4]
  assign valid_5_53 = io_inValid_53 & _T_19738; // @[Switch.scala 30:36:@1780.4]
  assign _T_19741 = io_inAddr_54 == 6'h5; // @[Switch.scala 30:53:@1782.4]
  assign valid_5_54 = io_inValid_54 & _T_19741; // @[Switch.scala 30:36:@1783.4]
  assign _T_19744 = io_inAddr_55 == 6'h5; // @[Switch.scala 30:53:@1785.4]
  assign valid_5_55 = io_inValid_55 & _T_19744; // @[Switch.scala 30:36:@1786.4]
  assign _T_19747 = io_inAddr_56 == 6'h5; // @[Switch.scala 30:53:@1788.4]
  assign valid_5_56 = io_inValid_56 & _T_19747; // @[Switch.scala 30:36:@1789.4]
  assign _T_19750 = io_inAddr_57 == 6'h5; // @[Switch.scala 30:53:@1791.4]
  assign valid_5_57 = io_inValid_57 & _T_19750; // @[Switch.scala 30:36:@1792.4]
  assign _T_19753 = io_inAddr_58 == 6'h5; // @[Switch.scala 30:53:@1794.4]
  assign valid_5_58 = io_inValid_58 & _T_19753; // @[Switch.scala 30:36:@1795.4]
  assign _T_19756 = io_inAddr_59 == 6'h5; // @[Switch.scala 30:53:@1797.4]
  assign valid_5_59 = io_inValid_59 & _T_19756; // @[Switch.scala 30:36:@1798.4]
  assign _T_19759 = io_inAddr_60 == 6'h5; // @[Switch.scala 30:53:@1800.4]
  assign valid_5_60 = io_inValid_60 & _T_19759; // @[Switch.scala 30:36:@1801.4]
  assign _T_19762 = io_inAddr_61 == 6'h5; // @[Switch.scala 30:53:@1803.4]
  assign valid_5_61 = io_inValid_61 & _T_19762; // @[Switch.scala 30:36:@1804.4]
  assign _T_19765 = io_inAddr_62 == 6'h5; // @[Switch.scala 30:53:@1806.4]
  assign valid_5_62 = io_inValid_62 & _T_19765; // @[Switch.scala 30:36:@1807.4]
  assign _T_19768 = io_inAddr_63 == 6'h5; // @[Switch.scala 30:53:@1809.4]
  assign valid_5_63 = io_inValid_63 & _T_19768; // @[Switch.scala 30:36:@1810.4]
  assign _T_19834 = valid_5_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@1812.4]
  assign _T_19835 = valid_5_61 ? 6'h3d : _T_19834; // @[Mux.scala 31:69:@1813.4]
  assign _T_19836 = valid_5_60 ? 6'h3c : _T_19835; // @[Mux.scala 31:69:@1814.4]
  assign _T_19837 = valid_5_59 ? 6'h3b : _T_19836; // @[Mux.scala 31:69:@1815.4]
  assign _T_19838 = valid_5_58 ? 6'h3a : _T_19837; // @[Mux.scala 31:69:@1816.4]
  assign _T_19839 = valid_5_57 ? 6'h39 : _T_19838; // @[Mux.scala 31:69:@1817.4]
  assign _T_19840 = valid_5_56 ? 6'h38 : _T_19839; // @[Mux.scala 31:69:@1818.4]
  assign _T_19841 = valid_5_55 ? 6'h37 : _T_19840; // @[Mux.scala 31:69:@1819.4]
  assign _T_19842 = valid_5_54 ? 6'h36 : _T_19841; // @[Mux.scala 31:69:@1820.4]
  assign _T_19843 = valid_5_53 ? 6'h35 : _T_19842; // @[Mux.scala 31:69:@1821.4]
  assign _T_19844 = valid_5_52 ? 6'h34 : _T_19843; // @[Mux.scala 31:69:@1822.4]
  assign _T_19845 = valid_5_51 ? 6'h33 : _T_19844; // @[Mux.scala 31:69:@1823.4]
  assign _T_19846 = valid_5_50 ? 6'h32 : _T_19845; // @[Mux.scala 31:69:@1824.4]
  assign _T_19847 = valid_5_49 ? 6'h31 : _T_19846; // @[Mux.scala 31:69:@1825.4]
  assign _T_19848 = valid_5_48 ? 6'h30 : _T_19847; // @[Mux.scala 31:69:@1826.4]
  assign _T_19849 = valid_5_47 ? 6'h2f : _T_19848; // @[Mux.scala 31:69:@1827.4]
  assign _T_19850 = valid_5_46 ? 6'h2e : _T_19849; // @[Mux.scala 31:69:@1828.4]
  assign _T_19851 = valid_5_45 ? 6'h2d : _T_19850; // @[Mux.scala 31:69:@1829.4]
  assign _T_19852 = valid_5_44 ? 6'h2c : _T_19851; // @[Mux.scala 31:69:@1830.4]
  assign _T_19853 = valid_5_43 ? 6'h2b : _T_19852; // @[Mux.scala 31:69:@1831.4]
  assign _T_19854 = valid_5_42 ? 6'h2a : _T_19853; // @[Mux.scala 31:69:@1832.4]
  assign _T_19855 = valid_5_41 ? 6'h29 : _T_19854; // @[Mux.scala 31:69:@1833.4]
  assign _T_19856 = valid_5_40 ? 6'h28 : _T_19855; // @[Mux.scala 31:69:@1834.4]
  assign _T_19857 = valid_5_39 ? 6'h27 : _T_19856; // @[Mux.scala 31:69:@1835.4]
  assign _T_19858 = valid_5_38 ? 6'h26 : _T_19857; // @[Mux.scala 31:69:@1836.4]
  assign _T_19859 = valid_5_37 ? 6'h25 : _T_19858; // @[Mux.scala 31:69:@1837.4]
  assign _T_19860 = valid_5_36 ? 6'h24 : _T_19859; // @[Mux.scala 31:69:@1838.4]
  assign _T_19861 = valid_5_35 ? 6'h23 : _T_19860; // @[Mux.scala 31:69:@1839.4]
  assign _T_19862 = valid_5_34 ? 6'h22 : _T_19861; // @[Mux.scala 31:69:@1840.4]
  assign _T_19863 = valid_5_33 ? 6'h21 : _T_19862; // @[Mux.scala 31:69:@1841.4]
  assign _T_19864 = valid_5_32 ? 6'h20 : _T_19863; // @[Mux.scala 31:69:@1842.4]
  assign _T_19865 = valid_5_31 ? 6'h1f : _T_19864; // @[Mux.scala 31:69:@1843.4]
  assign _T_19866 = valid_5_30 ? 6'h1e : _T_19865; // @[Mux.scala 31:69:@1844.4]
  assign _T_19867 = valid_5_29 ? 6'h1d : _T_19866; // @[Mux.scala 31:69:@1845.4]
  assign _T_19868 = valid_5_28 ? 6'h1c : _T_19867; // @[Mux.scala 31:69:@1846.4]
  assign _T_19869 = valid_5_27 ? 6'h1b : _T_19868; // @[Mux.scala 31:69:@1847.4]
  assign _T_19870 = valid_5_26 ? 6'h1a : _T_19869; // @[Mux.scala 31:69:@1848.4]
  assign _T_19871 = valid_5_25 ? 6'h19 : _T_19870; // @[Mux.scala 31:69:@1849.4]
  assign _T_19872 = valid_5_24 ? 6'h18 : _T_19871; // @[Mux.scala 31:69:@1850.4]
  assign _T_19873 = valid_5_23 ? 6'h17 : _T_19872; // @[Mux.scala 31:69:@1851.4]
  assign _T_19874 = valid_5_22 ? 6'h16 : _T_19873; // @[Mux.scala 31:69:@1852.4]
  assign _T_19875 = valid_5_21 ? 6'h15 : _T_19874; // @[Mux.scala 31:69:@1853.4]
  assign _T_19876 = valid_5_20 ? 6'h14 : _T_19875; // @[Mux.scala 31:69:@1854.4]
  assign _T_19877 = valid_5_19 ? 6'h13 : _T_19876; // @[Mux.scala 31:69:@1855.4]
  assign _T_19878 = valid_5_18 ? 6'h12 : _T_19877; // @[Mux.scala 31:69:@1856.4]
  assign _T_19879 = valid_5_17 ? 6'h11 : _T_19878; // @[Mux.scala 31:69:@1857.4]
  assign _T_19880 = valid_5_16 ? 6'h10 : _T_19879; // @[Mux.scala 31:69:@1858.4]
  assign _T_19881 = valid_5_15 ? 6'hf : _T_19880; // @[Mux.scala 31:69:@1859.4]
  assign _T_19882 = valid_5_14 ? 6'he : _T_19881; // @[Mux.scala 31:69:@1860.4]
  assign _T_19883 = valid_5_13 ? 6'hd : _T_19882; // @[Mux.scala 31:69:@1861.4]
  assign _T_19884 = valid_5_12 ? 6'hc : _T_19883; // @[Mux.scala 31:69:@1862.4]
  assign _T_19885 = valid_5_11 ? 6'hb : _T_19884; // @[Mux.scala 31:69:@1863.4]
  assign _T_19886 = valid_5_10 ? 6'ha : _T_19885; // @[Mux.scala 31:69:@1864.4]
  assign _T_19887 = valid_5_9 ? 6'h9 : _T_19886; // @[Mux.scala 31:69:@1865.4]
  assign _T_19888 = valid_5_8 ? 6'h8 : _T_19887; // @[Mux.scala 31:69:@1866.4]
  assign _T_19889 = valid_5_7 ? 6'h7 : _T_19888; // @[Mux.scala 31:69:@1867.4]
  assign _T_19890 = valid_5_6 ? 6'h6 : _T_19889; // @[Mux.scala 31:69:@1868.4]
  assign _T_19891 = valid_5_5 ? 6'h5 : _T_19890; // @[Mux.scala 31:69:@1869.4]
  assign _T_19892 = valid_5_4 ? 6'h4 : _T_19891; // @[Mux.scala 31:69:@1870.4]
  assign _T_19893 = valid_5_3 ? 6'h3 : _T_19892; // @[Mux.scala 31:69:@1871.4]
  assign _T_19894 = valid_5_2 ? 6'h2 : _T_19893; // @[Mux.scala 31:69:@1872.4]
  assign _T_19895 = valid_5_1 ? 6'h1 : _T_19894; // @[Mux.scala 31:69:@1873.4]
  assign select_5 = valid_5_0 ? 6'h0 : _T_19895; // @[Mux.scala 31:69:@1874.4]
  assign _GEN_321 = 6'h1 == select_5 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_322 = 6'h2 == select_5 ? io_inData_2 : _GEN_321; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_323 = 6'h3 == select_5 ? io_inData_3 : _GEN_322; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_324 = 6'h4 == select_5 ? io_inData_4 : _GEN_323; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_325 = 6'h5 == select_5 ? io_inData_5 : _GEN_324; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_326 = 6'h6 == select_5 ? io_inData_6 : _GEN_325; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_327 = 6'h7 == select_5 ? io_inData_7 : _GEN_326; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_328 = 6'h8 == select_5 ? io_inData_8 : _GEN_327; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_329 = 6'h9 == select_5 ? io_inData_9 : _GEN_328; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_330 = 6'ha == select_5 ? io_inData_10 : _GEN_329; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_331 = 6'hb == select_5 ? io_inData_11 : _GEN_330; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_332 = 6'hc == select_5 ? io_inData_12 : _GEN_331; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_333 = 6'hd == select_5 ? io_inData_13 : _GEN_332; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_334 = 6'he == select_5 ? io_inData_14 : _GEN_333; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_335 = 6'hf == select_5 ? io_inData_15 : _GEN_334; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_336 = 6'h10 == select_5 ? io_inData_16 : _GEN_335; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_337 = 6'h11 == select_5 ? io_inData_17 : _GEN_336; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_338 = 6'h12 == select_5 ? io_inData_18 : _GEN_337; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_339 = 6'h13 == select_5 ? io_inData_19 : _GEN_338; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_340 = 6'h14 == select_5 ? io_inData_20 : _GEN_339; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_341 = 6'h15 == select_5 ? io_inData_21 : _GEN_340; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_342 = 6'h16 == select_5 ? io_inData_22 : _GEN_341; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_343 = 6'h17 == select_5 ? io_inData_23 : _GEN_342; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_344 = 6'h18 == select_5 ? io_inData_24 : _GEN_343; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_345 = 6'h19 == select_5 ? io_inData_25 : _GEN_344; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_346 = 6'h1a == select_5 ? io_inData_26 : _GEN_345; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_347 = 6'h1b == select_5 ? io_inData_27 : _GEN_346; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_348 = 6'h1c == select_5 ? io_inData_28 : _GEN_347; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_349 = 6'h1d == select_5 ? io_inData_29 : _GEN_348; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_350 = 6'h1e == select_5 ? io_inData_30 : _GEN_349; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_351 = 6'h1f == select_5 ? io_inData_31 : _GEN_350; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_352 = 6'h20 == select_5 ? io_inData_32 : _GEN_351; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_353 = 6'h21 == select_5 ? io_inData_33 : _GEN_352; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_354 = 6'h22 == select_5 ? io_inData_34 : _GEN_353; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_355 = 6'h23 == select_5 ? io_inData_35 : _GEN_354; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_356 = 6'h24 == select_5 ? io_inData_36 : _GEN_355; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_357 = 6'h25 == select_5 ? io_inData_37 : _GEN_356; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_358 = 6'h26 == select_5 ? io_inData_38 : _GEN_357; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_359 = 6'h27 == select_5 ? io_inData_39 : _GEN_358; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_360 = 6'h28 == select_5 ? io_inData_40 : _GEN_359; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_361 = 6'h29 == select_5 ? io_inData_41 : _GEN_360; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_362 = 6'h2a == select_5 ? io_inData_42 : _GEN_361; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_363 = 6'h2b == select_5 ? io_inData_43 : _GEN_362; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_364 = 6'h2c == select_5 ? io_inData_44 : _GEN_363; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_365 = 6'h2d == select_5 ? io_inData_45 : _GEN_364; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_366 = 6'h2e == select_5 ? io_inData_46 : _GEN_365; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_367 = 6'h2f == select_5 ? io_inData_47 : _GEN_366; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_368 = 6'h30 == select_5 ? io_inData_48 : _GEN_367; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_369 = 6'h31 == select_5 ? io_inData_49 : _GEN_368; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_370 = 6'h32 == select_5 ? io_inData_50 : _GEN_369; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_371 = 6'h33 == select_5 ? io_inData_51 : _GEN_370; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_372 = 6'h34 == select_5 ? io_inData_52 : _GEN_371; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_373 = 6'h35 == select_5 ? io_inData_53 : _GEN_372; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_374 = 6'h36 == select_5 ? io_inData_54 : _GEN_373; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_375 = 6'h37 == select_5 ? io_inData_55 : _GEN_374; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_376 = 6'h38 == select_5 ? io_inData_56 : _GEN_375; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_377 = 6'h39 == select_5 ? io_inData_57 : _GEN_376; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_378 = 6'h3a == select_5 ? io_inData_58 : _GEN_377; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_379 = 6'h3b == select_5 ? io_inData_59 : _GEN_378; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_380 = 6'h3c == select_5 ? io_inData_60 : _GEN_379; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_381 = 6'h3d == select_5 ? io_inData_61 : _GEN_380; // @[Switch.scala 33:19:@1876.4]
  assign _GEN_382 = 6'h3e == select_5 ? io_inData_62 : _GEN_381; // @[Switch.scala 33:19:@1876.4]
  assign _T_19904 = {valid_5_7,valid_5_6,valid_5_5,valid_5_4,valid_5_3,valid_5_2,valid_5_1,valid_5_0}; // @[Switch.scala 34:32:@1883.4]
  assign _T_19912 = {valid_5_15,valid_5_14,valid_5_13,valid_5_12,valid_5_11,valid_5_10,valid_5_9,valid_5_8,_T_19904}; // @[Switch.scala 34:32:@1891.4]
  assign _T_19919 = {valid_5_23,valid_5_22,valid_5_21,valid_5_20,valid_5_19,valid_5_18,valid_5_17,valid_5_16}; // @[Switch.scala 34:32:@1898.4]
  assign _T_19928 = {valid_5_31,valid_5_30,valid_5_29,valid_5_28,valid_5_27,valid_5_26,valid_5_25,valid_5_24,_T_19919,_T_19912}; // @[Switch.scala 34:32:@1907.4]
  assign _T_19935 = {valid_5_39,valid_5_38,valid_5_37,valid_5_36,valid_5_35,valid_5_34,valid_5_33,valid_5_32}; // @[Switch.scala 34:32:@1914.4]
  assign _T_19943 = {valid_5_47,valid_5_46,valid_5_45,valid_5_44,valid_5_43,valid_5_42,valid_5_41,valid_5_40,_T_19935}; // @[Switch.scala 34:32:@1922.4]
  assign _T_19950 = {valid_5_55,valid_5_54,valid_5_53,valid_5_52,valid_5_51,valid_5_50,valid_5_49,valid_5_48}; // @[Switch.scala 34:32:@1929.4]
  assign _T_19959 = {valid_5_63,valid_5_62,valid_5_61,valid_5_60,valid_5_59,valid_5_58,valid_5_57,valid_5_56,_T_19950,_T_19943}; // @[Switch.scala 34:32:@1938.4]
  assign _T_19960 = {_T_19959,_T_19928}; // @[Switch.scala 34:32:@1939.4]
  assign _T_19964 = io_inAddr_0 == 6'h6; // @[Switch.scala 30:53:@1942.4]
  assign valid_6_0 = io_inValid_0 & _T_19964; // @[Switch.scala 30:36:@1943.4]
  assign _T_19967 = io_inAddr_1 == 6'h6; // @[Switch.scala 30:53:@1945.4]
  assign valid_6_1 = io_inValid_1 & _T_19967; // @[Switch.scala 30:36:@1946.4]
  assign _T_19970 = io_inAddr_2 == 6'h6; // @[Switch.scala 30:53:@1948.4]
  assign valid_6_2 = io_inValid_2 & _T_19970; // @[Switch.scala 30:36:@1949.4]
  assign _T_19973 = io_inAddr_3 == 6'h6; // @[Switch.scala 30:53:@1951.4]
  assign valid_6_3 = io_inValid_3 & _T_19973; // @[Switch.scala 30:36:@1952.4]
  assign _T_19976 = io_inAddr_4 == 6'h6; // @[Switch.scala 30:53:@1954.4]
  assign valid_6_4 = io_inValid_4 & _T_19976; // @[Switch.scala 30:36:@1955.4]
  assign _T_19979 = io_inAddr_5 == 6'h6; // @[Switch.scala 30:53:@1957.4]
  assign valid_6_5 = io_inValid_5 & _T_19979; // @[Switch.scala 30:36:@1958.4]
  assign _T_19982 = io_inAddr_6 == 6'h6; // @[Switch.scala 30:53:@1960.4]
  assign valid_6_6 = io_inValid_6 & _T_19982; // @[Switch.scala 30:36:@1961.4]
  assign _T_19985 = io_inAddr_7 == 6'h6; // @[Switch.scala 30:53:@1963.4]
  assign valid_6_7 = io_inValid_7 & _T_19985; // @[Switch.scala 30:36:@1964.4]
  assign _T_19988 = io_inAddr_8 == 6'h6; // @[Switch.scala 30:53:@1966.4]
  assign valid_6_8 = io_inValid_8 & _T_19988; // @[Switch.scala 30:36:@1967.4]
  assign _T_19991 = io_inAddr_9 == 6'h6; // @[Switch.scala 30:53:@1969.4]
  assign valid_6_9 = io_inValid_9 & _T_19991; // @[Switch.scala 30:36:@1970.4]
  assign _T_19994 = io_inAddr_10 == 6'h6; // @[Switch.scala 30:53:@1972.4]
  assign valid_6_10 = io_inValid_10 & _T_19994; // @[Switch.scala 30:36:@1973.4]
  assign _T_19997 = io_inAddr_11 == 6'h6; // @[Switch.scala 30:53:@1975.4]
  assign valid_6_11 = io_inValid_11 & _T_19997; // @[Switch.scala 30:36:@1976.4]
  assign _T_20000 = io_inAddr_12 == 6'h6; // @[Switch.scala 30:53:@1978.4]
  assign valid_6_12 = io_inValid_12 & _T_20000; // @[Switch.scala 30:36:@1979.4]
  assign _T_20003 = io_inAddr_13 == 6'h6; // @[Switch.scala 30:53:@1981.4]
  assign valid_6_13 = io_inValid_13 & _T_20003; // @[Switch.scala 30:36:@1982.4]
  assign _T_20006 = io_inAddr_14 == 6'h6; // @[Switch.scala 30:53:@1984.4]
  assign valid_6_14 = io_inValid_14 & _T_20006; // @[Switch.scala 30:36:@1985.4]
  assign _T_20009 = io_inAddr_15 == 6'h6; // @[Switch.scala 30:53:@1987.4]
  assign valid_6_15 = io_inValid_15 & _T_20009; // @[Switch.scala 30:36:@1988.4]
  assign _T_20012 = io_inAddr_16 == 6'h6; // @[Switch.scala 30:53:@1990.4]
  assign valid_6_16 = io_inValid_16 & _T_20012; // @[Switch.scala 30:36:@1991.4]
  assign _T_20015 = io_inAddr_17 == 6'h6; // @[Switch.scala 30:53:@1993.4]
  assign valid_6_17 = io_inValid_17 & _T_20015; // @[Switch.scala 30:36:@1994.4]
  assign _T_20018 = io_inAddr_18 == 6'h6; // @[Switch.scala 30:53:@1996.4]
  assign valid_6_18 = io_inValid_18 & _T_20018; // @[Switch.scala 30:36:@1997.4]
  assign _T_20021 = io_inAddr_19 == 6'h6; // @[Switch.scala 30:53:@1999.4]
  assign valid_6_19 = io_inValid_19 & _T_20021; // @[Switch.scala 30:36:@2000.4]
  assign _T_20024 = io_inAddr_20 == 6'h6; // @[Switch.scala 30:53:@2002.4]
  assign valid_6_20 = io_inValid_20 & _T_20024; // @[Switch.scala 30:36:@2003.4]
  assign _T_20027 = io_inAddr_21 == 6'h6; // @[Switch.scala 30:53:@2005.4]
  assign valid_6_21 = io_inValid_21 & _T_20027; // @[Switch.scala 30:36:@2006.4]
  assign _T_20030 = io_inAddr_22 == 6'h6; // @[Switch.scala 30:53:@2008.4]
  assign valid_6_22 = io_inValid_22 & _T_20030; // @[Switch.scala 30:36:@2009.4]
  assign _T_20033 = io_inAddr_23 == 6'h6; // @[Switch.scala 30:53:@2011.4]
  assign valid_6_23 = io_inValid_23 & _T_20033; // @[Switch.scala 30:36:@2012.4]
  assign _T_20036 = io_inAddr_24 == 6'h6; // @[Switch.scala 30:53:@2014.4]
  assign valid_6_24 = io_inValid_24 & _T_20036; // @[Switch.scala 30:36:@2015.4]
  assign _T_20039 = io_inAddr_25 == 6'h6; // @[Switch.scala 30:53:@2017.4]
  assign valid_6_25 = io_inValid_25 & _T_20039; // @[Switch.scala 30:36:@2018.4]
  assign _T_20042 = io_inAddr_26 == 6'h6; // @[Switch.scala 30:53:@2020.4]
  assign valid_6_26 = io_inValid_26 & _T_20042; // @[Switch.scala 30:36:@2021.4]
  assign _T_20045 = io_inAddr_27 == 6'h6; // @[Switch.scala 30:53:@2023.4]
  assign valid_6_27 = io_inValid_27 & _T_20045; // @[Switch.scala 30:36:@2024.4]
  assign _T_20048 = io_inAddr_28 == 6'h6; // @[Switch.scala 30:53:@2026.4]
  assign valid_6_28 = io_inValid_28 & _T_20048; // @[Switch.scala 30:36:@2027.4]
  assign _T_20051 = io_inAddr_29 == 6'h6; // @[Switch.scala 30:53:@2029.4]
  assign valid_6_29 = io_inValid_29 & _T_20051; // @[Switch.scala 30:36:@2030.4]
  assign _T_20054 = io_inAddr_30 == 6'h6; // @[Switch.scala 30:53:@2032.4]
  assign valid_6_30 = io_inValid_30 & _T_20054; // @[Switch.scala 30:36:@2033.4]
  assign _T_20057 = io_inAddr_31 == 6'h6; // @[Switch.scala 30:53:@2035.4]
  assign valid_6_31 = io_inValid_31 & _T_20057; // @[Switch.scala 30:36:@2036.4]
  assign _T_20060 = io_inAddr_32 == 6'h6; // @[Switch.scala 30:53:@2038.4]
  assign valid_6_32 = io_inValid_32 & _T_20060; // @[Switch.scala 30:36:@2039.4]
  assign _T_20063 = io_inAddr_33 == 6'h6; // @[Switch.scala 30:53:@2041.4]
  assign valid_6_33 = io_inValid_33 & _T_20063; // @[Switch.scala 30:36:@2042.4]
  assign _T_20066 = io_inAddr_34 == 6'h6; // @[Switch.scala 30:53:@2044.4]
  assign valid_6_34 = io_inValid_34 & _T_20066; // @[Switch.scala 30:36:@2045.4]
  assign _T_20069 = io_inAddr_35 == 6'h6; // @[Switch.scala 30:53:@2047.4]
  assign valid_6_35 = io_inValid_35 & _T_20069; // @[Switch.scala 30:36:@2048.4]
  assign _T_20072 = io_inAddr_36 == 6'h6; // @[Switch.scala 30:53:@2050.4]
  assign valid_6_36 = io_inValid_36 & _T_20072; // @[Switch.scala 30:36:@2051.4]
  assign _T_20075 = io_inAddr_37 == 6'h6; // @[Switch.scala 30:53:@2053.4]
  assign valid_6_37 = io_inValid_37 & _T_20075; // @[Switch.scala 30:36:@2054.4]
  assign _T_20078 = io_inAddr_38 == 6'h6; // @[Switch.scala 30:53:@2056.4]
  assign valid_6_38 = io_inValid_38 & _T_20078; // @[Switch.scala 30:36:@2057.4]
  assign _T_20081 = io_inAddr_39 == 6'h6; // @[Switch.scala 30:53:@2059.4]
  assign valid_6_39 = io_inValid_39 & _T_20081; // @[Switch.scala 30:36:@2060.4]
  assign _T_20084 = io_inAddr_40 == 6'h6; // @[Switch.scala 30:53:@2062.4]
  assign valid_6_40 = io_inValid_40 & _T_20084; // @[Switch.scala 30:36:@2063.4]
  assign _T_20087 = io_inAddr_41 == 6'h6; // @[Switch.scala 30:53:@2065.4]
  assign valid_6_41 = io_inValid_41 & _T_20087; // @[Switch.scala 30:36:@2066.4]
  assign _T_20090 = io_inAddr_42 == 6'h6; // @[Switch.scala 30:53:@2068.4]
  assign valid_6_42 = io_inValid_42 & _T_20090; // @[Switch.scala 30:36:@2069.4]
  assign _T_20093 = io_inAddr_43 == 6'h6; // @[Switch.scala 30:53:@2071.4]
  assign valid_6_43 = io_inValid_43 & _T_20093; // @[Switch.scala 30:36:@2072.4]
  assign _T_20096 = io_inAddr_44 == 6'h6; // @[Switch.scala 30:53:@2074.4]
  assign valid_6_44 = io_inValid_44 & _T_20096; // @[Switch.scala 30:36:@2075.4]
  assign _T_20099 = io_inAddr_45 == 6'h6; // @[Switch.scala 30:53:@2077.4]
  assign valid_6_45 = io_inValid_45 & _T_20099; // @[Switch.scala 30:36:@2078.4]
  assign _T_20102 = io_inAddr_46 == 6'h6; // @[Switch.scala 30:53:@2080.4]
  assign valid_6_46 = io_inValid_46 & _T_20102; // @[Switch.scala 30:36:@2081.4]
  assign _T_20105 = io_inAddr_47 == 6'h6; // @[Switch.scala 30:53:@2083.4]
  assign valid_6_47 = io_inValid_47 & _T_20105; // @[Switch.scala 30:36:@2084.4]
  assign _T_20108 = io_inAddr_48 == 6'h6; // @[Switch.scala 30:53:@2086.4]
  assign valid_6_48 = io_inValid_48 & _T_20108; // @[Switch.scala 30:36:@2087.4]
  assign _T_20111 = io_inAddr_49 == 6'h6; // @[Switch.scala 30:53:@2089.4]
  assign valid_6_49 = io_inValid_49 & _T_20111; // @[Switch.scala 30:36:@2090.4]
  assign _T_20114 = io_inAddr_50 == 6'h6; // @[Switch.scala 30:53:@2092.4]
  assign valid_6_50 = io_inValid_50 & _T_20114; // @[Switch.scala 30:36:@2093.4]
  assign _T_20117 = io_inAddr_51 == 6'h6; // @[Switch.scala 30:53:@2095.4]
  assign valid_6_51 = io_inValid_51 & _T_20117; // @[Switch.scala 30:36:@2096.4]
  assign _T_20120 = io_inAddr_52 == 6'h6; // @[Switch.scala 30:53:@2098.4]
  assign valid_6_52 = io_inValid_52 & _T_20120; // @[Switch.scala 30:36:@2099.4]
  assign _T_20123 = io_inAddr_53 == 6'h6; // @[Switch.scala 30:53:@2101.4]
  assign valid_6_53 = io_inValid_53 & _T_20123; // @[Switch.scala 30:36:@2102.4]
  assign _T_20126 = io_inAddr_54 == 6'h6; // @[Switch.scala 30:53:@2104.4]
  assign valid_6_54 = io_inValid_54 & _T_20126; // @[Switch.scala 30:36:@2105.4]
  assign _T_20129 = io_inAddr_55 == 6'h6; // @[Switch.scala 30:53:@2107.4]
  assign valid_6_55 = io_inValid_55 & _T_20129; // @[Switch.scala 30:36:@2108.4]
  assign _T_20132 = io_inAddr_56 == 6'h6; // @[Switch.scala 30:53:@2110.4]
  assign valid_6_56 = io_inValid_56 & _T_20132; // @[Switch.scala 30:36:@2111.4]
  assign _T_20135 = io_inAddr_57 == 6'h6; // @[Switch.scala 30:53:@2113.4]
  assign valid_6_57 = io_inValid_57 & _T_20135; // @[Switch.scala 30:36:@2114.4]
  assign _T_20138 = io_inAddr_58 == 6'h6; // @[Switch.scala 30:53:@2116.4]
  assign valid_6_58 = io_inValid_58 & _T_20138; // @[Switch.scala 30:36:@2117.4]
  assign _T_20141 = io_inAddr_59 == 6'h6; // @[Switch.scala 30:53:@2119.4]
  assign valid_6_59 = io_inValid_59 & _T_20141; // @[Switch.scala 30:36:@2120.4]
  assign _T_20144 = io_inAddr_60 == 6'h6; // @[Switch.scala 30:53:@2122.4]
  assign valid_6_60 = io_inValid_60 & _T_20144; // @[Switch.scala 30:36:@2123.4]
  assign _T_20147 = io_inAddr_61 == 6'h6; // @[Switch.scala 30:53:@2125.4]
  assign valid_6_61 = io_inValid_61 & _T_20147; // @[Switch.scala 30:36:@2126.4]
  assign _T_20150 = io_inAddr_62 == 6'h6; // @[Switch.scala 30:53:@2128.4]
  assign valid_6_62 = io_inValid_62 & _T_20150; // @[Switch.scala 30:36:@2129.4]
  assign _T_20153 = io_inAddr_63 == 6'h6; // @[Switch.scala 30:53:@2131.4]
  assign valid_6_63 = io_inValid_63 & _T_20153; // @[Switch.scala 30:36:@2132.4]
  assign _T_20219 = valid_6_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@2134.4]
  assign _T_20220 = valid_6_61 ? 6'h3d : _T_20219; // @[Mux.scala 31:69:@2135.4]
  assign _T_20221 = valid_6_60 ? 6'h3c : _T_20220; // @[Mux.scala 31:69:@2136.4]
  assign _T_20222 = valid_6_59 ? 6'h3b : _T_20221; // @[Mux.scala 31:69:@2137.4]
  assign _T_20223 = valid_6_58 ? 6'h3a : _T_20222; // @[Mux.scala 31:69:@2138.4]
  assign _T_20224 = valid_6_57 ? 6'h39 : _T_20223; // @[Mux.scala 31:69:@2139.4]
  assign _T_20225 = valid_6_56 ? 6'h38 : _T_20224; // @[Mux.scala 31:69:@2140.4]
  assign _T_20226 = valid_6_55 ? 6'h37 : _T_20225; // @[Mux.scala 31:69:@2141.4]
  assign _T_20227 = valid_6_54 ? 6'h36 : _T_20226; // @[Mux.scala 31:69:@2142.4]
  assign _T_20228 = valid_6_53 ? 6'h35 : _T_20227; // @[Mux.scala 31:69:@2143.4]
  assign _T_20229 = valid_6_52 ? 6'h34 : _T_20228; // @[Mux.scala 31:69:@2144.4]
  assign _T_20230 = valid_6_51 ? 6'h33 : _T_20229; // @[Mux.scala 31:69:@2145.4]
  assign _T_20231 = valid_6_50 ? 6'h32 : _T_20230; // @[Mux.scala 31:69:@2146.4]
  assign _T_20232 = valid_6_49 ? 6'h31 : _T_20231; // @[Mux.scala 31:69:@2147.4]
  assign _T_20233 = valid_6_48 ? 6'h30 : _T_20232; // @[Mux.scala 31:69:@2148.4]
  assign _T_20234 = valid_6_47 ? 6'h2f : _T_20233; // @[Mux.scala 31:69:@2149.4]
  assign _T_20235 = valid_6_46 ? 6'h2e : _T_20234; // @[Mux.scala 31:69:@2150.4]
  assign _T_20236 = valid_6_45 ? 6'h2d : _T_20235; // @[Mux.scala 31:69:@2151.4]
  assign _T_20237 = valid_6_44 ? 6'h2c : _T_20236; // @[Mux.scala 31:69:@2152.4]
  assign _T_20238 = valid_6_43 ? 6'h2b : _T_20237; // @[Mux.scala 31:69:@2153.4]
  assign _T_20239 = valid_6_42 ? 6'h2a : _T_20238; // @[Mux.scala 31:69:@2154.4]
  assign _T_20240 = valid_6_41 ? 6'h29 : _T_20239; // @[Mux.scala 31:69:@2155.4]
  assign _T_20241 = valid_6_40 ? 6'h28 : _T_20240; // @[Mux.scala 31:69:@2156.4]
  assign _T_20242 = valid_6_39 ? 6'h27 : _T_20241; // @[Mux.scala 31:69:@2157.4]
  assign _T_20243 = valid_6_38 ? 6'h26 : _T_20242; // @[Mux.scala 31:69:@2158.4]
  assign _T_20244 = valid_6_37 ? 6'h25 : _T_20243; // @[Mux.scala 31:69:@2159.4]
  assign _T_20245 = valid_6_36 ? 6'h24 : _T_20244; // @[Mux.scala 31:69:@2160.4]
  assign _T_20246 = valid_6_35 ? 6'h23 : _T_20245; // @[Mux.scala 31:69:@2161.4]
  assign _T_20247 = valid_6_34 ? 6'h22 : _T_20246; // @[Mux.scala 31:69:@2162.4]
  assign _T_20248 = valid_6_33 ? 6'h21 : _T_20247; // @[Mux.scala 31:69:@2163.4]
  assign _T_20249 = valid_6_32 ? 6'h20 : _T_20248; // @[Mux.scala 31:69:@2164.4]
  assign _T_20250 = valid_6_31 ? 6'h1f : _T_20249; // @[Mux.scala 31:69:@2165.4]
  assign _T_20251 = valid_6_30 ? 6'h1e : _T_20250; // @[Mux.scala 31:69:@2166.4]
  assign _T_20252 = valid_6_29 ? 6'h1d : _T_20251; // @[Mux.scala 31:69:@2167.4]
  assign _T_20253 = valid_6_28 ? 6'h1c : _T_20252; // @[Mux.scala 31:69:@2168.4]
  assign _T_20254 = valid_6_27 ? 6'h1b : _T_20253; // @[Mux.scala 31:69:@2169.4]
  assign _T_20255 = valid_6_26 ? 6'h1a : _T_20254; // @[Mux.scala 31:69:@2170.4]
  assign _T_20256 = valid_6_25 ? 6'h19 : _T_20255; // @[Mux.scala 31:69:@2171.4]
  assign _T_20257 = valid_6_24 ? 6'h18 : _T_20256; // @[Mux.scala 31:69:@2172.4]
  assign _T_20258 = valid_6_23 ? 6'h17 : _T_20257; // @[Mux.scala 31:69:@2173.4]
  assign _T_20259 = valid_6_22 ? 6'h16 : _T_20258; // @[Mux.scala 31:69:@2174.4]
  assign _T_20260 = valid_6_21 ? 6'h15 : _T_20259; // @[Mux.scala 31:69:@2175.4]
  assign _T_20261 = valid_6_20 ? 6'h14 : _T_20260; // @[Mux.scala 31:69:@2176.4]
  assign _T_20262 = valid_6_19 ? 6'h13 : _T_20261; // @[Mux.scala 31:69:@2177.4]
  assign _T_20263 = valid_6_18 ? 6'h12 : _T_20262; // @[Mux.scala 31:69:@2178.4]
  assign _T_20264 = valid_6_17 ? 6'h11 : _T_20263; // @[Mux.scala 31:69:@2179.4]
  assign _T_20265 = valid_6_16 ? 6'h10 : _T_20264; // @[Mux.scala 31:69:@2180.4]
  assign _T_20266 = valid_6_15 ? 6'hf : _T_20265; // @[Mux.scala 31:69:@2181.4]
  assign _T_20267 = valid_6_14 ? 6'he : _T_20266; // @[Mux.scala 31:69:@2182.4]
  assign _T_20268 = valid_6_13 ? 6'hd : _T_20267; // @[Mux.scala 31:69:@2183.4]
  assign _T_20269 = valid_6_12 ? 6'hc : _T_20268; // @[Mux.scala 31:69:@2184.4]
  assign _T_20270 = valid_6_11 ? 6'hb : _T_20269; // @[Mux.scala 31:69:@2185.4]
  assign _T_20271 = valid_6_10 ? 6'ha : _T_20270; // @[Mux.scala 31:69:@2186.4]
  assign _T_20272 = valid_6_9 ? 6'h9 : _T_20271; // @[Mux.scala 31:69:@2187.4]
  assign _T_20273 = valid_6_8 ? 6'h8 : _T_20272; // @[Mux.scala 31:69:@2188.4]
  assign _T_20274 = valid_6_7 ? 6'h7 : _T_20273; // @[Mux.scala 31:69:@2189.4]
  assign _T_20275 = valid_6_6 ? 6'h6 : _T_20274; // @[Mux.scala 31:69:@2190.4]
  assign _T_20276 = valid_6_5 ? 6'h5 : _T_20275; // @[Mux.scala 31:69:@2191.4]
  assign _T_20277 = valid_6_4 ? 6'h4 : _T_20276; // @[Mux.scala 31:69:@2192.4]
  assign _T_20278 = valid_6_3 ? 6'h3 : _T_20277; // @[Mux.scala 31:69:@2193.4]
  assign _T_20279 = valid_6_2 ? 6'h2 : _T_20278; // @[Mux.scala 31:69:@2194.4]
  assign _T_20280 = valid_6_1 ? 6'h1 : _T_20279; // @[Mux.scala 31:69:@2195.4]
  assign select_6 = valid_6_0 ? 6'h0 : _T_20280; // @[Mux.scala 31:69:@2196.4]
  assign _GEN_385 = 6'h1 == select_6 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_386 = 6'h2 == select_6 ? io_inData_2 : _GEN_385; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_387 = 6'h3 == select_6 ? io_inData_3 : _GEN_386; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_388 = 6'h4 == select_6 ? io_inData_4 : _GEN_387; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_389 = 6'h5 == select_6 ? io_inData_5 : _GEN_388; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_390 = 6'h6 == select_6 ? io_inData_6 : _GEN_389; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_391 = 6'h7 == select_6 ? io_inData_7 : _GEN_390; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_392 = 6'h8 == select_6 ? io_inData_8 : _GEN_391; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_393 = 6'h9 == select_6 ? io_inData_9 : _GEN_392; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_394 = 6'ha == select_6 ? io_inData_10 : _GEN_393; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_395 = 6'hb == select_6 ? io_inData_11 : _GEN_394; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_396 = 6'hc == select_6 ? io_inData_12 : _GEN_395; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_397 = 6'hd == select_6 ? io_inData_13 : _GEN_396; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_398 = 6'he == select_6 ? io_inData_14 : _GEN_397; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_399 = 6'hf == select_6 ? io_inData_15 : _GEN_398; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_400 = 6'h10 == select_6 ? io_inData_16 : _GEN_399; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_401 = 6'h11 == select_6 ? io_inData_17 : _GEN_400; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_402 = 6'h12 == select_6 ? io_inData_18 : _GEN_401; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_403 = 6'h13 == select_6 ? io_inData_19 : _GEN_402; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_404 = 6'h14 == select_6 ? io_inData_20 : _GEN_403; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_405 = 6'h15 == select_6 ? io_inData_21 : _GEN_404; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_406 = 6'h16 == select_6 ? io_inData_22 : _GEN_405; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_407 = 6'h17 == select_6 ? io_inData_23 : _GEN_406; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_408 = 6'h18 == select_6 ? io_inData_24 : _GEN_407; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_409 = 6'h19 == select_6 ? io_inData_25 : _GEN_408; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_410 = 6'h1a == select_6 ? io_inData_26 : _GEN_409; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_411 = 6'h1b == select_6 ? io_inData_27 : _GEN_410; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_412 = 6'h1c == select_6 ? io_inData_28 : _GEN_411; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_413 = 6'h1d == select_6 ? io_inData_29 : _GEN_412; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_414 = 6'h1e == select_6 ? io_inData_30 : _GEN_413; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_415 = 6'h1f == select_6 ? io_inData_31 : _GEN_414; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_416 = 6'h20 == select_6 ? io_inData_32 : _GEN_415; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_417 = 6'h21 == select_6 ? io_inData_33 : _GEN_416; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_418 = 6'h22 == select_6 ? io_inData_34 : _GEN_417; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_419 = 6'h23 == select_6 ? io_inData_35 : _GEN_418; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_420 = 6'h24 == select_6 ? io_inData_36 : _GEN_419; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_421 = 6'h25 == select_6 ? io_inData_37 : _GEN_420; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_422 = 6'h26 == select_6 ? io_inData_38 : _GEN_421; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_423 = 6'h27 == select_6 ? io_inData_39 : _GEN_422; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_424 = 6'h28 == select_6 ? io_inData_40 : _GEN_423; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_425 = 6'h29 == select_6 ? io_inData_41 : _GEN_424; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_426 = 6'h2a == select_6 ? io_inData_42 : _GEN_425; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_427 = 6'h2b == select_6 ? io_inData_43 : _GEN_426; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_428 = 6'h2c == select_6 ? io_inData_44 : _GEN_427; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_429 = 6'h2d == select_6 ? io_inData_45 : _GEN_428; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_430 = 6'h2e == select_6 ? io_inData_46 : _GEN_429; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_431 = 6'h2f == select_6 ? io_inData_47 : _GEN_430; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_432 = 6'h30 == select_6 ? io_inData_48 : _GEN_431; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_433 = 6'h31 == select_6 ? io_inData_49 : _GEN_432; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_434 = 6'h32 == select_6 ? io_inData_50 : _GEN_433; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_435 = 6'h33 == select_6 ? io_inData_51 : _GEN_434; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_436 = 6'h34 == select_6 ? io_inData_52 : _GEN_435; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_437 = 6'h35 == select_6 ? io_inData_53 : _GEN_436; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_438 = 6'h36 == select_6 ? io_inData_54 : _GEN_437; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_439 = 6'h37 == select_6 ? io_inData_55 : _GEN_438; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_440 = 6'h38 == select_6 ? io_inData_56 : _GEN_439; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_441 = 6'h39 == select_6 ? io_inData_57 : _GEN_440; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_442 = 6'h3a == select_6 ? io_inData_58 : _GEN_441; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_443 = 6'h3b == select_6 ? io_inData_59 : _GEN_442; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_444 = 6'h3c == select_6 ? io_inData_60 : _GEN_443; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_445 = 6'h3d == select_6 ? io_inData_61 : _GEN_444; // @[Switch.scala 33:19:@2198.4]
  assign _GEN_446 = 6'h3e == select_6 ? io_inData_62 : _GEN_445; // @[Switch.scala 33:19:@2198.4]
  assign _T_20289 = {valid_6_7,valid_6_6,valid_6_5,valid_6_4,valid_6_3,valid_6_2,valid_6_1,valid_6_0}; // @[Switch.scala 34:32:@2205.4]
  assign _T_20297 = {valid_6_15,valid_6_14,valid_6_13,valid_6_12,valid_6_11,valid_6_10,valid_6_9,valid_6_8,_T_20289}; // @[Switch.scala 34:32:@2213.4]
  assign _T_20304 = {valid_6_23,valid_6_22,valid_6_21,valid_6_20,valid_6_19,valid_6_18,valid_6_17,valid_6_16}; // @[Switch.scala 34:32:@2220.4]
  assign _T_20313 = {valid_6_31,valid_6_30,valid_6_29,valid_6_28,valid_6_27,valid_6_26,valid_6_25,valid_6_24,_T_20304,_T_20297}; // @[Switch.scala 34:32:@2229.4]
  assign _T_20320 = {valid_6_39,valid_6_38,valid_6_37,valid_6_36,valid_6_35,valid_6_34,valid_6_33,valid_6_32}; // @[Switch.scala 34:32:@2236.4]
  assign _T_20328 = {valid_6_47,valid_6_46,valid_6_45,valid_6_44,valid_6_43,valid_6_42,valid_6_41,valid_6_40,_T_20320}; // @[Switch.scala 34:32:@2244.4]
  assign _T_20335 = {valid_6_55,valid_6_54,valid_6_53,valid_6_52,valid_6_51,valid_6_50,valid_6_49,valid_6_48}; // @[Switch.scala 34:32:@2251.4]
  assign _T_20344 = {valid_6_63,valid_6_62,valid_6_61,valid_6_60,valid_6_59,valid_6_58,valid_6_57,valid_6_56,_T_20335,_T_20328}; // @[Switch.scala 34:32:@2260.4]
  assign _T_20345 = {_T_20344,_T_20313}; // @[Switch.scala 34:32:@2261.4]
  assign _T_20349 = io_inAddr_0 == 6'h7; // @[Switch.scala 30:53:@2264.4]
  assign valid_7_0 = io_inValid_0 & _T_20349; // @[Switch.scala 30:36:@2265.4]
  assign _T_20352 = io_inAddr_1 == 6'h7; // @[Switch.scala 30:53:@2267.4]
  assign valid_7_1 = io_inValid_1 & _T_20352; // @[Switch.scala 30:36:@2268.4]
  assign _T_20355 = io_inAddr_2 == 6'h7; // @[Switch.scala 30:53:@2270.4]
  assign valid_7_2 = io_inValid_2 & _T_20355; // @[Switch.scala 30:36:@2271.4]
  assign _T_20358 = io_inAddr_3 == 6'h7; // @[Switch.scala 30:53:@2273.4]
  assign valid_7_3 = io_inValid_3 & _T_20358; // @[Switch.scala 30:36:@2274.4]
  assign _T_20361 = io_inAddr_4 == 6'h7; // @[Switch.scala 30:53:@2276.4]
  assign valid_7_4 = io_inValid_4 & _T_20361; // @[Switch.scala 30:36:@2277.4]
  assign _T_20364 = io_inAddr_5 == 6'h7; // @[Switch.scala 30:53:@2279.4]
  assign valid_7_5 = io_inValid_5 & _T_20364; // @[Switch.scala 30:36:@2280.4]
  assign _T_20367 = io_inAddr_6 == 6'h7; // @[Switch.scala 30:53:@2282.4]
  assign valid_7_6 = io_inValid_6 & _T_20367; // @[Switch.scala 30:36:@2283.4]
  assign _T_20370 = io_inAddr_7 == 6'h7; // @[Switch.scala 30:53:@2285.4]
  assign valid_7_7 = io_inValid_7 & _T_20370; // @[Switch.scala 30:36:@2286.4]
  assign _T_20373 = io_inAddr_8 == 6'h7; // @[Switch.scala 30:53:@2288.4]
  assign valid_7_8 = io_inValid_8 & _T_20373; // @[Switch.scala 30:36:@2289.4]
  assign _T_20376 = io_inAddr_9 == 6'h7; // @[Switch.scala 30:53:@2291.4]
  assign valid_7_9 = io_inValid_9 & _T_20376; // @[Switch.scala 30:36:@2292.4]
  assign _T_20379 = io_inAddr_10 == 6'h7; // @[Switch.scala 30:53:@2294.4]
  assign valid_7_10 = io_inValid_10 & _T_20379; // @[Switch.scala 30:36:@2295.4]
  assign _T_20382 = io_inAddr_11 == 6'h7; // @[Switch.scala 30:53:@2297.4]
  assign valid_7_11 = io_inValid_11 & _T_20382; // @[Switch.scala 30:36:@2298.4]
  assign _T_20385 = io_inAddr_12 == 6'h7; // @[Switch.scala 30:53:@2300.4]
  assign valid_7_12 = io_inValid_12 & _T_20385; // @[Switch.scala 30:36:@2301.4]
  assign _T_20388 = io_inAddr_13 == 6'h7; // @[Switch.scala 30:53:@2303.4]
  assign valid_7_13 = io_inValid_13 & _T_20388; // @[Switch.scala 30:36:@2304.4]
  assign _T_20391 = io_inAddr_14 == 6'h7; // @[Switch.scala 30:53:@2306.4]
  assign valid_7_14 = io_inValid_14 & _T_20391; // @[Switch.scala 30:36:@2307.4]
  assign _T_20394 = io_inAddr_15 == 6'h7; // @[Switch.scala 30:53:@2309.4]
  assign valid_7_15 = io_inValid_15 & _T_20394; // @[Switch.scala 30:36:@2310.4]
  assign _T_20397 = io_inAddr_16 == 6'h7; // @[Switch.scala 30:53:@2312.4]
  assign valid_7_16 = io_inValid_16 & _T_20397; // @[Switch.scala 30:36:@2313.4]
  assign _T_20400 = io_inAddr_17 == 6'h7; // @[Switch.scala 30:53:@2315.4]
  assign valid_7_17 = io_inValid_17 & _T_20400; // @[Switch.scala 30:36:@2316.4]
  assign _T_20403 = io_inAddr_18 == 6'h7; // @[Switch.scala 30:53:@2318.4]
  assign valid_7_18 = io_inValid_18 & _T_20403; // @[Switch.scala 30:36:@2319.4]
  assign _T_20406 = io_inAddr_19 == 6'h7; // @[Switch.scala 30:53:@2321.4]
  assign valid_7_19 = io_inValid_19 & _T_20406; // @[Switch.scala 30:36:@2322.4]
  assign _T_20409 = io_inAddr_20 == 6'h7; // @[Switch.scala 30:53:@2324.4]
  assign valid_7_20 = io_inValid_20 & _T_20409; // @[Switch.scala 30:36:@2325.4]
  assign _T_20412 = io_inAddr_21 == 6'h7; // @[Switch.scala 30:53:@2327.4]
  assign valid_7_21 = io_inValid_21 & _T_20412; // @[Switch.scala 30:36:@2328.4]
  assign _T_20415 = io_inAddr_22 == 6'h7; // @[Switch.scala 30:53:@2330.4]
  assign valid_7_22 = io_inValid_22 & _T_20415; // @[Switch.scala 30:36:@2331.4]
  assign _T_20418 = io_inAddr_23 == 6'h7; // @[Switch.scala 30:53:@2333.4]
  assign valid_7_23 = io_inValid_23 & _T_20418; // @[Switch.scala 30:36:@2334.4]
  assign _T_20421 = io_inAddr_24 == 6'h7; // @[Switch.scala 30:53:@2336.4]
  assign valid_7_24 = io_inValid_24 & _T_20421; // @[Switch.scala 30:36:@2337.4]
  assign _T_20424 = io_inAddr_25 == 6'h7; // @[Switch.scala 30:53:@2339.4]
  assign valid_7_25 = io_inValid_25 & _T_20424; // @[Switch.scala 30:36:@2340.4]
  assign _T_20427 = io_inAddr_26 == 6'h7; // @[Switch.scala 30:53:@2342.4]
  assign valid_7_26 = io_inValid_26 & _T_20427; // @[Switch.scala 30:36:@2343.4]
  assign _T_20430 = io_inAddr_27 == 6'h7; // @[Switch.scala 30:53:@2345.4]
  assign valid_7_27 = io_inValid_27 & _T_20430; // @[Switch.scala 30:36:@2346.4]
  assign _T_20433 = io_inAddr_28 == 6'h7; // @[Switch.scala 30:53:@2348.4]
  assign valid_7_28 = io_inValid_28 & _T_20433; // @[Switch.scala 30:36:@2349.4]
  assign _T_20436 = io_inAddr_29 == 6'h7; // @[Switch.scala 30:53:@2351.4]
  assign valid_7_29 = io_inValid_29 & _T_20436; // @[Switch.scala 30:36:@2352.4]
  assign _T_20439 = io_inAddr_30 == 6'h7; // @[Switch.scala 30:53:@2354.4]
  assign valid_7_30 = io_inValid_30 & _T_20439; // @[Switch.scala 30:36:@2355.4]
  assign _T_20442 = io_inAddr_31 == 6'h7; // @[Switch.scala 30:53:@2357.4]
  assign valid_7_31 = io_inValid_31 & _T_20442; // @[Switch.scala 30:36:@2358.4]
  assign _T_20445 = io_inAddr_32 == 6'h7; // @[Switch.scala 30:53:@2360.4]
  assign valid_7_32 = io_inValid_32 & _T_20445; // @[Switch.scala 30:36:@2361.4]
  assign _T_20448 = io_inAddr_33 == 6'h7; // @[Switch.scala 30:53:@2363.4]
  assign valid_7_33 = io_inValid_33 & _T_20448; // @[Switch.scala 30:36:@2364.4]
  assign _T_20451 = io_inAddr_34 == 6'h7; // @[Switch.scala 30:53:@2366.4]
  assign valid_7_34 = io_inValid_34 & _T_20451; // @[Switch.scala 30:36:@2367.4]
  assign _T_20454 = io_inAddr_35 == 6'h7; // @[Switch.scala 30:53:@2369.4]
  assign valid_7_35 = io_inValid_35 & _T_20454; // @[Switch.scala 30:36:@2370.4]
  assign _T_20457 = io_inAddr_36 == 6'h7; // @[Switch.scala 30:53:@2372.4]
  assign valid_7_36 = io_inValid_36 & _T_20457; // @[Switch.scala 30:36:@2373.4]
  assign _T_20460 = io_inAddr_37 == 6'h7; // @[Switch.scala 30:53:@2375.4]
  assign valid_7_37 = io_inValid_37 & _T_20460; // @[Switch.scala 30:36:@2376.4]
  assign _T_20463 = io_inAddr_38 == 6'h7; // @[Switch.scala 30:53:@2378.4]
  assign valid_7_38 = io_inValid_38 & _T_20463; // @[Switch.scala 30:36:@2379.4]
  assign _T_20466 = io_inAddr_39 == 6'h7; // @[Switch.scala 30:53:@2381.4]
  assign valid_7_39 = io_inValid_39 & _T_20466; // @[Switch.scala 30:36:@2382.4]
  assign _T_20469 = io_inAddr_40 == 6'h7; // @[Switch.scala 30:53:@2384.4]
  assign valid_7_40 = io_inValid_40 & _T_20469; // @[Switch.scala 30:36:@2385.4]
  assign _T_20472 = io_inAddr_41 == 6'h7; // @[Switch.scala 30:53:@2387.4]
  assign valid_7_41 = io_inValid_41 & _T_20472; // @[Switch.scala 30:36:@2388.4]
  assign _T_20475 = io_inAddr_42 == 6'h7; // @[Switch.scala 30:53:@2390.4]
  assign valid_7_42 = io_inValid_42 & _T_20475; // @[Switch.scala 30:36:@2391.4]
  assign _T_20478 = io_inAddr_43 == 6'h7; // @[Switch.scala 30:53:@2393.4]
  assign valid_7_43 = io_inValid_43 & _T_20478; // @[Switch.scala 30:36:@2394.4]
  assign _T_20481 = io_inAddr_44 == 6'h7; // @[Switch.scala 30:53:@2396.4]
  assign valid_7_44 = io_inValid_44 & _T_20481; // @[Switch.scala 30:36:@2397.4]
  assign _T_20484 = io_inAddr_45 == 6'h7; // @[Switch.scala 30:53:@2399.4]
  assign valid_7_45 = io_inValid_45 & _T_20484; // @[Switch.scala 30:36:@2400.4]
  assign _T_20487 = io_inAddr_46 == 6'h7; // @[Switch.scala 30:53:@2402.4]
  assign valid_7_46 = io_inValid_46 & _T_20487; // @[Switch.scala 30:36:@2403.4]
  assign _T_20490 = io_inAddr_47 == 6'h7; // @[Switch.scala 30:53:@2405.4]
  assign valid_7_47 = io_inValid_47 & _T_20490; // @[Switch.scala 30:36:@2406.4]
  assign _T_20493 = io_inAddr_48 == 6'h7; // @[Switch.scala 30:53:@2408.4]
  assign valid_7_48 = io_inValid_48 & _T_20493; // @[Switch.scala 30:36:@2409.4]
  assign _T_20496 = io_inAddr_49 == 6'h7; // @[Switch.scala 30:53:@2411.4]
  assign valid_7_49 = io_inValid_49 & _T_20496; // @[Switch.scala 30:36:@2412.4]
  assign _T_20499 = io_inAddr_50 == 6'h7; // @[Switch.scala 30:53:@2414.4]
  assign valid_7_50 = io_inValid_50 & _T_20499; // @[Switch.scala 30:36:@2415.4]
  assign _T_20502 = io_inAddr_51 == 6'h7; // @[Switch.scala 30:53:@2417.4]
  assign valid_7_51 = io_inValid_51 & _T_20502; // @[Switch.scala 30:36:@2418.4]
  assign _T_20505 = io_inAddr_52 == 6'h7; // @[Switch.scala 30:53:@2420.4]
  assign valid_7_52 = io_inValid_52 & _T_20505; // @[Switch.scala 30:36:@2421.4]
  assign _T_20508 = io_inAddr_53 == 6'h7; // @[Switch.scala 30:53:@2423.4]
  assign valid_7_53 = io_inValid_53 & _T_20508; // @[Switch.scala 30:36:@2424.4]
  assign _T_20511 = io_inAddr_54 == 6'h7; // @[Switch.scala 30:53:@2426.4]
  assign valid_7_54 = io_inValid_54 & _T_20511; // @[Switch.scala 30:36:@2427.4]
  assign _T_20514 = io_inAddr_55 == 6'h7; // @[Switch.scala 30:53:@2429.4]
  assign valid_7_55 = io_inValid_55 & _T_20514; // @[Switch.scala 30:36:@2430.4]
  assign _T_20517 = io_inAddr_56 == 6'h7; // @[Switch.scala 30:53:@2432.4]
  assign valid_7_56 = io_inValid_56 & _T_20517; // @[Switch.scala 30:36:@2433.4]
  assign _T_20520 = io_inAddr_57 == 6'h7; // @[Switch.scala 30:53:@2435.4]
  assign valid_7_57 = io_inValid_57 & _T_20520; // @[Switch.scala 30:36:@2436.4]
  assign _T_20523 = io_inAddr_58 == 6'h7; // @[Switch.scala 30:53:@2438.4]
  assign valid_7_58 = io_inValid_58 & _T_20523; // @[Switch.scala 30:36:@2439.4]
  assign _T_20526 = io_inAddr_59 == 6'h7; // @[Switch.scala 30:53:@2441.4]
  assign valid_7_59 = io_inValid_59 & _T_20526; // @[Switch.scala 30:36:@2442.4]
  assign _T_20529 = io_inAddr_60 == 6'h7; // @[Switch.scala 30:53:@2444.4]
  assign valid_7_60 = io_inValid_60 & _T_20529; // @[Switch.scala 30:36:@2445.4]
  assign _T_20532 = io_inAddr_61 == 6'h7; // @[Switch.scala 30:53:@2447.4]
  assign valid_7_61 = io_inValid_61 & _T_20532; // @[Switch.scala 30:36:@2448.4]
  assign _T_20535 = io_inAddr_62 == 6'h7; // @[Switch.scala 30:53:@2450.4]
  assign valid_7_62 = io_inValid_62 & _T_20535; // @[Switch.scala 30:36:@2451.4]
  assign _T_20538 = io_inAddr_63 == 6'h7; // @[Switch.scala 30:53:@2453.4]
  assign valid_7_63 = io_inValid_63 & _T_20538; // @[Switch.scala 30:36:@2454.4]
  assign _T_20604 = valid_7_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@2456.4]
  assign _T_20605 = valid_7_61 ? 6'h3d : _T_20604; // @[Mux.scala 31:69:@2457.4]
  assign _T_20606 = valid_7_60 ? 6'h3c : _T_20605; // @[Mux.scala 31:69:@2458.4]
  assign _T_20607 = valid_7_59 ? 6'h3b : _T_20606; // @[Mux.scala 31:69:@2459.4]
  assign _T_20608 = valid_7_58 ? 6'h3a : _T_20607; // @[Mux.scala 31:69:@2460.4]
  assign _T_20609 = valid_7_57 ? 6'h39 : _T_20608; // @[Mux.scala 31:69:@2461.4]
  assign _T_20610 = valid_7_56 ? 6'h38 : _T_20609; // @[Mux.scala 31:69:@2462.4]
  assign _T_20611 = valid_7_55 ? 6'h37 : _T_20610; // @[Mux.scala 31:69:@2463.4]
  assign _T_20612 = valid_7_54 ? 6'h36 : _T_20611; // @[Mux.scala 31:69:@2464.4]
  assign _T_20613 = valid_7_53 ? 6'h35 : _T_20612; // @[Mux.scala 31:69:@2465.4]
  assign _T_20614 = valid_7_52 ? 6'h34 : _T_20613; // @[Mux.scala 31:69:@2466.4]
  assign _T_20615 = valid_7_51 ? 6'h33 : _T_20614; // @[Mux.scala 31:69:@2467.4]
  assign _T_20616 = valid_7_50 ? 6'h32 : _T_20615; // @[Mux.scala 31:69:@2468.4]
  assign _T_20617 = valid_7_49 ? 6'h31 : _T_20616; // @[Mux.scala 31:69:@2469.4]
  assign _T_20618 = valid_7_48 ? 6'h30 : _T_20617; // @[Mux.scala 31:69:@2470.4]
  assign _T_20619 = valid_7_47 ? 6'h2f : _T_20618; // @[Mux.scala 31:69:@2471.4]
  assign _T_20620 = valid_7_46 ? 6'h2e : _T_20619; // @[Mux.scala 31:69:@2472.4]
  assign _T_20621 = valid_7_45 ? 6'h2d : _T_20620; // @[Mux.scala 31:69:@2473.4]
  assign _T_20622 = valid_7_44 ? 6'h2c : _T_20621; // @[Mux.scala 31:69:@2474.4]
  assign _T_20623 = valid_7_43 ? 6'h2b : _T_20622; // @[Mux.scala 31:69:@2475.4]
  assign _T_20624 = valid_7_42 ? 6'h2a : _T_20623; // @[Mux.scala 31:69:@2476.4]
  assign _T_20625 = valid_7_41 ? 6'h29 : _T_20624; // @[Mux.scala 31:69:@2477.4]
  assign _T_20626 = valid_7_40 ? 6'h28 : _T_20625; // @[Mux.scala 31:69:@2478.4]
  assign _T_20627 = valid_7_39 ? 6'h27 : _T_20626; // @[Mux.scala 31:69:@2479.4]
  assign _T_20628 = valid_7_38 ? 6'h26 : _T_20627; // @[Mux.scala 31:69:@2480.4]
  assign _T_20629 = valid_7_37 ? 6'h25 : _T_20628; // @[Mux.scala 31:69:@2481.4]
  assign _T_20630 = valid_7_36 ? 6'h24 : _T_20629; // @[Mux.scala 31:69:@2482.4]
  assign _T_20631 = valid_7_35 ? 6'h23 : _T_20630; // @[Mux.scala 31:69:@2483.4]
  assign _T_20632 = valid_7_34 ? 6'h22 : _T_20631; // @[Mux.scala 31:69:@2484.4]
  assign _T_20633 = valid_7_33 ? 6'h21 : _T_20632; // @[Mux.scala 31:69:@2485.4]
  assign _T_20634 = valid_7_32 ? 6'h20 : _T_20633; // @[Mux.scala 31:69:@2486.4]
  assign _T_20635 = valid_7_31 ? 6'h1f : _T_20634; // @[Mux.scala 31:69:@2487.4]
  assign _T_20636 = valid_7_30 ? 6'h1e : _T_20635; // @[Mux.scala 31:69:@2488.4]
  assign _T_20637 = valid_7_29 ? 6'h1d : _T_20636; // @[Mux.scala 31:69:@2489.4]
  assign _T_20638 = valid_7_28 ? 6'h1c : _T_20637; // @[Mux.scala 31:69:@2490.4]
  assign _T_20639 = valid_7_27 ? 6'h1b : _T_20638; // @[Mux.scala 31:69:@2491.4]
  assign _T_20640 = valid_7_26 ? 6'h1a : _T_20639; // @[Mux.scala 31:69:@2492.4]
  assign _T_20641 = valid_7_25 ? 6'h19 : _T_20640; // @[Mux.scala 31:69:@2493.4]
  assign _T_20642 = valid_7_24 ? 6'h18 : _T_20641; // @[Mux.scala 31:69:@2494.4]
  assign _T_20643 = valid_7_23 ? 6'h17 : _T_20642; // @[Mux.scala 31:69:@2495.4]
  assign _T_20644 = valid_7_22 ? 6'h16 : _T_20643; // @[Mux.scala 31:69:@2496.4]
  assign _T_20645 = valid_7_21 ? 6'h15 : _T_20644; // @[Mux.scala 31:69:@2497.4]
  assign _T_20646 = valid_7_20 ? 6'h14 : _T_20645; // @[Mux.scala 31:69:@2498.4]
  assign _T_20647 = valid_7_19 ? 6'h13 : _T_20646; // @[Mux.scala 31:69:@2499.4]
  assign _T_20648 = valid_7_18 ? 6'h12 : _T_20647; // @[Mux.scala 31:69:@2500.4]
  assign _T_20649 = valid_7_17 ? 6'h11 : _T_20648; // @[Mux.scala 31:69:@2501.4]
  assign _T_20650 = valid_7_16 ? 6'h10 : _T_20649; // @[Mux.scala 31:69:@2502.4]
  assign _T_20651 = valid_7_15 ? 6'hf : _T_20650; // @[Mux.scala 31:69:@2503.4]
  assign _T_20652 = valid_7_14 ? 6'he : _T_20651; // @[Mux.scala 31:69:@2504.4]
  assign _T_20653 = valid_7_13 ? 6'hd : _T_20652; // @[Mux.scala 31:69:@2505.4]
  assign _T_20654 = valid_7_12 ? 6'hc : _T_20653; // @[Mux.scala 31:69:@2506.4]
  assign _T_20655 = valid_7_11 ? 6'hb : _T_20654; // @[Mux.scala 31:69:@2507.4]
  assign _T_20656 = valid_7_10 ? 6'ha : _T_20655; // @[Mux.scala 31:69:@2508.4]
  assign _T_20657 = valid_7_9 ? 6'h9 : _T_20656; // @[Mux.scala 31:69:@2509.4]
  assign _T_20658 = valid_7_8 ? 6'h8 : _T_20657; // @[Mux.scala 31:69:@2510.4]
  assign _T_20659 = valid_7_7 ? 6'h7 : _T_20658; // @[Mux.scala 31:69:@2511.4]
  assign _T_20660 = valid_7_6 ? 6'h6 : _T_20659; // @[Mux.scala 31:69:@2512.4]
  assign _T_20661 = valid_7_5 ? 6'h5 : _T_20660; // @[Mux.scala 31:69:@2513.4]
  assign _T_20662 = valid_7_4 ? 6'h4 : _T_20661; // @[Mux.scala 31:69:@2514.4]
  assign _T_20663 = valid_7_3 ? 6'h3 : _T_20662; // @[Mux.scala 31:69:@2515.4]
  assign _T_20664 = valid_7_2 ? 6'h2 : _T_20663; // @[Mux.scala 31:69:@2516.4]
  assign _T_20665 = valid_7_1 ? 6'h1 : _T_20664; // @[Mux.scala 31:69:@2517.4]
  assign select_7 = valid_7_0 ? 6'h0 : _T_20665; // @[Mux.scala 31:69:@2518.4]
  assign _GEN_449 = 6'h1 == select_7 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_450 = 6'h2 == select_7 ? io_inData_2 : _GEN_449; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_451 = 6'h3 == select_7 ? io_inData_3 : _GEN_450; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_452 = 6'h4 == select_7 ? io_inData_4 : _GEN_451; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_453 = 6'h5 == select_7 ? io_inData_5 : _GEN_452; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_454 = 6'h6 == select_7 ? io_inData_6 : _GEN_453; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_455 = 6'h7 == select_7 ? io_inData_7 : _GEN_454; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_456 = 6'h8 == select_7 ? io_inData_8 : _GEN_455; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_457 = 6'h9 == select_7 ? io_inData_9 : _GEN_456; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_458 = 6'ha == select_7 ? io_inData_10 : _GEN_457; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_459 = 6'hb == select_7 ? io_inData_11 : _GEN_458; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_460 = 6'hc == select_7 ? io_inData_12 : _GEN_459; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_461 = 6'hd == select_7 ? io_inData_13 : _GEN_460; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_462 = 6'he == select_7 ? io_inData_14 : _GEN_461; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_463 = 6'hf == select_7 ? io_inData_15 : _GEN_462; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_464 = 6'h10 == select_7 ? io_inData_16 : _GEN_463; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_465 = 6'h11 == select_7 ? io_inData_17 : _GEN_464; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_466 = 6'h12 == select_7 ? io_inData_18 : _GEN_465; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_467 = 6'h13 == select_7 ? io_inData_19 : _GEN_466; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_468 = 6'h14 == select_7 ? io_inData_20 : _GEN_467; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_469 = 6'h15 == select_7 ? io_inData_21 : _GEN_468; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_470 = 6'h16 == select_7 ? io_inData_22 : _GEN_469; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_471 = 6'h17 == select_7 ? io_inData_23 : _GEN_470; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_472 = 6'h18 == select_7 ? io_inData_24 : _GEN_471; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_473 = 6'h19 == select_7 ? io_inData_25 : _GEN_472; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_474 = 6'h1a == select_7 ? io_inData_26 : _GEN_473; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_475 = 6'h1b == select_7 ? io_inData_27 : _GEN_474; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_476 = 6'h1c == select_7 ? io_inData_28 : _GEN_475; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_477 = 6'h1d == select_7 ? io_inData_29 : _GEN_476; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_478 = 6'h1e == select_7 ? io_inData_30 : _GEN_477; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_479 = 6'h1f == select_7 ? io_inData_31 : _GEN_478; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_480 = 6'h20 == select_7 ? io_inData_32 : _GEN_479; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_481 = 6'h21 == select_7 ? io_inData_33 : _GEN_480; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_482 = 6'h22 == select_7 ? io_inData_34 : _GEN_481; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_483 = 6'h23 == select_7 ? io_inData_35 : _GEN_482; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_484 = 6'h24 == select_7 ? io_inData_36 : _GEN_483; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_485 = 6'h25 == select_7 ? io_inData_37 : _GEN_484; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_486 = 6'h26 == select_7 ? io_inData_38 : _GEN_485; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_487 = 6'h27 == select_7 ? io_inData_39 : _GEN_486; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_488 = 6'h28 == select_7 ? io_inData_40 : _GEN_487; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_489 = 6'h29 == select_7 ? io_inData_41 : _GEN_488; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_490 = 6'h2a == select_7 ? io_inData_42 : _GEN_489; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_491 = 6'h2b == select_7 ? io_inData_43 : _GEN_490; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_492 = 6'h2c == select_7 ? io_inData_44 : _GEN_491; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_493 = 6'h2d == select_7 ? io_inData_45 : _GEN_492; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_494 = 6'h2e == select_7 ? io_inData_46 : _GEN_493; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_495 = 6'h2f == select_7 ? io_inData_47 : _GEN_494; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_496 = 6'h30 == select_7 ? io_inData_48 : _GEN_495; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_497 = 6'h31 == select_7 ? io_inData_49 : _GEN_496; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_498 = 6'h32 == select_7 ? io_inData_50 : _GEN_497; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_499 = 6'h33 == select_7 ? io_inData_51 : _GEN_498; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_500 = 6'h34 == select_7 ? io_inData_52 : _GEN_499; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_501 = 6'h35 == select_7 ? io_inData_53 : _GEN_500; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_502 = 6'h36 == select_7 ? io_inData_54 : _GEN_501; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_503 = 6'h37 == select_7 ? io_inData_55 : _GEN_502; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_504 = 6'h38 == select_7 ? io_inData_56 : _GEN_503; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_505 = 6'h39 == select_7 ? io_inData_57 : _GEN_504; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_506 = 6'h3a == select_7 ? io_inData_58 : _GEN_505; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_507 = 6'h3b == select_7 ? io_inData_59 : _GEN_506; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_508 = 6'h3c == select_7 ? io_inData_60 : _GEN_507; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_509 = 6'h3d == select_7 ? io_inData_61 : _GEN_508; // @[Switch.scala 33:19:@2520.4]
  assign _GEN_510 = 6'h3e == select_7 ? io_inData_62 : _GEN_509; // @[Switch.scala 33:19:@2520.4]
  assign _T_20674 = {valid_7_7,valid_7_6,valid_7_5,valid_7_4,valid_7_3,valid_7_2,valid_7_1,valid_7_0}; // @[Switch.scala 34:32:@2527.4]
  assign _T_20682 = {valid_7_15,valid_7_14,valid_7_13,valid_7_12,valid_7_11,valid_7_10,valid_7_9,valid_7_8,_T_20674}; // @[Switch.scala 34:32:@2535.4]
  assign _T_20689 = {valid_7_23,valid_7_22,valid_7_21,valid_7_20,valid_7_19,valid_7_18,valid_7_17,valid_7_16}; // @[Switch.scala 34:32:@2542.4]
  assign _T_20698 = {valid_7_31,valid_7_30,valid_7_29,valid_7_28,valid_7_27,valid_7_26,valid_7_25,valid_7_24,_T_20689,_T_20682}; // @[Switch.scala 34:32:@2551.4]
  assign _T_20705 = {valid_7_39,valid_7_38,valid_7_37,valid_7_36,valid_7_35,valid_7_34,valid_7_33,valid_7_32}; // @[Switch.scala 34:32:@2558.4]
  assign _T_20713 = {valid_7_47,valid_7_46,valid_7_45,valid_7_44,valid_7_43,valid_7_42,valid_7_41,valid_7_40,_T_20705}; // @[Switch.scala 34:32:@2566.4]
  assign _T_20720 = {valid_7_55,valid_7_54,valid_7_53,valid_7_52,valid_7_51,valid_7_50,valid_7_49,valid_7_48}; // @[Switch.scala 34:32:@2573.4]
  assign _T_20729 = {valid_7_63,valid_7_62,valid_7_61,valid_7_60,valid_7_59,valid_7_58,valid_7_57,valid_7_56,_T_20720,_T_20713}; // @[Switch.scala 34:32:@2582.4]
  assign _T_20730 = {_T_20729,_T_20698}; // @[Switch.scala 34:32:@2583.4]
  assign _T_20734 = io_inAddr_0 == 6'h8; // @[Switch.scala 30:53:@2586.4]
  assign valid_8_0 = io_inValid_0 & _T_20734; // @[Switch.scala 30:36:@2587.4]
  assign _T_20737 = io_inAddr_1 == 6'h8; // @[Switch.scala 30:53:@2589.4]
  assign valid_8_1 = io_inValid_1 & _T_20737; // @[Switch.scala 30:36:@2590.4]
  assign _T_20740 = io_inAddr_2 == 6'h8; // @[Switch.scala 30:53:@2592.4]
  assign valid_8_2 = io_inValid_2 & _T_20740; // @[Switch.scala 30:36:@2593.4]
  assign _T_20743 = io_inAddr_3 == 6'h8; // @[Switch.scala 30:53:@2595.4]
  assign valid_8_3 = io_inValid_3 & _T_20743; // @[Switch.scala 30:36:@2596.4]
  assign _T_20746 = io_inAddr_4 == 6'h8; // @[Switch.scala 30:53:@2598.4]
  assign valid_8_4 = io_inValid_4 & _T_20746; // @[Switch.scala 30:36:@2599.4]
  assign _T_20749 = io_inAddr_5 == 6'h8; // @[Switch.scala 30:53:@2601.4]
  assign valid_8_5 = io_inValid_5 & _T_20749; // @[Switch.scala 30:36:@2602.4]
  assign _T_20752 = io_inAddr_6 == 6'h8; // @[Switch.scala 30:53:@2604.4]
  assign valid_8_6 = io_inValid_6 & _T_20752; // @[Switch.scala 30:36:@2605.4]
  assign _T_20755 = io_inAddr_7 == 6'h8; // @[Switch.scala 30:53:@2607.4]
  assign valid_8_7 = io_inValid_7 & _T_20755; // @[Switch.scala 30:36:@2608.4]
  assign _T_20758 = io_inAddr_8 == 6'h8; // @[Switch.scala 30:53:@2610.4]
  assign valid_8_8 = io_inValid_8 & _T_20758; // @[Switch.scala 30:36:@2611.4]
  assign _T_20761 = io_inAddr_9 == 6'h8; // @[Switch.scala 30:53:@2613.4]
  assign valid_8_9 = io_inValid_9 & _T_20761; // @[Switch.scala 30:36:@2614.4]
  assign _T_20764 = io_inAddr_10 == 6'h8; // @[Switch.scala 30:53:@2616.4]
  assign valid_8_10 = io_inValid_10 & _T_20764; // @[Switch.scala 30:36:@2617.4]
  assign _T_20767 = io_inAddr_11 == 6'h8; // @[Switch.scala 30:53:@2619.4]
  assign valid_8_11 = io_inValid_11 & _T_20767; // @[Switch.scala 30:36:@2620.4]
  assign _T_20770 = io_inAddr_12 == 6'h8; // @[Switch.scala 30:53:@2622.4]
  assign valid_8_12 = io_inValid_12 & _T_20770; // @[Switch.scala 30:36:@2623.4]
  assign _T_20773 = io_inAddr_13 == 6'h8; // @[Switch.scala 30:53:@2625.4]
  assign valid_8_13 = io_inValid_13 & _T_20773; // @[Switch.scala 30:36:@2626.4]
  assign _T_20776 = io_inAddr_14 == 6'h8; // @[Switch.scala 30:53:@2628.4]
  assign valid_8_14 = io_inValid_14 & _T_20776; // @[Switch.scala 30:36:@2629.4]
  assign _T_20779 = io_inAddr_15 == 6'h8; // @[Switch.scala 30:53:@2631.4]
  assign valid_8_15 = io_inValid_15 & _T_20779; // @[Switch.scala 30:36:@2632.4]
  assign _T_20782 = io_inAddr_16 == 6'h8; // @[Switch.scala 30:53:@2634.4]
  assign valid_8_16 = io_inValid_16 & _T_20782; // @[Switch.scala 30:36:@2635.4]
  assign _T_20785 = io_inAddr_17 == 6'h8; // @[Switch.scala 30:53:@2637.4]
  assign valid_8_17 = io_inValid_17 & _T_20785; // @[Switch.scala 30:36:@2638.4]
  assign _T_20788 = io_inAddr_18 == 6'h8; // @[Switch.scala 30:53:@2640.4]
  assign valid_8_18 = io_inValid_18 & _T_20788; // @[Switch.scala 30:36:@2641.4]
  assign _T_20791 = io_inAddr_19 == 6'h8; // @[Switch.scala 30:53:@2643.4]
  assign valid_8_19 = io_inValid_19 & _T_20791; // @[Switch.scala 30:36:@2644.4]
  assign _T_20794 = io_inAddr_20 == 6'h8; // @[Switch.scala 30:53:@2646.4]
  assign valid_8_20 = io_inValid_20 & _T_20794; // @[Switch.scala 30:36:@2647.4]
  assign _T_20797 = io_inAddr_21 == 6'h8; // @[Switch.scala 30:53:@2649.4]
  assign valid_8_21 = io_inValid_21 & _T_20797; // @[Switch.scala 30:36:@2650.4]
  assign _T_20800 = io_inAddr_22 == 6'h8; // @[Switch.scala 30:53:@2652.4]
  assign valid_8_22 = io_inValid_22 & _T_20800; // @[Switch.scala 30:36:@2653.4]
  assign _T_20803 = io_inAddr_23 == 6'h8; // @[Switch.scala 30:53:@2655.4]
  assign valid_8_23 = io_inValid_23 & _T_20803; // @[Switch.scala 30:36:@2656.4]
  assign _T_20806 = io_inAddr_24 == 6'h8; // @[Switch.scala 30:53:@2658.4]
  assign valid_8_24 = io_inValid_24 & _T_20806; // @[Switch.scala 30:36:@2659.4]
  assign _T_20809 = io_inAddr_25 == 6'h8; // @[Switch.scala 30:53:@2661.4]
  assign valid_8_25 = io_inValid_25 & _T_20809; // @[Switch.scala 30:36:@2662.4]
  assign _T_20812 = io_inAddr_26 == 6'h8; // @[Switch.scala 30:53:@2664.4]
  assign valid_8_26 = io_inValid_26 & _T_20812; // @[Switch.scala 30:36:@2665.4]
  assign _T_20815 = io_inAddr_27 == 6'h8; // @[Switch.scala 30:53:@2667.4]
  assign valid_8_27 = io_inValid_27 & _T_20815; // @[Switch.scala 30:36:@2668.4]
  assign _T_20818 = io_inAddr_28 == 6'h8; // @[Switch.scala 30:53:@2670.4]
  assign valid_8_28 = io_inValid_28 & _T_20818; // @[Switch.scala 30:36:@2671.4]
  assign _T_20821 = io_inAddr_29 == 6'h8; // @[Switch.scala 30:53:@2673.4]
  assign valid_8_29 = io_inValid_29 & _T_20821; // @[Switch.scala 30:36:@2674.4]
  assign _T_20824 = io_inAddr_30 == 6'h8; // @[Switch.scala 30:53:@2676.4]
  assign valid_8_30 = io_inValid_30 & _T_20824; // @[Switch.scala 30:36:@2677.4]
  assign _T_20827 = io_inAddr_31 == 6'h8; // @[Switch.scala 30:53:@2679.4]
  assign valid_8_31 = io_inValid_31 & _T_20827; // @[Switch.scala 30:36:@2680.4]
  assign _T_20830 = io_inAddr_32 == 6'h8; // @[Switch.scala 30:53:@2682.4]
  assign valid_8_32 = io_inValid_32 & _T_20830; // @[Switch.scala 30:36:@2683.4]
  assign _T_20833 = io_inAddr_33 == 6'h8; // @[Switch.scala 30:53:@2685.4]
  assign valid_8_33 = io_inValid_33 & _T_20833; // @[Switch.scala 30:36:@2686.4]
  assign _T_20836 = io_inAddr_34 == 6'h8; // @[Switch.scala 30:53:@2688.4]
  assign valid_8_34 = io_inValid_34 & _T_20836; // @[Switch.scala 30:36:@2689.4]
  assign _T_20839 = io_inAddr_35 == 6'h8; // @[Switch.scala 30:53:@2691.4]
  assign valid_8_35 = io_inValid_35 & _T_20839; // @[Switch.scala 30:36:@2692.4]
  assign _T_20842 = io_inAddr_36 == 6'h8; // @[Switch.scala 30:53:@2694.4]
  assign valid_8_36 = io_inValid_36 & _T_20842; // @[Switch.scala 30:36:@2695.4]
  assign _T_20845 = io_inAddr_37 == 6'h8; // @[Switch.scala 30:53:@2697.4]
  assign valid_8_37 = io_inValid_37 & _T_20845; // @[Switch.scala 30:36:@2698.4]
  assign _T_20848 = io_inAddr_38 == 6'h8; // @[Switch.scala 30:53:@2700.4]
  assign valid_8_38 = io_inValid_38 & _T_20848; // @[Switch.scala 30:36:@2701.4]
  assign _T_20851 = io_inAddr_39 == 6'h8; // @[Switch.scala 30:53:@2703.4]
  assign valid_8_39 = io_inValid_39 & _T_20851; // @[Switch.scala 30:36:@2704.4]
  assign _T_20854 = io_inAddr_40 == 6'h8; // @[Switch.scala 30:53:@2706.4]
  assign valid_8_40 = io_inValid_40 & _T_20854; // @[Switch.scala 30:36:@2707.4]
  assign _T_20857 = io_inAddr_41 == 6'h8; // @[Switch.scala 30:53:@2709.4]
  assign valid_8_41 = io_inValid_41 & _T_20857; // @[Switch.scala 30:36:@2710.4]
  assign _T_20860 = io_inAddr_42 == 6'h8; // @[Switch.scala 30:53:@2712.4]
  assign valid_8_42 = io_inValid_42 & _T_20860; // @[Switch.scala 30:36:@2713.4]
  assign _T_20863 = io_inAddr_43 == 6'h8; // @[Switch.scala 30:53:@2715.4]
  assign valid_8_43 = io_inValid_43 & _T_20863; // @[Switch.scala 30:36:@2716.4]
  assign _T_20866 = io_inAddr_44 == 6'h8; // @[Switch.scala 30:53:@2718.4]
  assign valid_8_44 = io_inValid_44 & _T_20866; // @[Switch.scala 30:36:@2719.4]
  assign _T_20869 = io_inAddr_45 == 6'h8; // @[Switch.scala 30:53:@2721.4]
  assign valid_8_45 = io_inValid_45 & _T_20869; // @[Switch.scala 30:36:@2722.4]
  assign _T_20872 = io_inAddr_46 == 6'h8; // @[Switch.scala 30:53:@2724.4]
  assign valid_8_46 = io_inValid_46 & _T_20872; // @[Switch.scala 30:36:@2725.4]
  assign _T_20875 = io_inAddr_47 == 6'h8; // @[Switch.scala 30:53:@2727.4]
  assign valid_8_47 = io_inValid_47 & _T_20875; // @[Switch.scala 30:36:@2728.4]
  assign _T_20878 = io_inAddr_48 == 6'h8; // @[Switch.scala 30:53:@2730.4]
  assign valid_8_48 = io_inValid_48 & _T_20878; // @[Switch.scala 30:36:@2731.4]
  assign _T_20881 = io_inAddr_49 == 6'h8; // @[Switch.scala 30:53:@2733.4]
  assign valid_8_49 = io_inValid_49 & _T_20881; // @[Switch.scala 30:36:@2734.4]
  assign _T_20884 = io_inAddr_50 == 6'h8; // @[Switch.scala 30:53:@2736.4]
  assign valid_8_50 = io_inValid_50 & _T_20884; // @[Switch.scala 30:36:@2737.4]
  assign _T_20887 = io_inAddr_51 == 6'h8; // @[Switch.scala 30:53:@2739.4]
  assign valid_8_51 = io_inValid_51 & _T_20887; // @[Switch.scala 30:36:@2740.4]
  assign _T_20890 = io_inAddr_52 == 6'h8; // @[Switch.scala 30:53:@2742.4]
  assign valid_8_52 = io_inValid_52 & _T_20890; // @[Switch.scala 30:36:@2743.4]
  assign _T_20893 = io_inAddr_53 == 6'h8; // @[Switch.scala 30:53:@2745.4]
  assign valid_8_53 = io_inValid_53 & _T_20893; // @[Switch.scala 30:36:@2746.4]
  assign _T_20896 = io_inAddr_54 == 6'h8; // @[Switch.scala 30:53:@2748.4]
  assign valid_8_54 = io_inValid_54 & _T_20896; // @[Switch.scala 30:36:@2749.4]
  assign _T_20899 = io_inAddr_55 == 6'h8; // @[Switch.scala 30:53:@2751.4]
  assign valid_8_55 = io_inValid_55 & _T_20899; // @[Switch.scala 30:36:@2752.4]
  assign _T_20902 = io_inAddr_56 == 6'h8; // @[Switch.scala 30:53:@2754.4]
  assign valid_8_56 = io_inValid_56 & _T_20902; // @[Switch.scala 30:36:@2755.4]
  assign _T_20905 = io_inAddr_57 == 6'h8; // @[Switch.scala 30:53:@2757.4]
  assign valid_8_57 = io_inValid_57 & _T_20905; // @[Switch.scala 30:36:@2758.4]
  assign _T_20908 = io_inAddr_58 == 6'h8; // @[Switch.scala 30:53:@2760.4]
  assign valid_8_58 = io_inValid_58 & _T_20908; // @[Switch.scala 30:36:@2761.4]
  assign _T_20911 = io_inAddr_59 == 6'h8; // @[Switch.scala 30:53:@2763.4]
  assign valid_8_59 = io_inValid_59 & _T_20911; // @[Switch.scala 30:36:@2764.4]
  assign _T_20914 = io_inAddr_60 == 6'h8; // @[Switch.scala 30:53:@2766.4]
  assign valid_8_60 = io_inValid_60 & _T_20914; // @[Switch.scala 30:36:@2767.4]
  assign _T_20917 = io_inAddr_61 == 6'h8; // @[Switch.scala 30:53:@2769.4]
  assign valid_8_61 = io_inValid_61 & _T_20917; // @[Switch.scala 30:36:@2770.4]
  assign _T_20920 = io_inAddr_62 == 6'h8; // @[Switch.scala 30:53:@2772.4]
  assign valid_8_62 = io_inValid_62 & _T_20920; // @[Switch.scala 30:36:@2773.4]
  assign _T_20923 = io_inAddr_63 == 6'h8; // @[Switch.scala 30:53:@2775.4]
  assign valid_8_63 = io_inValid_63 & _T_20923; // @[Switch.scala 30:36:@2776.4]
  assign _T_20989 = valid_8_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@2778.4]
  assign _T_20990 = valid_8_61 ? 6'h3d : _T_20989; // @[Mux.scala 31:69:@2779.4]
  assign _T_20991 = valid_8_60 ? 6'h3c : _T_20990; // @[Mux.scala 31:69:@2780.4]
  assign _T_20992 = valid_8_59 ? 6'h3b : _T_20991; // @[Mux.scala 31:69:@2781.4]
  assign _T_20993 = valid_8_58 ? 6'h3a : _T_20992; // @[Mux.scala 31:69:@2782.4]
  assign _T_20994 = valid_8_57 ? 6'h39 : _T_20993; // @[Mux.scala 31:69:@2783.4]
  assign _T_20995 = valid_8_56 ? 6'h38 : _T_20994; // @[Mux.scala 31:69:@2784.4]
  assign _T_20996 = valid_8_55 ? 6'h37 : _T_20995; // @[Mux.scala 31:69:@2785.4]
  assign _T_20997 = valid_8_54 ? 6'h36 : _T_20996; // @[Mux.scala 31:69:@2786.4]
  assign _T_20998 = valid_8_53 ? 6'h35 : _T_20997; // @[Mux.scala 31:69:@2787.4]
  assign _T_20999 = valid_8_52 ? 6'h34 : _T_20998; // @[Mux.scala 31:69:@2788.4]
  assign _T_21000 = valid_8_51 ? 6'h33 : _T_20999; // @[Mux.scala 31:69:@2789.4]
  assign _T_21001 = valid_8_50 ? 6'h32 : _T_21000; // @[Mux.scala 31:69:@2790.4]
  assign _T_21002 = valid_8_49 ? 6'h31 : _T_21001; // @[Mux.scala 31:69:@2791.4]
  assign _T_21003 = valid_8_48 ? 6'h30 : _T_21002; // @[Mux.scala 31:69:@2792.4]
  assign _T_21004 = valid_8_47 ? 6'h2f : _T_21003; // @[Mux.scala 31:69:@2793.4]
  assign _T_21005 = valid_8_46 ? 6'h2e : _T_21004; // @[Mux.scala 31:69:@2794.4]
  assign _T_21006 = valid_8_45 ? 6'h2d : _T_21005; // @[Mux.scala 31:69:@2795.4]
  assign _T_21007 = valid_8_44 ? 6'h2c : _T_21006; // @[Mux.scala 31:69:@2796.4]
  assign _T_21008 = valid_8_43 ? 6'h2b : _T_21007; // @[Mux.scala 31:69:@2797.4]
  assign _T_21009 = valid_8_42 ? 6'h2a : _T_21008; // @[Mux.scala 31:69:@2798.4]
  assign _T_21010 = valid_8_41 ? 6'h29 : _T_21009; // @[Mux.scala 31:69:@2799.4]
  assign _T_21011 = valid_8_40 ? 6'h28 : _T_21010; // @[Mux.scala 31:69:@2800.4]
  assign _T_21012 = valid_8_39 ? 6'h27 : _T_21011; // @[Mux.scala 31:69:@2801.4]
  assign _T_21013 = valid_8_38 ? 6'h26 : _T_21012; // @[Mux.scala 31:69:@2802.4]
  assign _T_21014 = valid_8_37 ? 6'h25 : _T_21013; // @[Mux.scala 31:69:@2803.4]
  assign _T_21015 = valid_8_36 ? 6'h24 : _T_21014; // @[Mux.scala 31:69:@2804.4]
  assign _T_21016 = valid_8_35 ? 6'h23 : _T_21015; // @[Mux.scala 31:69:@2805.4]
  assign _T_21017 = valid_8_34 ? 6'h22 : _T_21016; // @[Mux.scala 31:69:@2806.4]
  assign _T_21018 = valid_8_33 ? 6'h21 : _T_21017; // @[Mux.scala 31:69:@2807.4]
  assign _T_21019 = valid_8_32 ? 6'h20 : _T_21018; // @[Mux.scala 31:69:@2808.4]
  assign _T_21020 = valid_8_31 ? 6'h1f : _T_21019; // @[Mux.scala 31:69:@2809.4]
  assign _T_21021 = valid_8_30 ? 6'h1e : _T_21020; // @[Mux.scala 31:69:@2810.4]
  assign _T_21022 = valid_8_29 ? 6'h1d : _T_21021; // @[Mux.scala 31:69:@2811.4]
  assign _T_21023 = valid_8_28 ? 6'h1c : _T_21022; // @[Mux.scala 31:69:@2812.4]
  assign _T_21024 = valid_8_27 ? 6'h1b : _T_21023; // @[Mux.scala 31:69:@2813.4]
  assign _T_21025 = valid_8_26 ? 6'h1a : _T_21024; // @[Mux.scala 31:69:@2814.4]
  assign _T_21026 = valid_8_25 ? 6'h19 : _T_21025; // @[Mux.scala 31:69:@2815.4]
  assign _T_21027 = valid_8_24 ? 6'h18 : _T_21026; // @[Mux.scala 31:69:@2816.4]
  assign _T_21028 = valid_8_23 ? 6'h17 : _T_21027; // @[Mux.scala 31:69:@2817.4]
  assign _T_21029 = valid_8_22 ? 6'h16 : _T_21028; // @[Mux.scala 31:69:@2818.4]
  assign _T_21030 = valid_8_21 ? 6'h15 : _T_21029; // @[Mux.scala 31:69:@2819.4]
  assign _T_21031 = valid_8_20 ? 6'h14 : _T_21030; // @[Mux.scala 31:69:@2820.4]
  assign _T_21032 = valid_8_19 ? 6'h13 : _T_21031; // @[Mux.scala 31:69:@2821.4]
  assign _T_21033 = valid_8_18 ? 6'h12 : _T_21032; // @[Mux.scala 31:69:@2822.4]
  assign _T_21034 = valid_8_17 ? 6'h11 : _T_21033; // @[Mux.scala 31:69:@2823.4]
  assign _T_21035 = valid_8_16 ? 6'h10 : _T_21034; // @[Mux.scala 31:69:@2824.4]
  assign _T_21036 = valid_8_15 ? 6'hf : _T_21035; // @[Mux.scala 31:69:@2825.4]
  assign _T_21037 = valid_8_14 ? 6'he : _T_21036; // @[Mux.scala 31:69:@2826.4]
  assign _T_21038 = valid_8_13 ? 6'hd : _T_21037; // @[Mux.scala 31:69:@2827.4]
  assign _T_21039 = valid_8_12 ? 6'hc : _T_21038; // @[Mux.scala 31:69:@2828.4]
  assign _T_21040 = valid_8_11 ? 6'hb : _T_21039; // @[Mux.scala 31:69:@2829.4]
  assign _T_21041 = valid_8_10 ? 6'ha : _T_21040; // @[Mux.scala 31:69:@2830.4]
  assign _T_21042 = valid_8_9 ? 6'h9 : _T_21041; // @[Mux.scala 31:69:@2831.4]
  assign _T_21043 = valid_8_8 ? 6'h8 : _T_21042; // @[Mux.scala 31:69:@2832.4]
  assign _T_21044 = valid_8_7 ? 6'h7 : _T_21043; // @[Mux.scala 31:69:@2833.4]
  assign _T_21045 = valid_8_6 ? 6'h6 : _T_21044; // @[Mux.scala 31:69:@2834.4]
  assign _T_21046 = valid_8_5 ? 6'h5 : _T_21045; // @[Mux.scala 31:69:@2835.4]
  assign _T_21047 = valid_8_4 ? 6'h4 : _T_21046; // @[Mux.scala 31:69:@2836.4]
  assign _T_21048 = valid_8_3 ? 6'h3 : _T_21047; // @[Mux.scala 31:69:@2837.4]
  assign _T_21049 = valid_8_2 ? 6'h2 : _T_21048; // @[Mux.scala 31:69:@2838.4]
  assign _T_21050 = valid_8_1 ? 6'h1 : _T_21049; // @[Mux.scala 31:69:@2839.4]
  assign select_8 = valid_8_0 ? 6'h0 : _T_21050; // @[Mux.scala 31:69:@2840.4]
  assign _GEN_513 = 6'h1 == select_8 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_514 = 6'h2 == select_8 ? io_inData_2 : _GEN_513; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_515 = 6'h3 == select_8 ? io_inData_3 : _GEN_514; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_516 = 6'h4 == select_8 ? io_inData_4 : _GEN_515; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_517 = 6'h5 == select_8 ? io_inData_5 : _GEN_516; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_518 = 6'h6 == select_8 ? io_inData_6 : _GEN_517; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_519 = 6'h7 == select_8 ? io_inData_7 : _GEN_518; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_520 = 6'h8 == select_8 ? io_inData_8 : _GEN_519; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_521 = 6'h9 == select_8 ? io_inData_9 : _GEN_520; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_522 = 6'ha == select_8 ? io_inData_10 : _GEN_521; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_523 = 6'hb == select_8 ? io_inData_11 : _GEN_522; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_524 = 6'hc == select_8 ? io_inData_12 : _GEN_523; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_525 = 6'hd == select_8 ? io_inData_13 : _GEN_524; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_526 = 6'he == select_8 ? io_inData_14 : _GEN_525; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_527 = 6'hf == select_8 ? io_inData_15 : _GEN_526; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_528 = 6'h10 == select_8 ? io_inData_16 : _GEN_527; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_529 = 6'h11 == select_8 ? io_inData_17 : _GEN_528; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_530 = 6'h12 == select_8 ? io_inData_18 : _GEN_529; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_531 = 6'h13 == select_8 ? io_inData_19 : _GEN_530; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_532 = 6'h14 == select_8 ? io_inData_20 : _GEN_531; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_533 = 6'h15 == select_8 ? io_inData_21 : _GEN_532; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_534 = 6'h16 == select_8 ? io_inData_22 : _GEN_533; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_535 = 6'h17 == select_8 ? io_inData_23 : _GEN_534; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_536 = 6'h18 == select_8 ? io_inData_24 : _GEN_535; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_537 = 6'h19 == select_8 ? io_inData_25 : _GEN_536; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_538 = 6'h1a == select_8 ? io_inData_26 : _GEN_537; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_539 = 6'h1b == select_8 ? io_inData_27 : _GEN_538; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_540 = 6'h1c == select_8 ? io_inData_28 : _GEN_539; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_541 = 6'h1d == select_8 ? io_inData_29 : _GEN_540; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_542 = 6'h1e == select_8 ? io_inData_30 : _GEN_541; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_543 = 6'h1f == select_8 ? io_inData_31 : _GEN_542; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_544 = 6'h20 == select_8 ? io_inData_32 : _GEN_543; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_545 = 6'h21 == select_8 ? io_inData_33 : _GEN_544; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_546 = 6'h22 == select_8 ? io_inData_34 : _GEN_545; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_547 = 6'h23 == select_8 ? io_inData_35 : _GEN_546; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_548 = 6'h24 == select_8 ? io_inData_36 : _GEN_547; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_549 = 6'h25 == select_8 ? io_inData_37 : _GEN_548; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_550 = 6'h26 == select_8 ? io_inData_38 : _GEN_549; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_551 = 6'h27 == select_8 ? io_inData_39 : _GEN_550; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_552 = 6'h28 == select_8 ? io_inData_40 : _GEN_551; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_553 = 6'h29 == select_8 ? io_inData_41 : _GEN_552; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_554 = 6'h2a == select_8 ? io_inData_42 : _GEN_553; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_555 = 6'h2b == select_8 ? io_inData_43 : _GEN_554; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_556 = 6'h2c == select_8 ? io_inData_44 : _GEN_555; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_557 = 6'h2d == select_8 ? io_inData_45 : _GEN_556; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_558 = 6'h2e == select_8 ? io_inData_46 : _GEN_557; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_559 = 6'h2f == select_8 ? io_inData_47 : _GEN_558; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_560 = 6'h30 == select_8 ? io_inData_48 : _GEN_559; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_561 = 6'h31 == select_8 ? io_inData_49 : _GEN_560; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_562 = 6'h32 == select_8 ? io_inData_50 : _GEN_561; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_563 = 6'h33 == select_8 ? io_inData_51 : _GEN_562; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_564 = 6'h34 == select_8 ? io_inData_52 : _GEN_563; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_565 = 6'h35 == select_8 ? io_inData_53 : _GEN_564; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_566 = 6'h36 == select_8 ? io_inData_54 : _GEN_565; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_567 = 6'h37 == select_8 ? io_inData_55 : _GEN_566; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_568 = 6'h38 == select_8 ? io_inData_56 : _GEN_567; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_569 = 6'h39 == select_8 ? io_inData_57 : _GEN_568; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_570 = 6'h3a == select_8 ? io_inData_58 : _GEN_569; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_571 = 6'h3b == select_8 ? io_inData_59 : _GEN_570; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_572 = 6'h3c == select_8 ? io_inData_60 : _GEN_571; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_573 = 6'h3d == select_8 ? io_inData_61 : _GEN_572; // @[Switch.scala 33:19:@2842.4]
  assign _GEN_574 = 6'h3e == select_8 ? io_inData_62 : _GEN_573; // @[Switch.scala 33:19:@2842.4]
  assign _T_21059 = {valid_8_7,valid_8_6,valid_8_5,valid_8_4,valid_8_3,valid_8_2,valid_8_1,valid_8_0}; // @[Switch.scala 34:32:@2849.4]
  assign _T_21067 = {valid_8_15,valid_8_14,valid_8_13,valid_8_12,valid_8_11,valid_8_10,valid_8_9,valid_8_8,_T_21059}; // @[Switch.scala 34:32:@2857.4]
  assign _T_21074 = {valid_8_23,valid_8_22,valid_8_21,valid_8_20,valid_8_19,valid_8_18,valid_8_17,valid_8_16}; // @[Switch.scala 34:32:@2864.4]
  assign _T_21083 = {valid_8_31,valid_8_30,valid_8_29,valid_8_28,valid_8_27,valid_8_26,valid_8_25,valid_8_24,_T_21074,_T_21067}; // @[Switch.scala 34:32:@2873.4]
  assign _T_21090 = {valid_8_39,valid_8_38,valid_8_37,valid_8_36,valid_8_35,valid_8_34,valid_8_33,valid_8_32}; // @[Switch.scala 34:32:@2880.4]
  assign _T_21098 = {valid_8_47,valid_8_46,valid_8_45,valid_8_44,valid_8_43,valid_8_42,valid_8_41,valid_8_40,_T_21090}; // @[Switch.scala 34:32:@2888.4]
  assign _T_21105 = {valid_8_55,valid_8_54,valid_8_53,valid_8_52,valid_8_51,valid_8_50,valid_8_49,valid_8_48}; // @[Switch.scala 34:32:@2895.4]
  assign _T_21114 = {valid_8_63,valid_8_62,valid_8_61,valid_8_60,valid_8_59,valid_8_58,valid_8_57,valid_8_56,_T_21105,_T_21098}; // @[Switch.scala 34:32:@2904.4]
  assign _T_21115 = {_T_21114,_T_21083}; // @[Switch.scala 34:32:@2905.4]
  assign _T_21119 = io_inAddr_0 == 6'h9; // @[Switch.scala 30:53:@2908.4]
  assign valid_9_0 = io_inValid_0 & _T_21119; // @[Switch.scala 30:36:@2909.4]
  assign _T_21122 = io_inAddr_1 == 6'h9; // @[Switch.scala 30:53:@2911.4]
  assign valid_9_1 = io_inValid_1 & _T_21122; // @[Switch.scala 30:36:@2912.4]
  assign _T_21125 = io_inAddr_2 == 6'h9; // @[Switch.scala 30:53:@2914.4]
  assign valid_9_2 = io_inValid_2 & _T_21125; // @[Switch.scala 30:36:@2915.4]
  assign _T_21128 = io_inAddr_3 == 6'h9; // @[Switch.scala 30:53:@2917.4]
  assign valid_9_3 = io_inValid_3 & _T_21128; // @[Switch.scala 30:36:@2918.4]
  assign _T_21131 = io_inAddr_4 == 6'h9; // @[Switch.scala 30:53:@2920.4]
  assign valid_9_4 = io_inValid_4 & _T_21131; // @[Switch.scala 30:36:@2921.4]
  assign _T_21134 = io_inAddr_5 == 6'h9; // @[Switch.scala 30:53:@2923.4]
  assign valid_9_5 = io_inValid_5 & _T_21134; // @[Switch.scala 30:36:@2924.4]
  assign _T_21137 = io_inAddr_6 == 6'h9; // @[Switch.scala 30:53:@2926.4]
  assign valid_9_6 = io_inValid_6 & _T_21137; // @[Switch.scala 30:36:@2927.4]
  assign _T_21140 = io_inAddr_7 == 6'h9; // @[Switch.scala 30:53:@2929.4]
  assign valid_9_7 = io_inValid_7 & _T_21140; // @[Switch.scala 30:36:@2930.4]
  assign _T_21143 = io_inAddr_8 == 6'h9; // @[Switch.scala 30:53:@2932.4]
  assign valid_9_8 = io_inValid_8 & _T_21143; // @[Switch.scala 30:36:@2933.4]
  assign _T_21146 = io_inAddr_9 == 6'h9; // @[Switch.scala 30:53:@2935.4]
  assign valid_9_9 = io_inValid_9 & _T_21146; // @[Switch.scala 30:36:@2936.4]
  assign _T_21149 = io_inAddr_10 == 6'h9; // @[Switch.scala 30:53:@2938.4]
  assign valid_9_10 = io_inValid_10 & _T_21149; // @[Switch.scala 30:36:@2939.4]
  assign _T_21152 = io_inAddr_11 == 6'h9; // @[Switch.scala 30:53:@2941.4]
  assign valid_9_11 = io_inValid_11 & _T_21152; // @[Switch.scala 30:36:@2942.4]
  assign _T_21155 = io_inAddr_12 == 6'h9; // @[Switch.scala 30:53:@2944.4]
  assign valid_9_12 = io_inValid_12 & _T_21155; // @[Switch.scala 30:36:@2945.4]
  assign _T_21158 = io_inAddr_13 == 6'h9; // @[Switch.scala 30:53:@2947.4]
  assign valid_9_13 = io_inValid_13 & _T_21158; // @[Switch.scala 30:36:@2948.4]
  assign _T_21161 = io_inAddr_14 == 6'h9; // @[Switch.scala 30:53:@2950.4]
  assign valid_9_14 = io_inValid_14 & _T_21161; // @[Switch.scala 30:36:@2951.4]
  assign _T_21164 = io_inAddr_15 == 6'h9; // @[Switch.scala 30:53:@2953.4]
  assign valid_9_15 = io_inValid_15 & _T_21164; // @[Switch.scala 30:36:@2954.4]
  assign _T_21167 = io_inAddr_16 == 6'h9; // @[Switch.scala 30:53:@2956.4]
  assign valid_9_16 = io_inValid_16 & _T_21167; // @[Switch.scala 30:36:@2957.4]
  assign _T_21170 = io_inAddr_17 == 6'h9; // @[Switch.scala 30:53:@2959.4]
  assign valid_9_17 = io_inValid_17 & _T_21170; // @[Switch.scala 30:36:@2960.4]
  assign _T_21173 = io_inAddr_18 == 6'h9; // @[Switch.scala 30:53:@2962.4]
  assign valid_9_18 = io_inValid_18 & _T_21173; // @[Switch.scala 30:36:@2963.4]
  assign _T_21176 = io_inAddr_19 == 6'h9; // @[Switch.scala 30:53:@2965.4]
  assign valid_9_19 = io_inValid_19 & _T_21176; // @[Switch.scala 30:36:@2966.4]
  assign _T_21179 = io_inAddr_20 == 6'h9; // @[Switch.scala 30:53:@2968.4]
  assign valid_9_20 = io_inValid_20 & _T_21179; // @[Switch.scala 30:36:@2969.4]
  assign _T_21182 = io_inAddr_21 == 6'h9; // @[Switch.scala 30:53:@2971.4]
  assign valid_9_21 = io_inValid_21 & _T_21182; // @[Switch.scala 30:36:@2972.4]
  assign _T_21185 = io_inAddr_22 == 6'h9; // @[Switch.scala 30:53:@2974.4]
  assign valid_9_22 = io_inValid_22 & _T_21185; // @[Switch.scala 30:36:@2975.4]
  assign _T_21188 = io_inAddr_23 == 6'h9; // @[Switch.scala 30:53:@2977.4]
  assign valid_9_23 = io_inValid_23 & _T_21188; // @[Switch.scala 30:36:@2978.4]
  assign _T_21191 = io_inAddr_24 == 6'h9; // @[Switch.scala 30:53:@2980.4]
  assign valid_9_24 = io_inValid_24 & _T_21191; // @[Switch.scala 30:36:@2981.4]
  assign _T_21194 = io_inAddr_25 == 6'h9; // @[Switch.scala 30:53:@2983.4]
  assign valid_9_25 = io_inValid_25 & _T_21194; // @[Switch.scala 30:36:@2984.4]
  assign _T_21197 = io_inAddr_26 == 6'h9; // @[Switch.scala 30:53:@2986.4]
  assign valid_9_26 = io_inValid_26 & _T_21197; // @[Switch.scala 30:36:@2987.4]
  assign _T_21200 = io_inAddr_27 == 6'h9; // @[Switch.scala 30:53:@2989.4]
  assign valid_9_27 = io_inValid_27 & _T_21200; // @[Switch.scala 30:36:@2990.4]
  assign _T_21203 = io_inAddr_28 == 6'h9; // @[Switch.scala 30:53:@2992.4]
  assign valid_9_28 = io_inValid_28 & _T_21203; // @[Switch.scala 30:36:@2993.4]
  assign _T_21206 = io_inAddr_29 == 6'h9; // @[Switch.scala 30:53:@2995.4]
  assign valid_9_29 = io_inValid_29 & _T_21206; // @[Switch.scala 30:36:@2996.4]
  assign _T_21209 = io_inAddr_30 == 6'h9; // @[Switch.scala 30:53:@2998.4]
  assign valid_9_30 = io_inValid_30 & _T_21209; // @[Switch.scala 30:36:@2999.4]
  assign _T_21212 = io_inAddr_31 == 6'h9; // @[Switch.scala 30:53:@3001.4]
  assign valid_9_31 = io_inValid_31 & _T_21212; // @[Switch.scala 30:36:@3002.4]
  assign _T_21215 = io_inAddr_32 == 6'h9; // @[Switch.scala 30:53:@3004.4]
  assign valid_9_32 = io_inValid_32 & _T_21215; // @[Switch.scala 30:36:@3005.4]
  assign _T_21218 = io_inAddr_33 == 6'h9; // @[Switch.scala 30:53:@3007.4]
  assign valid_9_33 = io_inValid_33 & _T_21218; // @[Switch.scala 30:36:@3008.4]
  assign _T_21221 = io_inAddr_34 == 6'h9; // @[Switch.scala 30:53:@3010.4]
  assign valid_9_34 = io_inValid_34 & _T_21221; // @[Switch.scala 30:36:@3011.4]
  assign _T_21224 = io_inAddr_35 == 6'h9; // @[Switch.scala 30:53:@3013.4]
  assign valid_9_35 = io_inValid_35 & _T_21224; // @[Switch.scala 30:36:@3014.4]
  assign _T_21227 = io_inAddr_36 == 6'h9; // @[Switch.scala 30:53:@3016.4]
  assign valid_9_36 = io_inValid_36 & _T_21227; // @[Switch.scala 30:36:@3017.4]
  assign _T_21230 = io_inAddr_37 == 6'h9; // @[Switch.scala 30:53:@3019.4]
  assign valid_9_37 = io_inValid_37 & _T_21230; // @[Switch.scala 30:36:@3020.4]
  assign _T_21233 = io_inAddr_38 == 6'h9; // @[Switch.scala 30:53:@3022.4]
  assign valid_9_38 = io_inValid_38 & _T_21233; // @[Switch.scala 30:36:@3023.4]
  assign _T_21236 = io_inAddr_39 == 6'h9; // @[Switch.scala 30:53:@3025.4]
  assign valid_9_39 = io_inValid_39 & _T_21236; // @[Switch.scala 30:36:@3026.4]
  assign _T_21239 = io_inAddr_40 == 6'h9; // @[Switch.scala 30:53:@3028.4]
  assign valid_9_40 = io_inValid_40 & _T_21239; // @[Switch.scala 30:36:@3029.4]
  assign _T_21242 = io_inAddr_41 == 6'h9; // @[Switch.scala 30:53:@3031.4]
  assign valid_9_41 = io_inValid_41 & _T_21242; // @[Switch.scala 30:36:@3032.4]
  assign _T_21245 = io_inAddr_42 == 6'h9; // @[Switch.scala 30:53:@3034.4]
  assign valid_9_42 = io_inValid_42 & _T_21245; // @[Switch.scala 30:36:@3035.4]
  assign _T_21248 = io_inAddr_43 == 6'h9; // @[Switch.scala 30:53:@3037.4]
  assign valid_9_43 = io_inValid_43 & _T_21248; // @[Switch.scala 30:36:@3038.4]
  assign _T_21251 = io_inAddr_44 == 6'h9; // @[Switch.scala 30:53:@3040.4]
  assign valid_9_44 = io_inValid_44 & _T_21251; // @[Switch.scala 30:36:@3041.4]
  assign _T_21254 = io_inAddr_45 == 6'h9; // @[Switch.scala 30:53:@3043.4]
  assign valid_9_45 = io_inValid_45 & _T_21254; // @[Switch.scala 30:36:@3044.4]
  assign _T_21257 = io_inAddr_46 == 6'h9; // @[Switch.scala 30:53:@3046.4]
  assign valid_9_46 = io_inValid_46 & _T_21257; // @[Switch.scala 30:36:@3047.4]
  assign _T_21260 = io_inAddr_47 == 6'h9; // @[Switch.scala 30:53:@3049.4]
  assign valid_9_47 = io_inValid_47 & _T_21260; // @[Switch.scala 30:36:@3050.4]
  assign _T_21263 = io_inAddr_48 == 6'h9; // @[Switch.scala 30:53:@3052.4]
  assign valid_9_48 = io_inValid_48 & _T_21263; // @[Switch.scala 30:36:@3053.4]
  assign _T_21266 = io_inAddr_49 == 6'h9; // @[Switch.scala 30:53:@3055.4]
  assign valid_9_49 = io_inValid_49 & _T_21266; // @[Switch.scala 30:36:@3056.4]
  assign _T_21269 = io_inAddr_50 == 6'h9; // @[Switch.scala 30:53:@3058.4]
  assign valid_9_50 = io_inValid_50 & _T_21269; // @[Switch.scala 30:36:@3059.4]
  assign _T_21272 = io_inAddr_51 == 6'h9; // @[Switch.scala 30:53:@3061.4]
  assign valid_9_51 = io_inValid_51 & _T_21272; // @[Switch.scala 30:36:@3062.4]
  assign _T_21275 = io_inAddr_52 == 6'h9; // @[Switch.scala 30:53:@3064.4]
  assign valid_9_52 = io_inValid_52 & _T_21275; // @[Switch.scala 30:36:@3065.4]
  assign _T_21278 = io_inAddr_53 == 6'h9; // @[Switch.scala 30:53:@3067.4]
  assign valid_9_53 = io_inValid_53 & _T_21278; // @[Switch.scala 30:36:@3068.4]
  assign _T_21281 = io_inAddr_54 == 6'h9; // @[Switch.scala 30:53:@3070.4]
  assign valid_9_54 = io_inValid_54 & _T_21281; // @[Switch.scala 30:36:@3071.4]
  assign _T_21284 = io_inAddr_55 == 6'h9; // @[Switch.scala 30:53:@3073.4]
  assign valid_9_55 = io_inValid_55 & _T_21284; // @[Switch.scala 30:36:@3074.4]
  assign _T_21287 = io_inAddr_56 == 6'h9; // @[Switch.scala 30:53:@3076.4]
  assign valid_9_56 = io_inValid_56 & _T_21287; // @[Switch.scala 30:36:@3077.4]
  assign _T_21290 = io_inAddr_57 == 6'h9; // @[Switch.scala 30:53:@3079.4]
  assign valid_9_57 = io_inValid_57 & _T_21290; // @[Switch.scala 30:36:@3080.4]
  assign _T_21293 = io_inAddr_58 == 6'h9; // @[Switch.scala 30:53:@3082.4]
  assign valid_9_58 = io_inValid_58 & _T_21293; // @[Switch.scala 30:36:@3083.4]
  assign _T_21296 = io_inAddr_59 == 6'h9; // @[Switch.scala 30:53:@3085.4]
  assign valid_9_59 = io_inValid_59 & _T_21296; // @[Switch.scala 30:36:@3086.4]
  assign _T_21299 = io_inAddr_60 == 6'h9; // @[Switch.scala 30:53:@3088.4]
  assign valid_9_60 = io_inValid_60 & _T_21299; // @[Switch.scala 30:36:@3089.4]
  assign _T_21302 = io_inAddr_61 == 6'h9; // @[Switch.scala 30:53:@3091.4]
  assign valid_9_61 = io_inValid_61 & _T_21302; // @[Switch.scala 30:36:@3092.4]
  assign _T_21305 = io_inAddr_62 == 6'h9; // @[Switch.scala 30:53:@3094.4]
  assign valid_9_62 = io_inValid_62 & _T_21305; // @[Switch.scala 30:36:@3095.4]
  assign _T_21308 = io_inAddr_63 == 6'h9; // @[Switch.scala 30:53:@3097.4]
  assign valid_9_63 = io_inValid_63 & _T_21308; // @[Switch.scala 30:36:@3098.4]
  assign _T_21374 = valid_9_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@3100.4]
  assign _T_21375 = valid_9_61 ? 6'h3d : _T_21374; // @[Mux.scala 31:69:@3101.4]
  assign _T_21376 = valid_9_60 ? 6'h3c : _T_21375; // @[Mux.scala 31:69:@3102.4]
  assign _T_21377 = valid_9_59 ? 6'h3b : _T_21376; // @[Mux.scala 31:69:@3103.4]
  assign _T_21378 = valid_9_58 ? 6'h3a : _T_21377; // @[Mux.scala 31:69:@3104.4]
  assign _T_21379 = valid_9_57 ? 6'h39 : _T_21378; // @[Mux.scala 31:69:@3105.4]
  assign _T_21380 = valid_9_56 ? 6'h38 : _T_21379; // @[Mux.scala 31:69:@3106.4]
  assign _T_21381 = valid_9_55 ? 6'h37 : _T_21380; // @[Mux.scala 31:69:@3107.4]
  assign _T_21382 = valid_9_54 ? 6'h36 : _T_21381; // @[Mux.scala 31:69:@3108.4]
  assign _T_21383 = valid_9_53 ? 6'h35 : _T_21382; // @[Mux.scala 31:69:@3109.4]
  assign _T_21384 = valid_9_52 ? 6'h34 : _T_21383; // @[Mux.scala 31:69:@3110.4]
  assign _T_21385 = valid_9_51 ? 6'h33 : _T_21384; // @[Mux.scala 31:69:@3111.4]
  assign _T_21386 = valid_9_50 ? 6'h32 : _T_21385; // @[Mux.scala 31:69:@3112.4]
  assign _T_21387 = valid_9_49 ? 6'h31 : _T_21386; // @[Mux.scala 31:69:@3113.4]
  assign _T_21388 = valid_9_48 ? 6'h30 : _T_21387; // @[Mux.scala 31:69:@3114.4]
  assign _T_21389 = valid_9_47 ? 6'h2f : _T_21388; // @[Mux.scala 31:69:@3115.4]
  assign _T_21390 = valid_9_46 ? 6'h2e : _T_21389; // @[Mux.scala 31:69:@3116.4]
  assign _T_21391 = valid_9_45 ? 6'h2d : _T_21390; // @[Mux.scala 31:69:@3117.4]
  assign _T_21392 = valid_9_44 ? 6'h2c : _T_21391; // @[Mux.scala 31:69:@3118.4]
  assign _T_21393 = valid_9_43 ? 6'h2b : _T_21392; // @[Mux.scala 31:69:@3119.4]
  assign _T_21394 = valid_9_42 ? 6'h2a : _T_21393; // @[Mux.scala 31:69:@3120.4]
  assign _T_21395 = valid_9_41 ? 6'h29 : _T_21394; // @[Mux.scala 31:69:@3121.4]
  assign _T_21396 = valid_9_40 ? 6'h28 : _T_21395; // @[Mux.scala 31:69:@3122.4]
  assign _T_21397 = valid_9_39 ? 6'h27 : _T_21396; // @[Mux.scala 31:69:@3123.4]
  assign _T_21398 = valid_9_38 ? 6'h26 : _T_21397; // @[Mux.scala 31:69:@3124.4]
  assign _T_21399 = valid_9_37 ? 6'h25 : _T_21398; // @[Mux.scala 31:69:@3125.4]
  assign _T_21400 = valid_9_36 ? 6'h24 : _T_21399; // @[Mux.scala 31:69:@3126.4]
  assign _T_21401 = valid_9_35 ? 6'h23 : _T_21400; // @[Mux.scala 31:69:@3127.4]
  assign _T_21402 = valid_9_34 ? 6'h22 : _T_21401; // @[Mux.scala 31:69:@3128.4]
  assign _T_21403 = valid_9_33 ? 6'h21 : _T_21402; // @[Mux.scala 31:69:@3129.4]
  assign _T_21404 = valid_9_32 ? 6'h20 : _T_21403; // @[Mux.scala 31:69:@3130.4]
  assign _T_21405 = valid_9_31 ? 6'h1f : _T_21404; // @[Mux.scala 31:69:@3131.4]
  assign _T_21406 = valid_9_30 ? 6'h1e : _T_21405; // @[Mux.scala 31:69:@3132.4]
  assign _T_21407 = valid_9_29 ? 6'h1d : _T_21406; // @[Mux.scala 31:69:@3133.4]
  assign _T_21408 = valid_9_28 ? 6'h1c : _T_21407; // @[Mux.scala 31:69:@3134.4]
  assign _T_21409 = valid_9_27 ? 6'h1b : _T_21408; // @[Mux.scala 31:69:@3135.4]
  assign _T_21410 = valid_9_26 ? 6'h1a : _T_21409; // @[Mux.scala 31:69:@3136.4]
  assign _T_21411 = valid_9_25 ? 6'h19 : _T_21410; // @[Mux.scala 31:69:@3137.4]
  assign _T_21412 = valid_9_24 ? 6'h18 : _T_21411; // @[Mux.scala 31:69:@3138.4]
  assign _T_21413 = valid_9_23 ? 6'h17 : _T_21412; // @[Mux.scala 31:69:@3139.4]
  assign _T_21414 = valid_9_22 ? 6'h16 : _T_21413; // @[Mux.scala 31:69:@3140.4]
  assign _T_21415 = valid_9_21 ? 6'h15 : _T_21414; // @[Mux.scala 31:69:@3141.4]
  assign _T_21416 = valid_9_20 ? 6'h14 : _T_21415; // @[Mux.scala 31:69:@3142.4]
  assign _T_21417 = valid_9_19 ? 6'h13 : _T_21416; // @[Mux.scala 31:69:@3143.4]
  assign _T_21418 = valid_9_18 ? 6'h12 : _T_21417; // @[Mux.scala 31:69:@3144.4]
  assign _T_21419 = valid_9_17 ? 6'h11 : _T_21418; // @[Mux.scala 31:69:@3145.4]
  assign _T_21420 = valid_9_16 ? 6'h10 : _T_21419; // @[Mux.scala 31:69:@3146.4]
  assign _T_21421 = valid_9_15 ? 6'hf : _T_21420; // @[Mux.scala 31:69:@3147.4]
  assign _T_21422 = valid_9_14 ? 6'he : _T_21421; // @[Mux.scala 31:69:@3148.4]
  assign _T_21423 = valid_9_13 ? 6'hd : _T_21422; // @[Mux.scala 31:69:@3149.4]
  assign _T_21424 = valid_9_12 ? 6'hc : _T_21423; // @[Mux.scala 31:69:@3150.4]
  assign _T_21425 = valid_9_11 ? 6'hb : _T_21424; // @[Mux.scala 31:69:@3151.4]
  assign _T_21426 = valid_9_10 ? 6'ha : _T_21425; // @[Mux.scala 31:69:@3152.4]
  assign _T_21427 = valid_9_9 ? 6'h9 : _T_21426; // @[Mux.scala 31:69:@3153.4]
  assign _T_21428 = valid_9_8 ? 6'h8 : _T_21427; // @[Mux.scala 31:69:@3154.4]
  assign _T_21429 = valid_9_7 ? 6'h7 : _T_21428; // @[Mux.scala 31:69:@3155.4]
  assign _T_21430 = valid_9_6 ? 6'h6 : _T_21429; // @[Mux.scala 31:69:@3156.4]
  assign _T_21431 = valid_9_5 ? 6'h5 : _T_21430; // @[Mux.scala 31:69:@3157.4]
  assign _T_21432 = valid_9_4 ? 6'h4 : _T_21431; // @[Mux.scala 31:69:@3158.4]
  assign _T_21433 = valid_9_3 ? 6'h3 : _T_21432; // @[Mux.scala 31:69:@3159.4]
  assign _T_21434 = valid_9_2 ? 6'h2 : _T_21433; // @[Mux.scala 31:69:@3160.4]
  assign _T_21435 = valid_9_1 ? 6'h1 : _T_21434; // @[Mux.scala 31:69:@3161.4]
  assign select_9 = valid_9_0 ? 6'h0 : _T_21435; // @[Mux.scala 31:69:@3162.4]
  assign _GEN_577 = 6'h1 == select_9 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_578 = 6'h2 == select_9 ? io_inData_2 : _GEN_577; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_579 = 6'h3 == select_9 ? io_inData_3 : _GEN_578; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_580 = 6'h4 == select_9 ? io_inData_4 : _GEN_579; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_581 = 6'h5 == select_9 ? io_inData_5 : _GEN_580; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_582 = 6'h6 == select_9 ? io_inData_6 : _GEN_581; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_583 = 6'h7 == select_9 ? io_inData_7 : _GEN_582; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_584 = 6'h8 == select_9 ? io_inData_8 : _GEN_583; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_585 = 6'h9 == select_9 ? io_inData_9 : _GEN_584; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_586 = 6'ha == select_9 ? io_inData_10 : _GEN_585; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_587 = 6'hb == select_9 ? io_inData_11 : _GEN_586; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_588 = 6'hc == select_9 ? io_inData_12 : _GEN_587; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_589 = 6'hd == select_9 ? io_inData_13 : _GEN_588; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_590 = 6'he == select_9 ? io_inData_14 : _GEN_589; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_591 = 6'hf == select_9 ? io_inData_15 : _GEN_590; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_592 = 6'h10 == select_9 ? io_inData_16 : _GEN_591; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_593 = 6'h11 == select_9 ? io_inData_17 : _GEN_592; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_594 = 6'h12 == select_9 ? io_inData_18 : _GEN_593; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_595 = 6'h13 == select_9 ? io_inData_19 : _GEN_594; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_596 = 6'h14 == select_9 ? io_inData_20 : _GEN_595; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_597 = 6'h15 == select_9 ? io_inData_21 : _GEN_596; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_598 = 6'h16 == select_9 ? io_inData_22 : _GEN_597; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_599 = 6'h17 == select_9 ? io_inData_23 : _GEN_598; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_600 = 6'h18 == select_9 ? io_inData_24 : _GEN_599; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_601 = 6'h19 == select_9 ? io_inData_25 : _GEN_600; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_602 = 6'h1a == select_9 ? io_inData_26 : _GEN_601; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_603 = 6'h1b == select_9 ? io_inData_27 : _GEN_602; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_604 = 6'h1c == select_9 ? io_inData_28 : _GEN_603; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_605 = 6'h1d == select_9 ? io_inData_29 : _GEN_604; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_606 = 6'h1e == select_9 ? io_inData_30 : _GEN_605; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_607 = 6'h1f == select_9 ? io_inData_31 : _GEN_606; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_608 = 6'h20 == select_9 ? io_inData_32 : _GEN_607; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_609 = 6'h21 == select_9 ? io_inData_33 : _GEN_608; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_610 = 6'h22 == select_9 ? io_inData_34 : _GEN_609; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_611 = 6'h23 == select_9 ? io_inData_35 : _GEN_610; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_612 = 6'h24 == select_9 ? io_inData_36 : _GEN_611; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_613 = 6'h25 == select_9 ? io_inData_37 : _GEN_612; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_614 = 6'h26 == select_9 ? io_inData_38 : _GEN_613; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_615 = 6'h27 == select_9 ? io_inData_39 : _GEN_614; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_616 = 6'h28 == select_9 ? io_inData_40 : _GEN_615; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_617 = 6'h29 == select_9 ? io_inData_41 : _GEN_616; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_618 = 6'h2a == select_9 ? io_inData_42 : _GEN_617; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_619 = 6'h2b == select_9 ? io_inData_43 : _GEN_618; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_620 = 6'h2c == select_9 ? io_inData_44 : _GEN_619; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_621 = 6'h2d == select_9 ? io_inData_45 : _GEN_620; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_622 = 6'h2e == select_9 ? io_inData_46 : _GEN_621; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_623 = 6'h2f == select_9 ? io_inData_47 : _GEN_622; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_624 = 6'h30 == select_9 ? io_inData_48 : _GEN_623; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_625 = 6'h31 == select_9 ? io_inData_49 : _GEN_624; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_626 = 6'h32 == select_9 ? io_inData_50 : _GEN_625; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_627 = 6'h33 == select_9 ? io_inData_51 : _GEN_626; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_628 = 6'h34 == select_9 ? io_inData_52 : _GEN_627; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_629 = 6'h35 == select_9 ? io_inData_53 : _GEN_628; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_630 = 6'h36 == select_9 ? io_inData_54 : _GEN_629; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_631 = 6'h37 == select_9 ? io_inData_55 : _GEN_630; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_632 = 6'h38 == select_9 ? io_inData_56 : _GEN_631; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_633 = 6'h39 == select_9 ? io_inData_57 : _GEN_632; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_634 = 6'h3a == select_9 ? io_inData_58 : _GEN_633; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_635 = 6'h3b == select_9 ? io_inData_59 : _GEN_634; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_636 = 6'h3c == select_9 ? io_inData_60 : _GEN_635; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_637 = 6'h3d == select_9 ? io_inData_61 : _GEN_636; // @[Switch.scala 33:19:@3164.4]
  assign _GEN_638 = 6'h3e == select_9 ? io_inData_62 : _GEN_637; // @[Switch.scala 33:19:@3164.4]
  assign _T_21444 = {valid_9_7,valid_9_6,valid_9_5,valid_9_4,valid_9_3,valid_9_2,valid_9_1,valid_9_0}; // @[Switch.scala 34:32:@3171.4]
  assign _T_21452 = {valid_9_15,valid_9_14,valid_9_13,valid_9_12,valid_9_11,valid_9_10,valid_9_9,valid_9_8,_T_21444}; // @[Switch.scala 34:32:@3179.4]
  assign _T_21459 = {valid_9_23,valid_9_22,valid_9_21,valid_9_20,valid_9_19,valid_9_18,valid_9_17,valid_9_16}; // @[Switch.scala 34:32:@3186.4]
  assign _T_21468 = {valid_9_31,valid_9_30,valid_9_29,valid_9_28,valid_9_27,valid_9_26,valid_9_25,valid_9_24,_T_21459,_T_21452}; // @[Switch.scala 34:32:@3195.4]
  assign _T_21475 = {valid_9_39,valid_9_38,valid_9_37,valid_9_36,valid_9_35,valid_9_34,valid_9_33,valid_9_32}; // @[Switch.scala 34:32:@3202.4]
  assign _T_21483 = {valid_9_47,valid_9_46,valid_9_45,valid_9_44,valid_9_43,valid_9_42,valid_9_41,valid_9_40,_T_21475}; // @[Switch.scala 34:32:@3210.4]
  assign _T_21490 = {valid_9_55,valid_9_54,valid_9_53,valid_9_52,valid_9_51,valid_9_50,valid_9_49,valid_9_48}; // @[Switch.scala 34:32:@3217.4]
  assign _T_21499 = {valid_9_63,valid_9_62,valid_9_61,valid_9_60,valid_9_59,valid_9_58,valid_9_57,valid_9_56,_T_21490,_T_21483}; // @[Switch.scala 34:32:@3226.4]
  assign _T_21500 = {_T_21499,_T_21468}; // @[Switch.scala 34:32:@3227.4]
  assign _T_21504 = io_inAddr_0 == 6'ha; // @[Switch.scala 30:53:@3230.4]
  assign valid_10_0 = io_inValid_0 & _T_21504; // @[Switch.scala 30:36:@3231.4]
  assign _T_21507 = io_inAddr_1 == 6'ha; // @[Switch.scala 30:53:@3233.4]
  assign valid_10_1 = io_inValid_1 & _T_21507; // @[Switch.scala 30:36:@3234.4]
  assign _T_21510 = io_inAddr_2 == 6'ha; // @[Switch.scala 30:53:@3236.4]
  assign valid_10_2 = io_inValid_2 & _T_21510; // @[Switch.scala 30:36:@3237.4]
  assign _T_21513 = io_inAddr_3 == 6'ha; // @[Switch.scala 30:53:@3239.4]
  assign valid_10_3 = io_inValid_3 & _T_21513; // @[Switch.scala 30:36:@3240.4]
  assign _T_21516 = io_inAddr_4 == 6'ha; // @[Switch.scala 30:53:@3242.4]
  assign valid_10_4 = io_inValid_4 & _T_21516; // @[Switch.scala 30:36:@3243.4]
  assign _T_21519 = io_inAddr_5 == 6'ha; // @[Switch.scala 30:53:@3245.4]
  assign valid_10_5 = io_inValid_5 & _T_21519; // @[Switch.scala 30:36:@3246.4]
  assign _T_21522 = io_inAddr_6 == 6'ha; // @[Switch.scala 30:53:@3248.4]
  assign valid_10_6 = io_inValid_6 & _T_21522; // @[Switch.scala 30:36:@3249.4]
  assign _T_21525 = io_inAddr_7 == 6'ha; // @[Switch.scala 30:53:@3251.4]
  assign valid_10_7 = io_inValid_7 & _T_21525; // @[Switch.scala 30:36:@3252.4]
  assign _T_21528 = io_inAddr_8 == 6'ha; // @[Switch.scala 30:53:@3254.4]
  assign valid_10_8 = io_inValid_8 & _T_21528; // @[Switch.scala 30:36:@3255.4]
  assign _T_21531 = io_inAddr_9 == 6'ha; // @[Switch.scala 30:53:@3257.4]
  assign valid_10_9 = io_inValid_9 & _T_21531; // @[Switch.scala 30:36:@3258.4]
  assign _T_21534 = io_inAddr_10 == 6'ha; // @[Switch.scala 30:53:@3260.4]
  assign valid_10_10 = io_inValid_10 & _T_21534; // @[Switch.scala 30:36:@3261.4]
  assign _T_21537 = io_inAddr_11 == 6'ha; // @[Switch.scala 30:53:@3263.4]
  assign valid_10_11 = io_inValid_11 & _T_21537; // @[Switch.scala 30:36:@3264.4]
  assign _T_21540 = io_inAddr_12 == 6'ha; // @[Switch.scala 30:53:@3266.4]
  assign valid_10_12 = io_inValid_12 & _T_21540; // @[Switch.scala 30:36:@3267.4]
  assign _T_21543 = io_inAddr_13 == 6'ha; // @[Switch.scala 30:53:@3269.4]
  assign valid_10_13 = io_inValid_13 & _T_21543; // @[Switch.scala 30:36:@3270.4]
  assign _T_21546 = io_inAddr_14 == 6'ha; // @[Switch.scala 30:53:@3272.4]
  assign valid_10_14 = io_inValid_14 & _T_21546; // @[Switch.scala 30:36:@3273.4]
  assign _T_21549 = io_inAddr_15 == 6'ha; // @[Switch.scala 30:53:@3275.4]
  assign valid_10_15 = io_inValid_15 & _T_21549; // @[Switch.scala 30:36:@3276.4]
  assign _T_21552 = io_inAddr_16 == 6'ha; // @[Switch.scala 30:53:@3278.4]
  assign valid_10_16 = io_inValid_16 & _T_21552; // @[Switch.scala 30:36:@3279.4]
  assign _T_21555 = io_inAddr_17 == 6'ha; // @[Switch.scala 30:53:@3281.4]
  assign valid_10_17 = io_inValid_17 & _T_21555; // @[Switch.scala 30:36:@3282.4]
  assign _T_21558 = io_inAddr_18 == 6'ha; // @[Switch.scala 30:53:@3284.4]
  assign valid_10_18 = io_inValid_18 & _T_21558; // @[Switch.scala 30:36:@3285.4]
  assign _T_21561 = io_inAddr_19 == 6'ha; // @[Switch.scala 30:53:@3287.4]
  assign valid_10_19 = io_inValid_19 & _T_21561; // @[Switch.scala 30:36:@3288.4]
  assign _T_21564 = io_inAddr_20 == 6'ha; // @[Switch.scala 30:53:@3290.4]
  assign valid_10_20 = io_inValid_20 & _T_21564; // @[Switch.scala 30:36:@3291.4]
  assign _T_21567 = io_inAddr_21 == 6'ha; // @[Switch.scala 30:53:@3293.4]
  assign valid_10_21 = io_inValid_21 & _T_21567; // @[Switch.scala 30:36:@3294.4]
  assign _T_21570 = io_inAddr_22 == 6'ha; // @[Switch.scala 30:53:@3296.4]
  assign valid_10_22 = io_inValid_22 & _T_21570; // @[Switch.scala 30:36:@3297.4]
  assign _T_21573 = io_inAddr_23 == 6'ha; // @[Switch.scala 30:53:@3299.4]
  assign valid_10_23 = io_inValid_23 & _T_21573; // @[Switch.scala 30:36:@3300.4]
  assign _T_21576 = io_inAddr_24 == 6'ha; // @[Switch.scala 30:53:@3302.4]
  assign valid_10_24 = io_inValid_24 & _T_21576; // @[Switch.scala 30:36:@3303.4]
  assign _T_21579 = io_inAddr_25 == 6'ha; // @[Switch.scala 30:53:@3305.4]
  assign valid_10_25 = io_inValid_25 & _T_21579; // @[Switch.scala 30:36:@3306.4]
  assign _T_21582 = io_inAddr_26 == 6'ha; // @[Switch.scala 30:53:@3308.4]
  assign valid_10_26 = io_inValid_26 & _T_21582; // @[Switch.scala 30:36:@3309.4]
  assign _T_21585 = io_inAddr_27 == 6'ha; // @[Switch.scala 30:53:@3311.4]
  assign valid_10_27 = io_inValid_27 & _T_21585; // @[Switch.scala 30:36:@3312.4]
  assign _T_21588 = io_inAddr_28 == 6'ha; // @[Switch.scala 30:53:@3314.4]
  assign valid_10_28 = io_inValid_28 & _T_21588; // @[Switch.scala 30:36:@3315.4]
  assign _T_21591 = io_inAddr_29 == 6'ha; // @[Switch.scala 30:53:@3317.4]
  assign valid_10_29 = io_inValid_29 & _T_21591; // @[Switch.scala 30:36:@3318.4]
  assign _T_21594 = io_inAddr_30 == 6'ha; // @[Switch.scala 30:53:@3320.4]
  assign valid_10_30 = io_inValid_30 & _T_21594; // @[Switch.scala 30:36:@3321.4]
  assign _T_21597 = io_inAddr_31 == 6'ha; // @[Switch.scala 30:53:@3323.4]
  assign valid_10_31 = io_inValid_31 & _T_21597; // @[Switch.scala 30:36:@3324.4]
  assign _T_21600 = io_inAddr_32 == 6'ha; // @[Switch.scala 30:53:@3326.4]
  assign valid_10_32 = io_inValid_32 & _T_21600; // @[Switch.scala 30:36:@3327.4]
  assign _T_21603 = io_inAddr_33 == 6'ha; // @[Switch.scala 30:53:@3329.4]
  assign valid_10_33 = io_inValid_33 & _T_21603; // @[Switch.scala 30:36:@3330.4]
  assign _T_21606 = io_inAddr_34 == 6'ha; // @[Switch.scala 30:53:@3332.4]
  assign valid_10_34 = io_inValid_34 & _T_21606; // @[Switch.scala 30:36:@3333.4]
  assign _T_21609 = io_inAddr_35 == 6'ha; // @[Switch.scala 30:53:@3335.4]
  assign valid_10_35 = io_inValid_35 & _T_21609; // @[Switch.scala 30:36:@3336.4]
  assign _T_21612 = io_inAddr_36 == 6'ha; // @[Switch.scala 30:53:@3338.4]
  assign valid_10_36 = io_inValid_36 & _T_21612; // @[Switch.scala 30:36:@3339.4]
  assign _T_21615 = io_inAddr_37 == 6'ha; // @[Switch.scala 30:53:@3341.4]
  assign valid_10_37 = io_inValid_37 & _T_21615; // @[Switch.scala 30:36:@3342.4]
  assign _T_21618 = io_inAddr_38 == 6'ha; // @[Switch.scala 30:53:@3344.4]
  assign valid_10_38 = io_inValid_38 & _T_21618; // @[Switch.scala 30:36:@3345.4]
  assign _T_21621 = io_inAddr_39 == 6'ha; // @[Switch.scala 30:53:@3347.4]
  assign valid_10_39 = io_inValid_39 & _T_21621; // @[Switch.scala 30:36:@3348.4]
  assign _T_21624 = io_inAddr_40 == 6'ha; // @[Switch.scala 30:53:@3350.4]
  assign valid_10_40 = io_inValid_40 & _T_21624; // @[Switch.scala 30:36:@3351.4]
  assign _T_21627 = io_inAddr_41 == 6'ha; // @[Switch.scala 30:53:@3353.4]
  assign valid_10_41 = io_inValid_41 & _T_21627; // @[Switch.scala 30:36:@3354.4]
  assign _T_21630 = io_inAddr_42 == 6'ha; // @[Switch.scala 30:53:@3356.4]
  assign valid_10_42 = io_inValid_42 & _T_21630; // @[Switch.scala 30:36:@3357.4]
  assign _T_21633 = io_inAddr_43 == 6'ha; // @[Switch.scala 30:53:@3359.4]
  assign valid_10_43 = io_inValid_43 & _T_21633; // @[Switch.scala 30:36:@3360.4]
  assign _T_21636 = io_inAddr_44 == 6'ha; // @[Switch.scala 30:53:@3362.4]
  assign valid_10_44 = io_inValid_44 & _T_21636; // @[Switch.scala 30:36:@3363.4]
  assign _T_21639 = io_inAddr_45 == 6'ha; // @[Switch.scala 30:53:@3365.4]
  assign valid_10_45 = io_inValid_45 & _T_21639; // @[Switch.scala 30:36:@3366.4]
  assign _T_21642 = io_inAddr_46 == 6'ha; // @[Switch.scala 30:53:@3368.4]
  assign valid_10_46 = io_inValid_46 & _T_21642; // @[Switch.scala 30:36:@3369.4]
  assign _T_21645 = io_inAddr_47 == 6'ha; // @[Switch.scala 30:53:@3371.4]
  assign valid_10_47 = io_inValid_47 & _T_21645; // @[Switch.scala 30:36:@3372.4]
  assign _T_21648 = io_inAddr_48 == 6'ha; // @[Switch.scala 30:53:@3374.4]
  assign valid_10_48 = io_inValid_48 & _T_21648; // @[Switch.scala 30:36:@3375.4]
  assign _T_21651 = io_inAddr_49 == 6'ha; // @[Switch.scala 30:53:@3377.4]
  assign valid_10_49 = io_inValid_49 & _T_21651; // @[Switch.scala 30:36:@3378.4]
  assign _T_21654 = io_inAddr_50 == 6'ha; // @[Switch.scala 30:53:@3380.4]
  assign valid_10_50 = io_inValid_50 & _T_21654; // @[Switch.scala 30:36:@3381.4]
  assign _T_21657 = io_inAddr_51 == 6'ha; // @[Switch.scala 30:53:@3383.4]
  assign valid_10_51 = io_inValid_51 & _T_21657; // @[Switch.scala 30:36:@3384.4]
  assign _T_21660 = io_inAddr_52 == 6'ha; // @[Switch.scala 30:53:@3386.4]
  assign valid_10_52 = io_inValid_52 & _T_21660; // @[Switch.scala 30:36:@3387.4]
  assign _T_21663 = io_inAddr_53 == 6'ha; // @[Switch.scala 30:53:@3389.4]
  assign valid_10_53 = io_inValid_53 & _T_21663; // @[Switch.scala 30:36:@3390.4]
  assign _T_21666 = io_inAddr_54 == 6'ha; // @[Switch.scala 30:53:@3392.4]
  assign valid_10_54 = io_inValid_54 & _T_21666; // @[Switch.scala 30:36:@3393.4]
  assign _T_21669 = io_inAddr_55 == 6'ha; // @[Switch.scala 30:53:@3395.4]
  assign valid_10_55 = io_inValid_55 & _T_21669; // @[Switch.scala 30:36:@3396.4]
  assign _T_21672 = io_inAddr_56 == 6'ha; // @[Switch.scala 30:53:@3398.4]
  assign valid_10_56 = io_inValid_56 & _T_21672; // @[Switch.scala 30:36:@3399.4]
  assign _T_21675 = io_inAddr_57 == 6'ha; // @[Switch.scala 30:53:@3401.4]
  assign valid_10_57 = io_inValid_57 & _T_21675; // @[Switch.scala 30:36:@3402.4]
  assign _T_21678 = io_inAddr_58 == 6'ha; // @[Switch.scala 30:53:@3404.4]
  assign valid_10_58 = io_inValid_58 & _T_21678; // @[Switch.scala 30:36:@3405.4]
  assign _T_21681 = io_inAddr_59 == 6'ha; // @[Switch.scala 30:53:@3407.4]
  assign valid_10_59 = io_inValid_59 & _T_21681; // @[Switch.scala 30:36:@3408.4]
  assign _T_21684 = io_inAddr_60 == 6'ha; // @[Switch.scala 30:53:@3410.4]
  assign valid_10_60 = io_inValid_60 & _T_21684; // @[Switch.scala 30:36:@3411.4]
  assign _T_21687 = io_inAddr_61 == 6'ha; // @[Switch.scala 30:53:@3413.4]
  assign valid_10_61 = io_inValid_61 & _T_21687; // @[Switch.scala 30:36:@3414.4]
  assign _T_21690 = io_inAddr_62 == 6'ha; // @[Switch.scala 30:53:@3416.4]
  assign valid_10_62 = io_inValid_62 & _T_21690; // @[Switch.scala 30:36:@3417.4]
  assign _T_21693 = io_inAddr_63 == 6'ha; // @[Switch.scala 30:53:@3419.4]
  assign valid_10_63 = io_inValid_63 & _T_21693; // @[Switch.scala 30:36:@3420.4]
  assign _T_21759 = valid_10_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@3422.4]
  assign _T_21760 = valid_10_61 ? 6'h3d : _T_21759; // @[Mux.scala 31:69:@3423.4]
  assign _T_21761 = valid_10_60 ? 6'h3c : _T_21760; // @[Mux.scala 31:69:@3424.4]
  assign _T_21762 = valid_10_59 ? 6'h3b : _T_21761; // @[Mux.scala 31:69:@3425.4]
  assign _T_21763 = valid_10_58 ? 6'h3a : _T_21762; // @[Mux.scala 31:69:@3426.4]
  assign _T_21764 = valid_10_57 ? 6'h39 : _T_21763; // @[Mux.scala 31:69:@3427.4]
  assign _T_21765 = valid_10_56 ? 6'h38 : _T_21764; // @[Mux.scala 31:69:@3428.4]
  assign _T_21766 = valid_10_55 ? 6'h37 : _T_21765; // @[Mux.scala 31:69:@3429.4]
  assign _T_21767 = valid_10_54 ? 6'h36 : _T_21766; // @[Mux.scala 31:69:@3430.4]
  assign _T_21768 = valid_10_53 ? 6'h35 : _T_21767; // @[Mux.scala 31:69:@3431.4]
  assign _T_21769 = valid_10_52 ? 6'h34 : _T_21768; // @[Mux.scala 31:69:@3432.4]
  assign _T_21770 = valid_10_51 ? 6'h33 : _T_21769; // @[Mux.scala 31:69:@3433.4]
  assign _T_21771 = valid_10_50 ? 6'h32 : _T_21770; // @[Mux.scala 31:69:@3434.4]
  assign _T_21772 = valid_10_49 ? 6'h31 : _T_21771; // @[Mux.scala 31:69:@3435.4]
  assign _T_21773 = valid_10_48 ? 6'h30 : _T_21772; // @[Mux.scala 31:69:@3436.4]
  assign _T_21774 = valid_10_47 ? 6'h2f : _T_21773; // @[Mux.scala 31:69:@3437.4]
  assign _T_21775 = valid_10_46 ? 6'h2e : _T_21774; // @[Mux.scala 31:69:@3438.4]
  assign _T_21776 = valid_10_45 ? 6'h2d : _T_21775; // @[Mux.scala 31:69:@3439.4]
  assign _T_21777 = valid_10_44 ? 6'h2c : _T_21776; // @[Mux.scala 31:69:@3440.4]
  assign _T_21778 = valid_10_43 ? 6'h2b : _T_21777; // @[Mux.scala 31:69:@3441.4]
  assign _T_21779 = valid_10_42 ? 6'h2a : _T_21778; // @[Mux.scala 31:69:@3442.4]
  assign _T_21780 = valid_10_41 ? 6'h29 : _T_21779; // @[Mux.scala 31:69:@3443.4]
  assign _T_21781 = valid_10_40 ? 6'h28 : _T_21780; // @[Mux.scala 31:69:@3444.4]
  assign _T_21782 = valid_10_39 ? 6'h27 : _T_21781; // @[Mux.scala 31:69:@3445.4]
  assign _T_21783 = valid_10_38 ? 6'h26 : _T_21782; // @[Mux.scala 31:69:@3446.4]
  assign _T_21784 = valid_10_37 ? 6'h25 : _T_21783; // @[Mux.scala 31:69:@3447.4]
  assign _T_21785 = valid_10_36 ? 6'h24 : _T_21784; // @[Mux.scala 31:69:@3448.4]
  assign _T_21786 = valid_10_35 ? 6'h23 : _T_21785; // @[Mux.scala 31:69:@3449.4]
  assign _T_21787 = valid_10_34 ? 6'h22 : _T_21786; // @[Mux.scala 31:69:@3450.4]
  assign _T_21788 = valid_10_33 ? 6'h21 : _T_21787; // @[Mux.scala 31:69:@3451.4]
  assign _T_21789 = valid_10_32 ? 6'h20 : _T_21788; // @[Mux.scala 31:69:@3452.4]
  assign _T_21790 = valid_10_31 ? 6'h1f : _T_21789; // @[Mux.scala 31:69:@3453.4]
  assign _T_21791 = valid_10_30 ? 6'h1e : _T_21790; // @[Mux.scala 31:69:@3454.4]
  assign _T_21792 = valid_10_29 ? 6'h1d : _T_21791; // @[Mux.scala 31:69:@3455.4]
  assign _T_21793 = valid_10_28 ? 6'h1c : _T_21792; // @[Mux.scala 31:69:@3456.4]
  assign _T_21794 = valid_10_27 ? 6'h1b : _T_21793; // @[Mux.scala 31:69:@3457.4]
  assign _T_21795 = valid_10_26 ? 6'h1a : _T_21794; // @[Mux.scala 31:69:@3458.4]
  assign _T_21796 = valid_10_25 ? 6'h19 : _T_21795; // @[Mux.scala 31:69:@3459.4]
  assign _T_21797 = valid_10_24 ? 6'h18 : _T_21796; // @[Mux.scala 31:69:@3460.4]
  assign _T_21798 = valid_10_23 ? 6'h17 : _T_21797; // @[Mux.scala 31:69:@3461.4]
  assign _T_21799 = valid_10_22 ? 6'h16 : _T_21798; // @[Mux.scala 31:69:@3462.4]
  assign _T_21800 = valid_10_21 ? 6'h15 : _T_21799; // @[Mux.scala 31:69:@3463.4]
  assign _T_21801 = valid_10_20 ? 6'h14 : _T_21800; // @[Mux.scala 31:69:@3464.4]
  assign _T_21802 = valid_10_19 ? 6'h13 : _T_21801; // @[Mux.scala 31:69:@3465.4]
  assign _T_21803 = valid_10_18 ? 6'h12 : _T_21802; // @[Mux.scala 31:69:@3466.4]
  assign _T_21804 = valid_10_17 ? 6'h11 : _T_21803; // @[Mux.scala 31:69:@3467.4]
  assign _T_21805 = valid_10_16 ? 6'h10 : _T_21804; // @[Mux.scala 31:69:@3468.4]
  assign _T_21806 = valid_10_15 ? 6'hf : _T_21805; // @[Mux.scala 31:69:@3469.4]
  assign _T_21807 = valid_10_14 ? 6'he : _T_21806; // @[Mux.scala 31:69:@3470.4]
  assign _T_21808 = valid_10_13 ? 6'hd : _T_21807; // @[Mux.scala 31:69:@3471.4]
  assign _T_21809 = valid_10_12 ? 6'hc : _T_21808; // @[Mux.scala 31:69:@3472.4]
  assign _T_21810 = valid_10_11 ? 6'hb : _T_21809; // @[Mux.scala 31:69:@3473.4]
  assign _T_21811 = valid_10_10 ? 6'ha : _T_21810; // @[Mux.scala 31:69:@3474.4]
  assign _T_21812 = valid_10_9 ? 6'h9 : _T_21811; // @[Mux.scala 31:69:@3475.4]
  assign _T_21813 = valid_10_8 ? 6'h8 : _T_21812; // @[Mux.scala 31:69:@3476.4]
  assign _T_21814 = valid_10_7 ? 6'h7 : _T_21813; // @[Mux.scala 31:69:@3477.4]
  assign _T_21815 = valid_10_6 ? 6'h6 : _T_21814; // @[Mux.scala 31:69:@3478.4]
  assign _T_21816 = valid_10_5 ? 6'h5 : _T_21815; // @[Mux.scala 31:69:@3479.4]
  assign _T_21817 = valid_10_4 ? 6'h4 : _T_21816; // @[Mux.scala 31:69:@3480.4]
  assign _T_21818 = valid_10_3 ? 6'h3 : _T_21817; // @[Mux.scala 31:69:@3481.4]
  assign _T_21819 = valid_10_2 ? 6'h2 : _T_21818; // @[Mux.scala 31:69:@3482.4]
  assign _T_21820 = valid_10_1 ? 6'h1 : _T_21819; // @[Mux.scala 31:69:@3483.4]
  assign select_10 = valid_10_0 ? 6'h0 : _T_21820; // @[Mux.scala 31:69:@3484.4]
  assign _GEN_641 = 6'h1 == select_10 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_642 = 6'h2 == select_10 ? io_inData_2 : _GEN_641; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_643 = 6'h3 == select_10 ? io_inData_3 : _GEN_642; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_644 = 6'h4 == select_10 ? io_inData_4 : _GEN_643; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_645 = 6'h5 == select_10 ? io_inData_5 : _GEN_644; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_646 = 6'h6 == select_10 ? io_inData_6 : _GEN_645; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_647 = 6'h7 == select_10 ? io_inData_7 : _GEN_646; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_648 = 6'h8 == select_10 ? io_inData_8 : _GEN_647; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_649 = 6'h9 == select_10 ? io_inData_9 : _GEN_648; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_650 = 6'ha == select_10 ? io_inData_10 : _GEN_649; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_651 = 6'hb == select_10 ? io_inData_11 : _GEN_650; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_652 = 6'hc == select_10 ? io_inData_12 : _GEN_651; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_653 = 6'hd == select_10 ? io_inData_13 : _GEN_652; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_654 = 6'he == select_10 ? io_inData_14 : _GEN_653; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_655 = 6'hf == select_10 ? io_inData_15 : _GEN_654; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_656 = 6'h10 == select_10 ? io_inData_16 : _GEN_655; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_657 = 6'h11 == select_10 ? io_inData_17 : _GEN_656; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_658 = 6'h12 == select_10 ? io_inData_18 : _GEN_657; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_659 = 6'h13 == select_10 ? io_inData_19 : _GEN_658; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_660 = 6'h14 == select_10 ? io_inData_20 : _GEN_659; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_661 = 6'h15 == select_10 ? io_inData_21 : _GEN_660; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_662 = 6'h16 == select_10 ? io_inData_22 : _GEN_661; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_663 = 6'h17 == select_10 ? io_inData_23 : _GEN_662; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_664 = 6'h18 == select_10 ? io_inData_24 : _GEN_663; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_665 = 6'h19 == select_10 ? io_inData_25 : _GEN_664; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_666 = 6'h1a == select_10 ? io_inData_26 : _GEN_665; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_667 = 6'h1b == select_10 ? io_inData_27 : _GEN_666; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_668 = 6'h1c == select_10 ? io_inData_28 : _GEN_667; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_669 = 6'h1d == select_10 ? io_inData_29 : _GEN_668; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_670 = 6'h1e == select_10 ? io_inData_30 : _GEN_669; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_671 = 6'h1f == select_10 ? io_inData_31 : _GEN_670; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_672 = 6'h20 == select_10 ? io_inData_32 : _GEN_671; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_673 = 6'h21 == select_10 ? io_inData_33 : _GEN_672; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_674 = 6'h22 == select_10 ? io_inData_34 : _GEN_673; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_675 = 6'h23 == select_10 ? io_inData_35 : _GEN_674; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_676 = 6'h24 == select_10 ? io_inData_36 : _GEN_675; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_677 = 6'h25 == select_10 ? io_inData_37 : _GEN_676; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_678 = 6'h26 == select_10 ? io_inData_38 : _GEN_677; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_679 = 6'h27 == select_10 ? io_inData_39 : _GEN_678; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_680 = 6'h28 == select_10 ? io_inData_40 : _GEN_679; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_681 = 6'h29 == select_10 ? io_inData_41 : _GEN_680; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_682 = 6'h2a == select_10 ? io_inData_42 : _GEN_681; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_683 = 6'h2b == select_10 ? io_inData_43 : _GEN_682; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_684 = 6'h2c == select_10 ? io_inData_44 : _GEN_683; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_685 = 6'h2d == select_10 ? io_inData_45 : _GEN_684; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_686 = 6'h2e == select_10 ? io_inData_46 : _GEN_685; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_687 = 6'h2f == select_10 ? io_inData_47 : _GEN_686; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_688 = 6'h30 == select_10 ? io_inData_48 : _GEN_687; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_689 = 6'h31 == select_10 ? io_inData_49 : _GEN_688; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_690 = 6'h32 == select_10 ? io_inData_50 : _GEN_689; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_691 = 6'h33 == select_10 ? io_inData_51 : _GEN_690; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_692 = 6'h34 == select_10 ? io_inData_52 : _GEN_691; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_693 = 6'h35 == select_10 ? io_inData_53 : _GEN_692; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_694 = 6'h36 == select_10 ? io_inData_54 : _GEN_693; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_695 = 6'h37 == select_10 ? io_inData_55 : _GEN_694; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_696 = 6'h38 == select_10 ? io_inData_56 : _GEN_695; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_697 = 6'h39 == select_10 ? io_inData_57 : _GEN_696; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_698 = 6'h3a == select_10 ? io_inData_58 : _GEN_697; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_699 = 6'h3b == select_10 ? io_inData_59 : _GEN_698; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_700 = 6'h3c == select_10 ? io_inData_60 : _GEN_699; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_701 = 6'h3d == select_10 ? io_inData_61 : _GEN_700; // @[Switch.scala 33:19:@3486.4]
  assign _GEN_702 = 6'h3e == select_10 ? io_inData_62 : _GEN_701; // @[Switch.scala 33:19:@3486.4]
  assign _T_21829 = {valid_10_7,valid_10_6,valid_10_5,valid_10_4,valid_10_3,valid_10_2,valid_10_1,valid_10_0}; // @[Switch.scala 34:32:@3493.4]
  assign _T_21837 = {valid_10_15,valid_10_14,valid_10_13,valid_10_12,valid_10_11,valid_10_10,valid_10_9,valid_10_8,_T_21829}; // @[Switch.scala 34:32:@3501.4]
  assign _T_21844 = {valid_10_23,valid_10_22,valid_10_21,valid_10_20,valid_10_19,valid_10_18,valid_10_17,valid_10_16}; // @[Switch.scala 34:32:@3508.4]
  assign _T_21853 = {valid_10_31,valid_10_30,valid_10_29,valid_10_28,valid_10_27,valid_10_26,valid_10_25,valid_10_24,_T_21844,_T_21837}; // @[Switch.scala 34:32:@3517.4]
  assign _T_21860 = {valid_10_39,valid_10_38,valid_10_37,valid_10_36,valid_10_35,valid_10_34,valid_10_33,valid_10_32}; // @[Switch.scala 34:32:@3524.4]
  assign _T_21868 = {valid_10_47,valid_10_46,valid_10_45,valid_10_44,valid_10_43,valid_10_42,valid_10_41,valid_10_40,_T_21860}; // @[Switch.scala 34:32:@3532.4]
  assign _T_21875 = {valid_10_55,valid_10_54,valid_10_53,valid_10_52,valid_10_51,valid_10_50,valid_10_49,valid_10_48}; // @[Switch.scala 34:32:@3539.4]
  assign _T_21884 = {valid_10_63,valid_10_62,valid_10_61,valid_10_60,valid_10_59,valid_10_58,valid_10_57,valid_10_56,_T_21875,_T_21868}; // @[Switch.scala 34:32:@3548.4]
  assign _T_21885 = {_T_21884,_T_21853}; // @[Switch.scala 34:32:@3549.4]
  assign _T_21889 = io_inAddr_0 == 6'hb; // @[Switch.scala 30:53:@3552.4]
  assign valid_11_0 = io_inValid_0 & _T_21889; // @[Switch.scala 30:36:@3553.4]
  assign _T_21892 = io_inAddr_1 == 6'hb; // @[Switch.scala 30:53:@3555.4]
  assign valid_11_1 = io_inValid_1 & _T_21892; // @[Switch.scala 30:36:@3556.4]
  assign _T_21895 = io_inAddr_2 == 6'hb; // @[Switch.scala 30:53:@3558.4]
  assign valid_11_2 = io_inValid_2 & _T_21895; // @[Switch.scala 30:36:@3559.4]
  assign _T_21898 = io_inAddr_3 == 6'hb; // @[Switch.scala 30:53:@3561.4]
  assign valid_11_3 = io_inValid_3 & _T_21898; // @[Switch.scala 30:36:@3562.4]
  assign _T_21901 = io_inAddr_4 == 6'hb; // @[Switch.scala 30:53:@3564.4]
  assign valid_11_4 = io_inValid_4 & _T_21901; // @[Switch.scala 30:36:@3565.4]
  assign _T_21904 = io_inAddr_5 == 6'hb; // @[Switch.scala 30:53:@3567.4]
  assign valid_11_5 = io_inValid_5 & _T_21904; // @[Switch.scala 30:36:@3568.4]
  assign _T_21907 = io_inAddr_6 == 6'hb; // @[Switch.scala 30:53:@3570.4]
  assign valid_11_6 = io_inValid_6 & _T_21907; // @[Switch.scala 30:36:@3571.4]
  assign _T_21910 = io_inAddr_7 == 6'hb; // @[Switch.scala 30:53:@3573.4]
  assign valid_11_7 = io_inValid_7 & _T_21910; // @[Switch.scala 30:36:@3574.4]
  assign _T_21913 = io_inAddr_8 == 6'hb; // @[Switch.scala 30:53:@3576.4]
  assign valid_11_8 = io_inValid_8 & _T_21913; // @[Switch.scala 30:36:@3577.4]
  assign _T_21916 = io_inAddr_9 == 6'hb; // @[Switch.scala 30:53:@3579.4]
  assign valid_11_9 = io_inValid_9 & _T_21916; // @[Switch.scala 30:36:@3580.4]
  assign _T_21919 = io_inAddr_10 == 6'hb; // @[Switch.scala 30:53:@3582.4]
  assign valid_11_10 = io_inValid_10 & _T_21919; // @[Switch.scala 30:36:@3583.4]
  assign _T_21922 = io_inAddr_11 == 6'hb; // @[Switch.scala 30:53:@3585.4]
  assign valid_11_11 = io_inValid_11 & _T_21922; // @[Switch.scala 30:36:@3586.4]
  assign _T_21925 = io_inAddr_12 == 6'hb; // @[Switch.scala 30:53:@3588.4]
  assign valid_11_12 = io_inValid_12 & _T_21925; // @[Switch.scala 30:36:@3589.4]
  assign _T_21928 = io_inAddr_13 == 6'hb; // @[Switch.scala 30:53:@3591.4]
  assign valid_11_13 = io_inValid_13 & _T_21928; // @[Switch.scala 30:36:@3592.4]
  assign _T_21931 = io_inAddr_14 == 6'hb; // @[Switch.scala 30:53:@3594.4]
  assign valid_11_14 = io_inValid_14 & _T_21931; // @[Switch.scala 30:36:@3595.4]
  assign _T_21934 = io_inAddr_15 == 6'hb; // @[Switch.scala 30:53:@3597.4]
  assign valid_11_15 = io_inValid_15 & _T_21934; // @[Switch.scala 30:36:@3598.4]
  assign _T_21937 = io_inAddr_16 == 6'hb; // @[Switch.scala 30:53:@3600.4]
  assign valid_11_16 = io_inValid_16 & _T_21937; // @[Switch.scala 30:36:@3601.4]
  assign _T_21940 = io_inAddr_17 == 6'hb; // @[Switch.scala 30:53:@3603.4]
  assign valid_11_17 = io_inValid_17 & _T_21940; // @[Switch.scala 30:36:@3604.4]
  assign _T_21943 = io_inAddr_18 == 6'hb; // @[Switch.scala 30:53:@3606.4]
  assign valid_11_18 = io_inValid_18 & _T_21943; // @[Switch.scala 30:36:@3607.4]
  assign _T_21946 = io_inAddr_19 == 6'hb; // @[Switch.scala 30:53:@3609.4]
  assign valid_11_19 = io_inValid_19 & _T_21946; // @[Switch.scala 30:36:@3610.4]
  assign _T_21949 = io_inAddr_20 == 6'hb; // @[Switch.scala 30:53:@3612.4]
  assign valid_11_20 = io_inValid_20 & _T_21949; // @[Switch.scala 30:36:@3613.4]
  assign _T_21952 = io_inAddr_21 == 6'hb; // @[Switch.scala 30:53:@3615.4]
  assign valid_11_21 = io_inValid_21 & _T_21952; // @[Switch.scala 30:36:@3616.4]
  assign _T_21955 = io_inAddr_22 == 6'hb; // @[Switch.scala 30:53:@3618.4]
  assign valid_11_22 = io_inValid_22 & _T_21955; // @[Switch.scala 30:36:@3619.4]
  assign _T_21958 = io_inAddr_23 == 6'hb; // @[Switch.scala 30:53:@3621.4]
  assign valid_11_23 = io_inValid_23 & _T_21958; // @[Switch.scala 30:36:@3622.4]
  assign _T_21961 = io_inAddr_24 == 6'hb; // @[Switch.scala 30:53:@3624.4]
  assign valid_11_24 = io_inValid_24 & _T_21961; // @[Switch.scala 30:36:@3625.4]
  assign _T_21964 = io_inAddr_25 == 6'hb; // @[Switch.scala 30:53:@3627.4]
  assign valid_11_25 = io_inValid_25 & _T_21964; // @[Switch.scala 30:36:@3628.4]
  assign _T_21967 = io_inAddr_26 == 6'hb; // @[Switch.scala 30:53:@3630.4]
  assign valid_11_26 = io_inValid_26 & _T_21967; // @[Switch.scala 30:36:@3631.4]
  assign _T_21970 = io_inAddr_27 == 6'hb; // @[Switch.scala 30:53:@3633.4]
  assign valid_11_27 = io_inValid_27 & _T_21970; // @[Switch.scala 30:36:@3634.4]
  assign _T_21973 = io_inAddr_28 == 6'hb; // @[Switch.scala 30:53:@3636.4]
  assign valid_11_28 = io_inValid_28 & _T_21973; // @[Switch.scala 30:36:@3637.4]
  assign _T_21976 = io_inAddr_29 == 6'hb; // @[Switch.scala 30:53:@3639.4]
  assign valid_11_29 = io_inValid_29 & _T_21976; // @[Switch.scala 30:36:@3640.4]
  assign _T_21979 = io_inAddr_30 == 6'hb; // @[Switch.scala 30:53:@3642.4]
  assign valid_11_30 = io_inValid_30 & _T_21979; // @[Switch.scala 30:36:@3643.4]
  assign _T_21982 = io_inAddr_31 == 6'hb; // @[Switch.scala 30:53:@3645.4]
  assign valid_11_31 = io_inValid_31 & _T_21982; // @[Switch.scala 30:36:@3646.4]
  assign _T_21985 = io_inAddr_32 == 6'hb; // @[Switch.scala 30:53:@3648.4]
  assign valid_11_32 = io_inValid_32 & _T_21985; // @[Switch.scala 30:36:@3649.4]
  assign _T_21988 = io_inAddr_33 == 6'hb; // @[Switch.scala 30:53:@3651.4]
  assign valid_11_33 = io_inValid_33 & _T_21988; // @[Switch.scala 30:36:@3652.4]
  assign _T_21991 = io_inAddr_34 == 6'hb; // @[Switch.scala 30:53:@3654.4]
  assign valid_11_34 = io_inValid_34 & _T_21991; // @[Switch.scala 30:36:@3655.4]
  assign _T_21994 = io_inAddr_35 == 6'hb; // @[Switch.scala 30:53:@3657.4]
  assign valid_11_35 = io_inValid_35 & _T_21994; // @[Switch.scala 30:36:@3658.4]
  assign _T_21997 = io_inAddr_36 == 6'hb; // @[Switch.scala 30:53:@3660.4]
  assign valid_11_36 = io_inValid_36 & _T_21997; // @[Switch.scala 30:36:@3661.4]
  assign _T_22000 = io_inAddr_37 == 6'hb; // @[Switch.scala 30:53:@3663.4]
  assign valid_11_37 = io_inValid_37 & _T_22000; // @[Switch.scala 30:36:@3664.4]
  assign _T_22003 = io_inAddr_38 == 6'hb; // @[Switch.scala 30:53:@3666.4]
  assign valid_11_38 = io_inValid_38 & _T_22003; // @[Switch.scala 30:36:@3667.4]
  assign _T_22006 = io_inAddr_39 == 6'hb; // @[Switch.scala 30:53:@3669.4]
  assign valid_11_39 = io_inValid_39 & _T_22006; // @[Switch.scala 30:36:@3670.4]
  assign _T_22009 = io_inAddr_40 == 6'hb; // @[Switch.scala 30:53:@3672.4]
  assign valid_11_40 = io_inValid_40 & _T_22009; // @[Switch.scala 30:36:@3673.4]
  assign _T_22012 = io_inAddr_41 == 6'hb; // @[Switch.scala 30:53:@3675.4]
  assign valid_11_41 = io_inValid_41 & _T_22012; // @[Switch.scala 30:36:@3676.4]
  assign _T_22015 = io_inAddr_42 == 6'hb; // @[Switch.scala 30:53:@3678.4]
  assign valid_11_42 = io_inValid_42 & _T_22015; // @[Switch.scala 30:36:@3679.4]
  assign _T_22018 = io_inAddr_43 == 6'hb; // @[Switch.scala 30:53:@3681.4]
  assign valid_11_43 = io_inValid_43 & _T_22018; // @[Switch.scala 30:36:@3682.4]
  assign _T_22021 = io_inAddr_44 == 6'hb; // @[Switch.scala 30:53:@3684.4]
  assign valid_11_44 = io_inValid_44 & _T_22021; // @[Switch.scala 30:36:@3685.4]
  assign _T_22024 = io_inAddr_45 == 6'hb; // @[Switch.scala 30:53:@3687.4]
  assign valid_11_45 = io_inValid_45 & _T_22024; // @[Switch.scala 30:36:@3688.4]
  assign _T_22027 = io_inAddr_46 == 6'hb; // @[Switch.scala 30:53:@3690.4]
  assign valid_11_46 = io_inValid_46 & _T_22027; // @[Switch.scala 30:36:@3691.4]
  assign _T_22030 = io_inAddr_47 == 6'hb; // @[Switch.scala 30:53:@3693.4]
  assign valid_11_47 = io_inValid_47 & _T_22030; // @[Switch.scala 30:36:@3694.4]
  assign _T_22033 = io_inAddr_48 == 6'hb; // @[Switch.scala 30:53:@3696.4]
  assign valid_11_48 = io_inValid_48 & _T_22033; // @[Switch.scala 30:36:@3697.4]
  assign _T_22036 = io_inAddr_49 == 6'hb; // @[Switch.scala 30:53:@3699.4]
  assign valid_11_49 = io_inValid_49 & _T_22036; // @[Switch.scala 30:36:@3700.4]
  assign _T_22039 = io_inAddr_50 == 6'hb; // @[Switch.scala 30:53:@3702.4]
  assign valid_11_50 = io_inValid_50 & _T_22039; // @[Switch.scala 30:36:@3703.4]
  assign _T_22042 = io_inAddr_51 == 6'hb; // @[Switch.scala 30:53:@3705.4]
  assign valid_11_51 = io_inValid_51 & _T_22042; // @[Switch.scala 30:36:@3706.4]
  assign _T_22045 = io_inAddr_52 == 6'hb; // @[Switch.scala 30:53:@3708.4]
  assign valid_11_52 = io_inValid_52 & _T_22045; // @[Switch.scala 30:36:@3709.4]
  assign _T_22048 = io_inAddr_53 == 6'hb; // @[Switch.scala 30:53:@3711.4]
  assign valid_11_53 = io_inValid_53 & _T_22048; // @[Switch.scala 30:36:@3712.4]
  assign _T_22051 = io_inAddr_54 == 6'hb; // @[Switch.scala 30:53:@3714.4]
  assign valid_11_54 = io_inValid_54 & _T_22051; // @[Switch.scala 30:36:@3715.4]
  assign _T_22054 = io_inAddr_55 == 6'hb; // @[Switch.scala 30:53:@3717.4]
  assign valid_11_55 = io_inValid_55 & _T_22054; // @[Switch.scala 30:36:@3718.4]
  assign _T_22057 = io_inAddr_56 == 6'hb; // @[Switch.scala 30:53:@3720.4]
  assign valid_11_56 = io_inValid_56 & _T_22057; // @[Switch.scala 30:36:@3721.4]
  assign _T_22060 = io_inAddr_57 == 6'hb; // @[Switch.scala 30:53:@3723.4]
  assign valid_11_57 = io_inValid_57 & _T_22060; // @[Switch.scala 30:36:@3724.4]
  assign _T_22063 = io_inAddr_58 == 6'hb; // @[Switch.scala 30:53:@3726.4]
  assign valid_11_58 = io_inValid_58 & _T_22063; // @[Switch.scala 30:36:@3727.4]
  assign _T_22066 = io_inAddr_59 == 6'hb; // @[Switch.scala 30:53:@3729.4]
  assign valid_11_59 = io_inValid_59 & _T_22066; // @[Switch.scala 30:36:@3730.4]
  assign _T_22069 = io_inAddr_60 == 6'hb; // @[Switch.scala 30:53:@3732.4]
  assign valid_11_60 = io_inValid_60 & _T_22069; // @[Switch.scala 30:36:@3733.4]
  assign _T_22072 = io_inAddr_61 == 6'hb; // @[Switch.scala 30:53:@3735.4]
  assign valid_11_61 = io_inValid_61 & _T_22072; // @[Switch.scala 30:36:@3736.4]
  assign _T_22075 = io_inAddr_62 == 6'hb; // @[Switch.scala 30:53:@3738.4]
  assign valid_11_62 = io_inValid_62 & _T_22075; // @[Switch.scala 30:36:@3739.4]
  assign _T_22078 = io_inAddr_63 == 6'hb; // @[Switch.scala 30:53:@3741.4]
  assign valid_11_63 = io_inValid_63 & _T_22078; // @[Switch.scala 30:36:@3742.4]
  assign _T_22144 = valid_11_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@3744.4]
  assign _T_22145 = valid_11_61 ? 6'h3d : _T_22144; // @[Mux.scala 31:69:@3745.4]
  assign _T_22146 = valid_11_60 ? 6'h3c : _T_22145; // @[Mux.scala 31:69:@3746.4]
  assign _T_22147 = valid_11_59 ? 6'h3b : _T_22146; // @[Mux.scala 31:69:@3747.4]
  assign _T_22148 = valid_11_58 ? 6'h3a : _T_22147; // @[Mux.scala 31:69:@3748.4]
  assign _T_22149 = valid_11_57 ? 6'h39 : _T_22148; // @[Mux.scala 31:69:@3749.4]
  assign _T_22150 = valid_11_56 ? 6'h38 : _T_22149; // @[Mux.scala 31:69:@3750.4]
  assign _T_22151 = valid_11_55 ? 6'h37 : _T_22150; // @[Mux.scala 31:69:@3751.4]
  assign _T_22152 = valid_11_54 ? 6'h36 : _T_22151; // @[Mux.scala 31:69:@3752.4]
  assign _T_22153 = valid_11_53 ? 6'h35 : _T_22152; // @[Mux.scala 31:69:@3753.4]
  assign _T_22154 = valid_11_52 ? 6'h34 : _T_22153; // @[Mux.scala 31:69:@3754.4]
  assign _T_22155 = valid_11_51 ? 6'h33 : _T_22154; // @[Mux.scala 31:69:@3755.4]
  assign _T_22156 = valid_11_50 ? 6'h32 : _T_22155; // @[Mux.scala 31:69:@3756.4]
  assign _T_22157 = valid_11_49 ? 6'h31 : _T_22156; // @[Mux.scala 31:69:@3757.4]
  assign _T_22158 = valid_11_48 ? 6'h30 : _T_22157; // @[Mux.scala 31:69:@3758.4]
  assign _T_22159 = valid_11_47 ? 6'h2f : _T_22158; // @[Mux.scala 31:69:@3759.4]
  assign _T_22160 = valid_11_46 ? 6'h2e : _T_22159; // @[Mux.scala 31:69:@3760.4]
  assign _T_22161 = valid_11_45 ? 6'h2d : _T_22160; // @[Mux.scala 31:69:@3761.4]
  assign _T_22162 = valid_11_44 ? 6'h2c : _T_22161; // @[Mux.scala 31:69:@3762.4]
  assign _T_22163 = valid_11_43 ? 6'h2b : _T_22162; // @[Mux.scala 31:69:@3763.4]
  assign _T_22164 = valid_11_42 ? 6'h2a : _T_22163; // @[Mux.scala 31:69:@3764.4]
  assign _T_22165 = valid_11_41 ? 6'h29 : _T_22164; // @[Mux.scala 31:69:@3765.4]
  assign _T_22166 = valid_11_40 ? 6'h28 : _T_22165; // @[Mux.scala 31:69:@3766.4]
  assign _T_22167 = valid_11_39 ? 6'h27 : _T_22166; // @[Mux.scala 31:69:@3767.4]
  assign _T_22168 = valid_11_38 ? 6'h26 : _T_22167; // @[Mux.scala 31:69:@3768.4]
  assign _T_22169 = valid_11_37 ? 6'h25 : _T_22168; // @[Mux.scala 31:69:@3769.4]
  assign _T_22170 = valid_11_36 ? 6'h24 : _T_22169; // @[Mux.scala 31:69:@3770.4]
  assign _T_22171 = valid_11_35 ? 6'h23 : _T_22170; // @[Mux.scala 31:69:@3771.4]
  assign _T_22172 = valid_11_34 ? 6'h22 : _T_22171; // @[Mux.scala 31:69:@3772.4]
  assign _T_22173 = valid_11_33 ? 6'h21 : _T_22172; // @[Mux.scala 31:69:@3773.4]
  assign _T_22174 = valid_11_32 ? 6'h20 : _T_22173; // @[Mux.scala 31:69:@3774.4]
  assign _T_22175 = valid_11_31 ? 6'h1f : _T_22174; // @[Mux.scala 31:69:@3775.4]
  assign _T_22176 = valid_11_30 ? 6'h1e : _T_22175; // @[Mux.scala 31:69:@3776.4]
  assign _T_22177 = valid_11_29 ? 6'h1d : _T_22176; // @[Mux.scala 31:69:@3777.4]
  assign _T_22178 = valid_11_28 ? 6'h1c : _T_22177; // @[Mux.scala 31:69:@3778.4]
  assign _T_22179 = valid_11_27 ? 6'h1b : _T_22178; // @[Mux.scala 31:69:@3779.4]
  assign _T_22180 = valid_11_26 ? 6'h1a : _T_22179; // @[Mux.scala 31:69:@3780.4]
  assign _T_22181 = valid_11_25 ? 6'h19 : _T_22180; // @[Mux.scala 31:69:@3781.4]
  assign _T_22182 = valid_11_24 ? 6'h18 : _T_22181; // @[Mux.scala 31:69:@3782.4]
  assign _T_22183 = valid_11_23 ? 6'h17 : _T_22182; // @[Mux.scala 31:69:@3783.4]
  assign _T_22184 = valid_11_22 ? 6'h16 : _T_22183; // @[Mux.scala 31:69:@3784.4]
  assign _T_22185 = valid_11_21 ? 6'h15 : _T_22184; // @[Mux.scala 31:69:@3785.4]
  assign _T_22186 = valid_11_20 ? 6'h14 : _T_22185; // @[Mux.scala 31:69:@3786.4]
  assign _T_22187 = valid_11_19 ? 6'h13 : _T_22186; // @[Mux.scala 31:69:@3787.4]
  assign _T_22188 = valid_11_18 ? 6'h12 : _T_22187; // @[Mux.scala 31:69:@3788.4]
  assign _T_22189 = valid_11_17 ? 6'h11 : _T_22188; // @[Mux.scala 31:69:@3789.4]
  assign _T_22190 = valid_11_16 ? 6'h10 : _T_22189; // @[Mux.scala 31:69:@3790.4]
  assign _T_22191 = valid_11_15 ? 6'hf : _T_22190; // @[Mux.scala 31:69:@3791.4]
  assign _T_22192 = valid_11_14 ? 6'he : _T_22191; // @[Mux.scala 31:69:@3792.4]
  assign _T_22193 = valid_11_13 ? 6'hd : _T_22192; // @[Mux.scala 31:69:@3793.4]
  assign _T_22194 = valid_11_12 ? 6'hc : _T_22193; // @[Mux.scala 31:69:@3794.4]
  assign _T_22195 = valid_11_11 ? 6'hb : _T_22194; // @[Mux.scala 31:69:@3795.4]
  assign _T_22196 = valid_11_10 ? 6'ha : _T_22195; // @[Mux.scala 31:69:@3796.4]
  assign _T_22197 = valid_11_9 ? 6'h9 : _T_22196; // @[Mux.scala 31:69:@3797.4]
  assign _T_22198 = valid_11_8 ? 6'h8 : _T_22197; // @[Mux.scala 31:69:@3798.4]
  assign _T_22199 = valid_11_7 ? 6'h7 : _T_22198; // @[Mux.scala 31:69:@3799.4]
  assign _T_22200 = valid_11_6 ? 6'h6 : _T_22199; // @[Mux.scala 31:69:@3800.4]
  assign _T_22201 = valid_11_5 ? 6'h5 : _T_22200; // @[Mux.scala 31:69:@3801.4]
  assign _T_22202 = valid_11_4 ? 6'h4 : _T_22201; // @[Mux.scala 31:69:@3802.4]
  assign _T_22203 = valid_11_3 ? 6'h3 : _T_22202; // @[Mux.scala 31:69:@3803.4]
  assign _T_22204 = valid_11_2 ? 6'h2 : _T_22203; // @[Mux.scala 31:69:@3804.4]
  assign _T_22205 = valid_11_1 ? 6'h1 : _T_22204; // @[Mux.scala 31:69:@3805.4]
  assign select_11 = valid_11_0 ? 6'h0 : _T_22205; // @[Mux.scala 31:69:@3806.4]
  assign _GEN_705 = 6'h1 == select_11 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_706 = 6'h2 == select_11 ? io_inData_2 : _GEN_705; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_707 = 6'h3 == select_11 ? io_inData_3 : _GEN_706; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_708 = 6'h4 == select_11 ? io_inData_4 : _GEN_707; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_709 = 6'h5 == select_11 ? io_inData_5 : _GEN_708; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_710 = 6'h6 == select_11 ? io_inData_6 : _GEN_709; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_711 = 6'h7 == select_11 ? io_inData_7 : _GEN_710; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_712 = 6'h8 == select_11 ? io_inData_8 : _GEN_711; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_713 = 6'h9 == select_11 ? io_inData_9 : _GEN_712; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_714 = 6'ha == select_11 ? io_inData_10 : _GEN_713; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_715 = 6'hb == select_11 ? io_inData_11 : _GEN_714; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_716 = 6'hc == select_11 ? io_inData_12 : _GEN_715; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_717 = 6'hd == select_11 ? io_inData_13 : _GEN_716; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_718 = 6'he == select_11 ? io_inData_14 : _GEN_717; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_719 = 6'hf == select_11 ? io_inData_15 : _GEN_718; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_720 = 6'h10 == select_11 ? io_inData_16 : _GEN_719; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_721 = 6'h11 == select_11 ? io_inData_17 : _GEN_720; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_722 = 6'h12 == select_11 ? io_inData_18 : _GEN_721; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_723 = 6'h13 == select_11 ? io_inData_19 : _GEN_722; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_724 = 6'h14 == select_11 ? io_inData_20 : _GEN_723; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_725 = 6'h15 == select_11 ? io_inData_21 : _GEN_724; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_726 = 6'h16 == select_11 ? io_inData_22 : _GEN_725; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_727 = 6'h17 == select_11 ? io_inData_23 : _GEN_726; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_728 = 6'h18 == select_11 ? io_inData_24 : _GEN_727; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_729 = 6'h19 == select_11 ? io_inData_25 : _GEN_728; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_730 = 6'h1a == select_11 ? io_inData_26 : _GEN_729; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_731 = 6'h1b == select_11 ? io_inData_27 : _GEN_730; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_732 = 6'h1c == select_11 ? io_inData_28 : _GEN_731; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_733 = 6'h1d == select_11 ? io_inData_29 : _GEN_732; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_734 = 6'h1e == select_11 ? io_inData_30 : _GEN_733; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_735 = 6'h1f == select_11 ? io_inData_31 : _GEN_734; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_736 = 6'h20 == select_11 ? io_inData_32 : _GEN_735; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_737 = 6'h21 == select_11 ? io_inData_33 : _GEN_736; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_738 = 6'h22 == select_11 ? io_inData_34 : _GEN_737; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_739 = 6'h23 == select_11 ? io_inData_35 : _GEN_738; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_740 = 6'h24 == select_11 ? io_inData_36 : _GEN_739; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_741 = 6'h25 == select_11 ? io_inData_37 : _GEN_740; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_742 = 6'h26 == select_11 ? io_inData_38 : _GEN_741; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_743 = 6'h27 == select_11 ? io_inData_39 : _GEN_742; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_744 = 6'h28 == select_11 ? io_inData_40 : _GEN_743; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_745 = 6'h29 == select_11 ? io_inData_41 : _GEN_744; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_746 = 6'h2a == select_11 ? io_inData_42 : _GEN_745; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_747 = 6'h2b == select_11 ? io_inData_43 : _GEN_746; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_748 = 6'h2c == select_11 ? io_inData_44 : _GEN_747; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_749 = 6'h2d == select_11 ? io_inData_45 : _GEN_748; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_750 = 6'h2e == select_11 ? io_inData_46 : _GEN_749; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_751 = 6'h2f == select_11 ? io_inData_47 : _GEN_750; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_752 = 6'h30 == select_11 ? io_inData_48 : _GEN_751; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_753 = 6'h31 == select_11 ? io_inData_49 : _GEN_752; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_754 = 6'h32 == select_11 ? io_inData_50 : _GEN_753; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_755 = 6'h33 == select_11 ? io_inData_51 : _GEN_754; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_756 = 6'h34 == select_11 ? io_inData_52 : _GEN_755; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_757 = 6'h35 == select_11 ? io_inData_53 : _GEN_756; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_758 = 6'h36 == select_11 ? io_inData_54 : _GEN_757; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_759 = 6'h37 == select_11 ? io_inData_55 : _GEN_758; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_760 = 6'h38 == select_11 ? io_inData_56 : _GEN_759; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_761 = 6'h39 == select_11 ? io_inData_57 : _GEN_760; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_762 = 6'h3a == select_11 ? io_inData_58 : _GEN_761; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_763 = 6'h3b == select_11 ? io_inData_59 : _GEN_762; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_764 = 6'h3c == select_11 ? io_inData_60 : _GEN_763; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_765 = 6'h3d == select_11 ? io_inData_61 : _GEN_764; // @[Switch.scala 33:19:@3808.4]
  assign _GEN_766 = 6'h3e == select_11 ? io_inData_62 : _GEN_765; // @[Switch.scala 33:19:@3808.4]
  assign _T_22214 = {valid_11_7,valid_11_6,valid_11_5,valid_11_4,valid_11_3,valid_11_2,valid_11_1,valid_11_0}; // @[Switch.scala 34:32:@3815.4]
  assign _T_22222 = {valid_11_15,valid_11_14,valid_11_13,valid_11_12,valid_11_11,valid_11_10,valid_11_9,valid_11_8,_T_22214}; // @[Switch.scala 34:32:@3823.4]
  assign _T_22229 = {valid_11_23,valid_11_22,valid_11_21,valid_11_20,valid_11_19,valid_11_18,valid_11_17,valid_11_16}; // @[Switch.scala 34:32:@3830.4]
  assign _T_22238 = {valid_11_31,valid_11_30,valid_11_29,valid_11_28,valid_11_27,valid_11_26,valid_11_25,valid_11_24,_T_22229,_T_22222}; // @[Switch.scala 34:32:@3839.4]
  assign _T_22245 = {valid_11_39,valid_11_38,valid_11_37,valid_11_36,valid_11_35,valid_11_34,valid_11_33,valid_11_32}; // @[Switch.scala 34:32:@3846.4]
  assign _T_22253 = {valid_11_47,valid_11_46,valid_11_45,valid_11_44,valid_11_43,valid_11_42,valid_11_41,valid_11_40,_T_22245}; // @[Switch.scala 34:32:@3854.4]
  assign _T_22260 = {valid_11_55,valid_11_54,valid_11_53,valid_11_52,valid_11_51,valid_11_50,valid_11_49,valid_11_48}; // @[Switch.scala 34:32:@3861.4]
  assign _T_22269 = {valid_11_63,valid_11_62,valid_11_61,valid_11_60,valid_11_59,valid_11_58,valid_11_57,valid_11_56,_T_22260,_T_22253}; // @[Switch.scala 34:32:@3870.4]
  assign _T_22270 = {_T_22269,_T_22238}; // @[Switch.scala 34:32:@3871.4]
  assign _T_22274 = io_inAddr_0 == 6'hc; // @[Switch.scala 30:53:@3874.4]
  assign valid_12_0 = io_inValid_0 & _T_22274; // @[Switch.scala 30:36:@3875.4]
  assign _T_22277 = io_inAddr_1 == 6'hc; // @[Switch.scala 30:53:@3877.4]
  assign valid_12_1 = io_inValid_1 & _T_22277; // @[Switch.scala 30:36:@3878.4]
  assign _T_22280 = io_inAddr_2 == 6'hc; // @[Switch.scala 30:53:@3880.4]
  assign valid_12_2 = io_inValid_2 & _T_22280; // @[Switch.scala 30:36:@3881.4]
  assign _T_22283 = io_inAddr_3 == 6'hc; // @[Switch.scala 30:53:@3883.4]
  assign valid_12_3 = io_inValid_3 & _T_22283; // @[Switch.scala 30:36:@3884.4]
  assign _T_22286 = io_inAddr_4 == 6'hc; // @[Switch.scala 30:53:@3886.4]
  assign valid_12_4 = io_inValid_4 & _T_22286; // @[Switch.scala 30:36:@3887.4]
  assign _T_22289 = io_inAddr_5 == 6'hc; // @[Switch.scala 30:53:@3889.4]
  assign valid_12_5 = io_inValid_5 & _T_22289; // @[Switch.scala 30:36:@3890.4]
  assign _T_22292 = io_inAddr_6 == 6'hc; // @[Switch.scala 30:53:@3892.4]
  assign valid_12_6 = io_inValid_6 & _T_22292; // @[Switch.scala 30:36:@3893.4]
  assign _T_22295 = io_inAddr_7 == 6'hc; // @[Switch.scala 30:53:@3895.4]
  assign valid_12_7 = io_inValid_7 & _T_22295; // @[Switch.scala 30:36:@3896.4]
  assign _T_22298 = io_inAddr_8 == 6'hc; // @[Switch.scala 30:53:@3898.4]
  assign valid_12_8 = io_inValid_8 & _T_22298; // @[Switch.scala 30:36:@3899.4]
  assign _T_22301 = io_inAddr_9 == 6'hc; // @[Switch.scala 30:53:@3901.4]
  assign valid_12_9 = io_inValid_9 & _T_22301; // @[Switch.scala 30:36:@3902.4]
  assign _T_22304 = io_inAddr_10 == 6'hc; // @[Switch.scala 30:53:@3904.4]
  assign valid_12_10 = io_inValid_10 & _T_22304; // @[Switch.scala 30:36:@3905.4]
  assign _T_22307 = io_inAddr_11 == 6'hc; // @[Switch.scala 30:53:@3907.4]
  assign valid_12_11 = io_inValid_11 & _T_22307; // @[Switch.scala 30:36:@3908.4]
  assign _T_22310 = io_inAddr_12 == 6'hc; // @[Switch.scala 30:53:@3910.4]
  assign valid_12_12 = io_inValid_12 & _T_22310; // @[Switch.scala 30:36:@3911.4]
  assign _T_22313 = io_inAddr_13 == 6'hc; // @[Switch.scala 30:53:@3913.4]
  assign valid_12_13 = io_inValid_13 & _T_22313; // @[Switch.scala 30:36:@3914.4]
  assign _T_22316 = io_inAddr_14 == 6'hc; // @[Switch.scala 30:53:@3916.4]
  assign valid_12_14 = io_inValid_14 & _T_22316; // @[Switch.scala 30:36:@3917.4]
  assign _T_22319 = io_inAddr_15 == 6'hc; // @[Switch.scala 30:53:@3919.4]
  assign valid_12_15 = io_inValid_15 & _T_22319; // @[Switch.scala 30:36:@3920.4]
  assign _T_22322 = io_inAddr_16 == 6'hc; // @[Switch.scala 30:53:@3922.4]
  assign valid_12_16 = io_inValid_16 & _T_22322; // @[Switch.scala 30:36:@3923.4]
  assign _T_22325 = io_inAddr_17 == 6'hc; // @[Switch.scala 30:53:@3925.4]
  assign valid_12_17 = io_inValid_17 & _T_22325; // @[Switch.scala 30:36:@3926.4]
  assign _T_22328 = io_inAddr_18 == 6'hc; // @[Switch.scala 30:53:@3928.4]
  assign valid_12_18 = io_inValid_18 & _T_22328; // @[Switch.scala 30:36:@3929.4]
  assign _T_22331 = io_inAddr_19 == 6'hc; // @[Switch.scala 30:53:@3931.4]
  assign valid_12_19 = io_inValid_19 & _T_22331; // @[Switch.scala 30:36:@3932.4]
  assign _T_22334 = io_inAddr_20 == 6'hc; // @[Switch.scala 30:53:@3934.4]
  assign valid_12_20 = io_inValid_20 & _T_22334; // @[Switch.scala 30:36:@3935.4]
  assign _T_22337 = io_inAddr_21 == 6'hc; // @[Switch.scala 30:53:@3937.4]
  assign valid_12_21 = io_inValid_21 & _T_22337; // @[Switch.scala 30:36:@3938.4]
  assign _T_22340 = io_inAddr_22 == 6'hc; // @[Switch.scala 30:53:@3940.4]
  assign valid_12_22 = io_inValid_22 & _T_22340; // @[Switch.scala 30:36:@3941.4]
  assign _T_22343 = io_inAddr_23 == 6'hc; // @[Switch.scala 30:53:@3943.4]
  assign valid_12_23 = io_inValid_23 & _T_22343; // @[Switch.scala 30:36:@3944.4]
  assign _T_22346 = io_inAddr_24 == 6'hc; // @[Switch.scala 30:53:@3946.4]
  assign valid_12_24 = io_inValid_24 & _T_22346; // @[Switch.scala 30:36:@3947.4]
  assign _T_22349 = io_inAddr_25 == 6'hc; // @[Switch.scala 30:53:@3949.4]
  assign valid_12_25 = io_inValid_25 & _T_22349; // @[Switch.scala 30:36:@3950.4]
  assign _T_22352 = io_inAddr_26 == 6'hc; // @[Switch.scala 30:53:@3952.4]
  assign valid_12_26 = io_inValid_26 & _T_22352; // @[Switch.scala 30:36:@3953.4]
  assign _T_22355 = io_inAddr_27 == 6'hc; // @[Switch.scala 30:53:@3955.4]
  assign valid_12_27 = io_inValid_27 & _T_22355; // @[Switch.scala 30:36:@3956.4]
  assign _T_22358 = io_inAddr_28 == 6'hc; // @[Switch.scala 30:53:@3958.4]
  assign valid_12_28 = io_inValid_28 & _T_22358; // @[Switch.scala 30:36:@3959.4]
  assign _T_22361 = io_inAddr_29 == 6'hc; // @[Switch.scala 30:53:@3961.4]
  assign valid_12_29 = io_inValid_29 & _T_22361; // @[Switch.scala 30:36:@3962.4]
  assign _T_22364 = io_inAddr_30 == 6'hc; // @[Switch.scala 30:53:@3964.4]
  assign valid_12_30 = io_inValid_30 & _T_22364; // @[Switch.scala 30:36:@3965.4]
  assign _T_22367 = io_inAddr_31 == 6'hc; // @[Switch.scala 30:53:@3967.4]
  assign valid_12_31 = io_inValid_31 & _T_22367; // @[Switch.scala 30:36:@3968.4]
  assign _T_22370 = io_inAddr_32 == 6'hc; // @[Switch.scala 30:53:@3970.4]
  assign valid_12_32 = io_inValid_32 & _T_22370; // @[Switch.scala 30:36:@3971.4]
  assign _T_22373 = io_inAddr_33 == 6'hc; // @[Switch.scala 30:53:@3973.4]
  assign valid_12_33 = io_inValid_33 & _T_22373; // @[Switch.scala 30:36:@3974.4]
  assign _T_22376 = io_inAddr_34 == 6'hc; // @[Switch.scala 30:53:@3976.4]
  assign valid_12_34 = io_inValid_34 & _T_22376; // @[Switch.scala 30:36:@3977.4]
  assign _T_22379 = io_inAddr_35 == 6'hc; // @[Switch.scala 30:53:@3979.4]
  assign valid_12_35 = io_inValid_35 & _T_22379; // @[Switch.scala 30:36:@3980.4]
  assign _T_22382 = io_inAddr_36 == 6'hc; // @[Switch.scala 30:53:@3982.4]
  assign valid_12_36 = io_inValid_36 & _T_22382; // @[Switch.scala 30:36:@3983.4]
  assign _T_22385 = io_inAddr_37 == 6'hc; // @[Switch.scala 30:53:@3985.4]
  assign valid_12_37 = io_inValid_37 & _T_22385; // @[Switch.scala 30:36:@3986.4]
  assign _T_22388 = io_inAddr_38 == 6'hc; // @[Switch.scala 30:53:@3988.4]
  assign valid_12_38 = io_inValid_38 & _T_22388; // @[Switch.scala 30:36:@3989.4]
  assign _T_22391 = io_inAddr_39 == 6'hc; // @[Switch.scala 30:53:@3991.4]
  assign valid_12_39 = io_inValid_39 & _T_22391; // @[Switch.scala 30:36:@3992.4]
  assign _T_22394 = io_inAddr_40 == 6'hc; // @[Switch.scala 30:53:@3994.4]
  assign valid_12_40 = io_inValid_40 & _T_22394; // @[Switch.scala 30:36:@3995.4]
  assign _T_22397 = io_inAddr_41 == 6'hc; // @[Switch.scala 30:53:@3997.4]
  assign valid_12_41 = io_inValid_41 & _T_22397; // @[Switch.scala 30:36:@3998.4]
  assign _T_22400 = io_inAddr_42 == 6'hc; // @[Switch.scala 30:53:@4000.4]
  assign valid_12_42 = io_inValid_42 & _T_22400; // @[Switch.scala 30:36:@4001.4]
  assign _T_22403 = io_inAddr_43 == 6'hc; // @[Switch.scala 30:53:@4003.4]
  assign valid_12_43 = io_inValid_43 & _T_22403; // @[Switch.scala 30:36:@4004.4]
  assign _T_22406 = io_inAddr_44 == 6'hc; // @[Switch.scala 30:53:@4006.4]
  assign valid_12_44 = io_inValid_44 & _T_22406; // @[Switch.scala 30:36:@4007.4]
  assign _T_22409 = io_inAddr_45 == 6'hc; // @[Switch.scala 30:53:@4009.4]
  assign valid_12_45 = io_inValid_45 & _T_22409; // @[Switch.scala 30:36:@4010.4]
  assign _T_22412 = io_inAddr_46 == 6'hc; // @[Switch.scala 30:53:@4012.4]
  assign valid_12_46 = io_inValid_46 & _T_22412; // @[Switch.scala 30:36:@4013.4]
  assign _T_22415 = io_inAddr_47 == 6'hc; // @[Switch.scala 30:53:@4015.4]
  assign valid_12_47 = io_inValid_47 & _T_22415; // @[Switch.scala 30:36:@4016.4]
  assign _T_22418 = io_inAddr_48 == 6'hc; // @[Switch.scala 30:53:@4018.4]
  assign valid_12_48 = io_inValid_48 & _T_22418; // @[Switch.scala 30:36:@4019.4]
  assign _T_22421 = io_inAddr_49 == 6'hc; // @[Switch.scala 30:53:@4021.4]
  assign valid_12_49 = io_inValid_49 & _T_22421; // @[Switch.scala 30:36:@4022.4]
  assign _T_22424 = io_inAddr_50 == 6'hc; // @[Switch.scala 30:53:@4024.4]
  assign valid_12_50 = io_inValid_50 & _T_22424; // @[Switch.scala 30:36:@4025.4]
  assign _T_22427 = io_inAddr_51 == 6'hc; // @[Switch.scala 30:53:@4027.4]
  assign valid_12_51 = io_inValid_51 & _T_22427; // @[Switch.scala 30:36:@4028.4]
  assign _T_22430 = io_inAddr_52 == 6'hc; // @[Switch.scala 30:53:@4030.4]
  assign valid_12_52 = io_inValid_52 & _T_22430; // @[Switch.scala 30:36:@4031.4]
  assign _T_22433 = io_inAddr_53 == 6'hc; // @[Switch.scala 30:53:@4033.4]
  assign valid_12_53 = io_inValid_53 & _T_22433; // @[Switch.scala 30:36:@4034.4]
  assign _T_22436 = io_inAddr_54 == 6'hc; // @[Switch.scala 30:53:@4036.4]
  assign valid_12_54 = io_inValid_54 & _T_22436; // @[Switch.scala 30:36:@4037.4]
  assign _T_22439 = io_inAddr_55 == 6'hc; // @[Switch.scala 30:53:@4039.4]
  assign valid_12_55 = io_inValid_55 & _T_22439; // @[Switch.scala 30:36:@4040.4]
  assign _T_22442 = io_inAddr_56 == 6'hc; // @[Switch.scala 30:53:@4042.4]
  assign valid_12_56 = io_inValid_56 & _T_22442; // @[Switch.scala 30:36:@4043.4]
  assign _T_22445 = io_inAddr_57 == 6'hc; // @[Switch.scala 30:53:@4045.4]
  assign valid_12_57 = io_inValid_57 & _T_22445; // @[Switch.scala 30:36:@4046.4]
  assign _T_22448 = io_inAddr_58 == 6'hc; // @[Switch.scala 30:53:@4048.4]
  assign valid_12_58 = io_inValid_58 & _T_22448; // @[Switch.scala 30:36:@4049.4]
  assign _T_22451 = io_inAddr_59 == 6'hc; // @[Switch.scala 30:53:@4051.4]
  assign valid_12_59 = io_inValid_59 & _T_22451; // @[Switch.scala 30:36:@4052.4]
  assign _T_22454 = io_inAddr_60 == 6'hc; // @[Switch.scala 30:53:@4054.4]
  assign valid_12_60 = io_inValid_60 & _T_22454; // @[Switch.scala 30:36:@4055.4]
  assign _T_22457 = io_inAddr_61 == 6'hc; // @[Switch.scala 30:53:@4057.4]
  assign valid_12_61 = io_inValid_61 & _T_22457; // @[Switch.scala 30:36:@4058.4]
  assign _T_22460 = io_inAddr_62 == 6'hc; // @[Switch.scala 30:53:@4060.4]
  assign valid_12_62 = io_inValid_62 & _T_22460; // @[Switch.scala 30:36:@4061.4]
  assign _T_22463 = io_inAddr_63 == 6'hc; // @[Switch.scala 30:53:@4063.4]
  assign valid_12_63 = io_inValid_63 & _T_22463; // @[Switch.scala 30:36:@4064.4]
  assign _T_22529 = valid_12_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@4066.4]
  assign _T_22530 = valid_12_61 ? 6'h3d : _T_22529; // @[Mux.scala 31:69:@4067.4]
  assign _T_22531 = valid_12_60 ? 6'h3c : _T_22530; // @[Mux.scala 31:69:@4068.4]
  assign _T_22532 = valid_12_59 ? 6'h3b : _T_22531; // @[Mux.scala 31:69:@4069.4]
  assign _T_22533 = valid_12_58 ? 6'h3a : _T_22532; // @[Mux.scala 31:69:@4070.4]
  assign _T_22534 = valid_12_57 ? 6'h39 : _T_22533; // @[Mux.scala 31:69:@4071.4]
  assign _T_22535 = valid_12_56 ? 6'h38 : _T_22534; // @[Mux.scala 31:69:@4072.4]
  assign _T_22536 = valid_12_55 ? 6'h37 : _T_22535; // @[Mux.scala 31:69:@4073.4]
  assign _T_22537 = valid_12_54 ? 6'h36 : _T_22536; // @[Mux.scala 31:69:@4074.4]
  assign _T_22538 = valid_12_53 ? 6'h35 : _T_22537; // @[Mux.scala 31:69:@4075.4]
  assign _T_22539 = valid_12_52 ? 6'h34 : _T_22538; // @[Mux.scala 31:69:@4076.4]
  assign _T_22540 = valid_12_51 ? 6'h33 : _T_22539; // @[Mux.scala 31:69:@4077.4]
  assign _T_22541 = valid_12_50 ? 6'h32 : _T_22540; // @[Mux.scala 31:69:@4078.4]
  assign _T_22542 = valid_12_49 ? 6'h31 : _T_22541; // @[Mux.scala 31:69:@4079.4]
  assign _T_22543 = valid_12_48 ? 6'h30 : _T_22542; // @[Mux.scala 31:69:@4080.4]
  assign _T_22544 = valid_12_47 ? 6'h2f : _T_22543; // @[Mux.scala 31:69:@4081.4]
  assign _T_22545 = valid_12_46 ? 6'h2e : _T_22544; // @[Mux.scala 31:69:@4082.4]
  assign _T_22546 = valid_12_45 ? 6'h2d : _T_22545; // @[Mux.scala 31:69:@4083.4]
  assign _T_22547 = valid_12_44 ? 6'h2c : _T_22546; // @[Mux.scala 31:69:@4084.4]
  assign _T_22548 = valid_12_43 ? 6'h2b : _T_22547; // @[Mux.scala 31:69:@4085.4]
  assign _T_22549 = valid_12_42 ? 6'h2a : _T_22548; // @[Mux.scala 31:69:@4086.4]
  assign _T_22550 = valid_12_41 ? 6'h29 : _T_22549; // @[Mux.scala 31:69:@4087.4]
  assign _T_22551 = valid_12_40 ? 6'h28 : _T_22550; // @[Mux.scala 31:69:@4088.4]
  assign _T_22552 = valid_12_39 ? 6'h27 : _T_22551; // @[Mux.scala 31:69:@4089.4]
  assign _T_22553 = valid_12_38 ? 6'h26 : _T_22552; // @[Mux.scala 31:69:@4090.4]
  assign _T_22554 = valid_12_37 ? 6'h25 : _T_22553; // @[Mux.scala 31:69:@4091.4]
  assign _T_22555 = valid_12_36 ? 6'h24 : _T_22554; // @[Mux.scala 31:69:@4092.4]
  assign _T_22556 = valid_12_35 ? 6'h23 : _T_22555; // @[Mux.scala 31:69:@4093.4]
  assign _T_22557 = valid_12_34 ? 6'h22 : _T_22556; // @[Mux.scala 31:69:@4094.4]
  assign _T_22558 = valid_12_33 ? 6'h21 : _T_22557; // @[Mux.scala 31:69:@4095.4]
  assign _T_22559 = valid_12_32 ? 6'h20 : _T_22558; // @[Mux.scala 31:69:@4096.4]
  assign _T_22560 = valid_12_31 ? 6'h1f : _T_22559; // @[Mux.scala 31:69:@4097.4]
  assign _T_22561 = valid_12_30 ? 6'h1e : _T_22560; // @[Mux.scala 31:69:@4098.4]
  assign _T_22562 = valid_12_29 ? 6'h1d : _T_22561; // @[Mux.scala 31:69:@4099.4]
  assign _T_22563 = valid_12_28 ? 6'h1c : _T_22562; // @[Mux.scala 31:69:@4100.4]
  assign _T_22564 = valid_12_27 ? 6'h1b : _T_22563; // @[Mux.scala 31:69:@4101.4]
  assign _T_22565 = valid_12_26 ? 6'h1a : _T_22564; // @[Mux.scala 31:69:@4102.4]
  assign _T_22566 = valid_12_25 ? 6'h19 : _T_22565; // @[Mux.scala 31:69:@4103.4]
  assign _T_22567 = valid_12_24 ? 6'h18 : _T_22566; // @[Mux.scala 31:69:@4104.4]
  assign _T_22568 = valid_12_23 ? 6'h17 : _T_22567; // @[Mux.scala 31:69:@4105.4]
  assign _T_22569 = valid_12_22 ? 6'h16 : _T_22568; // @[Mux.scala 31:69:@4106.4]
  assign _T_22570 = valid_12_21 ? 6'h15 : _T_22569; // @[Mux.scala 31:69:@4107.4]
  assign _T_22571 = valid_12_20 ? 6'h14 : _T_22570; // @[Mux.scala 31:69:@4108.4]
  assign _T_22572 = valid_12_19 ? 6'h13 : _T_22571; // @[Mux.scala 31:69:@4109.4]
  assign _T_22573 = valid_12_18 ? 6'h12 : _T_22572; // @[Mux.scala 31:69:@4110.4]
  assign _T_22574 = valid_12_17 ? 6'h11 : _T_22573; // @[Mux.scala 31:69:@4111.4]
  assign _T_22575 = valid_12_16 ? 6'h10 : _T_22574; // @[Mux.scala 31:69:@4112.4]
  assign _T_22576 = valid_12_15 ? 6'hf : _T_22575; // @[Mux.scala 31:69:@4113.4]
  assign _T_22577 = valid_12_14 ? 6'he : _T_22576; // @[Mux.scala 31:69:@4114.4]
  assign _T_22578 = valid_12_13 ? 6'hd : _T_22577; // @[Mux.scala 31:69:@4115.4]
  assign _T_22579 = valid_12_12 ? 6'hc : _T_22578; // @[Mux.scala 31:69:@4116.4]
  assign _T_22580 = valid_12_11 ? 6'hb : _T_22579; // @[Mux.scala 31:69:@4117.4]
  assign _T_22581 = valid_12_10 ? 6'ha : _T_22580; // @[Mux.scala 31:69:@4118.4]
  assign _T_22582 = valid_12_9 ? 6'h9 : _T_22581; // @[Mux.scala 31:69:@4119.4]
  assign _T_22583 = valid_12_8 ? 6'h8 : _T_22582; // @[Mux.scala 31:69:@4120.4]
  assign _T_22584 = valid_12_7 ? 6'h7 : _T_22583; // @[Mux.scala 31:69:@4121.4]
  assign _T_22585 = valid_12_6 ? 6'h6 : _T_22584; // @[Mux.scala 31:69:@4122.4]
  assign _T_22586 = valid_12_5 ? 6'h5 : _T_22585; // @[Mux.scala 31:69:@4123.4]
  assign _T_22587 = valid_12_4 ? 6'h4 : _T_22586; // @[Mux.scala 31:69:@4124.4]
  assign _T_22588 = valid_12_3 ? 6'h3 : _T_22587; // @[Mux.scala 31:69:@4125.4]
  assign _T_22589 = valid_12_2 ? 6'h2 : _T_22588; // @[Mux.scala 31:69:@4126.4]
  assign _T_22590 = valid_12_1 ? 6'h1 : _T_22589; // @[Mux.scala 31:69:@4127.4]
  assign select_12 = valid_12_0 ? 6'h0 : _T_22590; // @[Mux.scala 31:69:@4128.4]
  assign _GEN_769 = 6'h1 == select_12 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_770 = 6'h2 == select_12 ? io_inData_2 : _GEN_769; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_771 = 6'h3 == select_12 ? io_inData_3 : _GEN_770; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_772 = 6'h4 == select_12 ? io_inData_4 : _GEN_771; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_773 = 6'h5 == select_12 ? io_inData_5 : _GEN_772; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_774 = 6'h6 == select_12 ? io_inData_6 : _GEN_773; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_775 = 6'h7 == select_12 ? io_inData_7 : _GEN_774; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_776 = 6'h8 == select_12 ? io_inData_8 : _GEN_775; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_777 = 6'h9 == select_12 ? io_inData_9 : _GEN_776; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_778 = 6'ha == select_12 ? io_inData_10 : _GEN_777; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_779 = 6'hb == select_12 ? io_inData_11 : _GEN_778; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_780 = 6'hc == select_12 ? io_inData_12 : _GEN_779; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_781 = 6'hd == select_12 ? io_inData_13 : _GEN_780; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_782 = 6'he == select_12 ? io_inData_14 : _GEN_781; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_783 = 6'hf == select_12 ? io_inData_15 : _GEN_782; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_784 = 6'h10 == select_12 ? io_inData_16 : _GEN_783; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_785 = 6'h11 == select_12 ? io_inData_17 : _GEN_784; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_786 = 6'h12 == select_12 ? io_inData_18 : _GEN_785; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_787 = 6'h13 == select_12 ? io_inData_19 : _GEN_786; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_788 = 6'h14 == select_12 ? io_inData_20 : _GEN_787; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_789 = 6'h15 == select_12 ? io_inData_21 : _GEN_788; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_790 = 6'h16 == select_12 ? io_inData_22 : _GEN_789; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_791 = 6'h17 == select_12 ? io_inData_23 : _GEN_790; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_792 = 6'h18 == select_12 ? io_inData_24 : _GEN_791; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_793 = 6'h19 == select_12 ? io_inData_25 : _GEN_792; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_794 = 6'h1a == select_12 ? io_inData_26 : _GEN_793; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_795 = 6'h1b == select_12 ? io_inData_27 : _GEN_794; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_796 = 6'h1c == select_12 ? io_inData_28 : _GEN_795; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_797 = 6'h1d == select_12 ? io_inData_29 : _GEN_796; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_798 = 6'h1e == select_12 ? io_inData_30 : _GEN_797; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_799 = 6'h1f == select_12 ? io_inData_31 : _GEN_798; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_800 = 6'h20 == select_12 ? io_inData_32 : _GEN_799; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_801 = 6'h21 == select_12 ? io_inData_33 : _GEN_800; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_802 = 6'h22 == select_12 ? io_inData_34 : _GEN_801; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_803 = 6'h23 == select_12 ? io_inData_35 : _GEN_802; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_804 = 6'h24 == select_12 ? io_inData_36 : _GEN_803; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_805 = 6'h25 == select_12 ? io_inData_37 : _GEN_804; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_806 = 6'h26 == select_12 ? io_inData_38 : _GEN_805; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_807 = 6'h27 == select_12 ? io_inData_39 : _GEN_806; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_808 = 6'h28 == select_12 ? io_inData_40 : _GEN_807; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_809 = 6'h29 == select_12 ? io_inData_41 : _GEN_808; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_810 = 6'h2a == select_12 ? io_inData_42 : _GEN_809; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_811 = 6'h2b == select_12 ? io_inData_43 : _GEN_810; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_812 = 6'h2c == select_12 ? io_inData_44 : _GEN_811; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_813 = 6'h2d == select_12 ? io_inData_45 : _GEN_812; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_814 = 6'h2e == select_12 ? io_inData_46 : _GEN_813; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_815 = 6'h2f == select_12 ? io_inData_47 : _GEN_814; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_816 = 6'h30 == select_12 ? io_inData_48 : _GEN_815; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_817 = 6'h31 == select_12 ? io_inData_49 : _GEN_816; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_818 = 6'h32 == select_12 ? io_inData_50 : _GEN_817; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_819 = 6'h33 == select_12 ? io_inData_51 : _GEN_818; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_820 = 6'h34 == select_12 ? io_inData_52 : _GEN_819; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_821 = 6'h35 == select_12 ? io_inData_53 : _GEN_820; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_822 = 6'h36 == select_12 ? io_inData_54 : _GEN_821; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_823 = 6'h37 == select_12 ? io_inData_55 : _GEN_822; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_824 = 6'h38 == select_12 ? io_inData_56 : _GEN_823; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_825 = 6'h39 == select_12 ? io_inData_57 : _GEN_824; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_826 = 6'h3a == select_12 ? io_inData_58 : _GEN_825; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_827 = 6'h3b == select_12 ? io_inData_59 : _GEN_826; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_828 = 6'h3c == select_12 ? io_inData_60 : _GEN_827; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_829 = 6'h3d == select_12 ? io_inData_61 : _GEN_828; // @[Switch.scala 33:19:@4130.4]
  assign _GEN_830 = 6'h3e == select_12 ? io_inData_62 : _GEN_829; // @[Switch.scala 33:19:@4130.4]
  assign _T_22599 = {valid_12_7,valid_12_6,valid_12_5,valid_12_4,valid_12_3,valid_12_2,valid_12_1,valid_12_0}; // @[Switch.scala 34:32:@4137.4]
  assign _T_22607 = {valid_12_15,valid_12_14,valid_12_13,valid_12_12,valid_12_11,valid_12_10,valid_12_9,valid_12_8,_T_22599}; // @[Switch.scala 34:32:@4145.4]
  assign _T_22614 = {valid_12_23,valid_12_22,valid_12_21,valid_12_20,valid_12_19,valid_12_18,valid_12_17,valid_12_16}; // @[Switch.scala 34:32:@4152.4]
  assign _T_22623 = {valid_12_31,valid_12_30,valid_12_29,valid_12_28,valid_12_27,valid_12_26,valid_12_25,valid_12_24,_T_22614,_T_22607}; // @[Switch.scala 34:32:@4161.4]
  assign _T_22630 = {valid_12_39,valid_12_38,valid_12_37,valid_12_36,valid_12_35,valid_12_34,valid_12_33,valid_12_32}; // @[Switch.scala 34:32:@4168.4]
  assign _T_22638 = {valid_12_47,valid_12_46,valid_12_45,valid_12_44,valid_12_43,valid_12_42,valid_12_41,valid_12_40,_T_22630}; // @[Switch.scala 34:32:@4176.4]
  assign _T_22645 = {valid_12_55,valid_12_54,valid_12_53,valid_12_52,valid_12_51,valid_12_50,valid_12_49,valid_12_48}; // @[Switch.scala 34:32:@4183.4]
  assign _T_22654 = {valid_12_63,valid_12_62,valid_12_61,valid_12_60,valid_12_59,valid_12_58,valid_12_57,valid_12_56,_T_22645,_T_22638}; // @[Switch.scala 34:32:@4192.4]
  assign _T_22655 = {_T_22654,_T_22623}; // @[Switch.scala 34:32:@4193.4]
  assign _T_22659 = io_inAddr_0 == 6'hd; // @[Switch.scala 30:53:@4196.4]
  assign valid_13_0 = io_inValid_0 & _T_22659; // @[Switch.scala 30:36:@4197.4]
  assign _T_22662 = io_inAddr_1 == 6'hd; // @[Switch.scala 30:53:@4199.4]
  assign valid_13_1 = io_inValid_1 & _T_22662; // @[Switch.scala 30:36:@4200.4]
  assign _T_22665 = io_inAddr_2 == 6'hd; // @[Switch.scala 30:53:@4202.4]
  assign valid_13_2 = io_inValid_2 & _T_22665; // @[Switch.scala 30:36:@4203.4]
  assign _T_22668 = io_inAddr_3 == 6'hd; // @[Switch.scala 30:53:@4205.4]
  assign valid_13_3 = io_inValid_3 & _T_22668; // @[Switch.scala 30:36:@4206.4]
  assign _T_22671 = io_inAddr_4 == 6'hd; // @[Switch.scala 30:53:@4208.4]
  assign valid_13_4 = io_inValid_4 & _T_22671; // @[Switch.scala 30:36:@4209.4]
  assign _T_22674 = io_inAddr_5 == 6'hd; // @[Switch.scala 30:53:@4211.4]
  assign valid_13_5 = io_inValid_5 & _T_22674; // @[Switch.scala 30:36:@4212.4]
  assign _T_22677 = io_inAddr_6 == 6'hd; // @[Switch.scala 30:53:@4214.4]
  assign valid_13_6 = io_inValid_6 & _T_22677; // @[Switch.scala 30:36:@4215.4]
  assign _T_22680 = io_inAddr_7 == 6'hd; // @[Switch.scala 30:53:@4217.4]
  assign valid_13_7 = io_inValid_7 & _T_22680; // @[Switch.scala 30:36:@4218.4]
  assign _T_22683 = io_inAddr_8 == 6'hd; // @[Switch.scala 30:53:@4220.4]
  assign valid_13_8 = io_inValid_8 & _T_22683; // @[Switch.scala 30:36:@4221.4]
  assign _T_22686 = io_inAddr_9 == 6'hd; // @[Switch.scala 30:53:@4223.4]
  assign valid_13_9 = io_inValid_9 & _T_22686; // @[Switch.scala 30:36:@4224.4]
  assign _T_22689 = io_inAddr_10 == 6'hd; // @[Switch.scala 30:53:@4226.4]
  assign valid_13_10 = io_inValid_10 & _T_22689; // @[Switch.scala 30:36:@4227.4]
  assign _T_22692 = io_inAddr_11 == 6'hd; // @[Switch.scala 30:53:@4229.4]
  assign valid_13_11 = io_inValid_11 & _T_22692; // @[Switch.scala 30:36:@4230.4]
  assign _T_22695 = io_inAddr_12 == 6'hd; // @[Switch.scala 30:53:@4232.4]
  assign valid_13_12 = io_inValid_12 & _T_22695; // @[Switch.scala 30:36:@4233.4]
  assign _T_22698 = io_inAddr_13 == 6'hd; // @[Switch.scala 30:53:@4235.4]
  assign valid_13_13 = io_inValid_13 & _T_22698; // @[Switch.scala 30:36:@4236.4]
  assign _T_22701 = io_inAddr_14 == 6'hd; // @[Switch.scala 30:53:@4238.4]
  assign valid_13_14 = io_inValid_14 & _T_22701; // @[Switch.scala 30:36:@4239.4]
  assign _T_22704 = io_inAddr_15 == 6'hd; // @[Switch.scala 30:53:@4241.4]
  assign valid_13_15 = io_inValid_15 & _T_22704; // @[Switch.scala 30:36:@4242.4]
  assign _T_22707 = io_inAddr_16 == 6'hd; // @[Switch.scala 30:53:@4244.4]
  assign valid_13_16 = io_inValid_16 & _T_22707; // @[Switch.scala 30:36:@4245.4]
  assign _T_22710 = io_inAddr_17 == 6'hd; // @[Switch.scala 30:53:@4247.4]
  assign valid_13_17 = io_inValid_17 & _T_22710; // @[Switch.scala 30:36:@4248.4]
  assign _T_22713 = io_inAddr_18 == 6'hd; // @[Switch.scala 30:53:@4250.4]
  assign valid_13_18 = io_inValid_18 & _T_22713; // @[Switch.scala 30:36:@4251.4]
  assign _T_22716 = io_inAddr_19 == 6'hd; // @[Switch.scala 30:53:@4253.4]
  assign valid_13_19 = io_inValid_19 & _T_22716; // @[Switch.scala 30:36:@4254.4]
  assign _T_22719 = io_inAddr_20 == 6'hd; // @[Switch.scala 30:53:@4256.4]
  assign valid_13_20 = io_inValid_20 & _T_22719; // @[Switch.scala 30:36:@4257.4]
  assign _T_22722 = io_inAddr_21 == 6'hd; // @[Switch.scala 30:53:@4259.4]
  assign valid_13_21 = io_inValid_21 & _T_22722; // @[Switch.scala 30:36:@4260.4]
  assign _T_22725 = io_inAddr_22 == 6'hd; // @[Switch.scala 30:53:@4262.4]
  assign valid_13_22 = io_inValid_22 & _T_22725; // @[Switch.scala 30:36:@4263.4]
  assign _T_22728 = io_inAddr_23 == 6'hd; // @[Switch.scala 30:53:@4265.4]
  assign valid_13_23 = io_inValid_23 & _T_22728; // @[Switch.scala 30:36:@4266.4]
  assign _T_22731 = io_inAddr_24 == 6'hd; // @[Switch.scala 30:53:@4268.4]
  assign valid_13_24 = io_inValid_24 & _T_22731; // @[Switch.scala 30:36:@4269.4]
  assign _T_22734 = io_inAddr_25 == 6'hd; // @[Switch.scala 30:53:@4271.4]
  assign valid_13_25 = io_inValid_25 & _T_22734; // @[Switch.scala 30:36:@4272.4]
  assign _T_22737 = io_inAddr_26 == 6'hd; // @[Switch.scala 30:53:@4274.4]
  assign valid_13_26 = io_inValid_26 & _T_22737; // @[Switch.scala 30:36:@4275.4]
  assign _T_22740 = io_inAddr_27 == 6'hd; // @[Switch.scala 30:53:@4277.4]
  assign valid_13_27 = io_inValid_27 & _T_22740; // @[Switch.scala 30:36:@4278.4]
  assign _T_22743 = io_inAddr_28 == 6'hd; // @[Switch.scala 30:53:@4280.4]
  assign valid_13_28 = io_inValid_28 & _T_22743; // @[Switch.scala 30:36:@4281.4]
  assign _T_22746 = io_inAddr_29 == 6'hd; // @[Switch.scala 30:53:@4283.4]
  assign valid_13_29 = io_inValid_29 & _T_22746; // @[Switch.scala 30:36:@4284.4]
  assign _T_22749 = io_inAddr_30 == 6'hd; // @[Switch.scala 30:53:@4286.4]
  assign valid_13_30 = io_inValid_30 & _T_22749; // @[Switch.scala 30:36:@4287.4]
  assign _T_22752 = io_inAddr_31 == 6'hd; // @[Switch.scala 30:53:@4289.4]
  assign valid_13_31 = io_inValid_31 & _T_22752; // @[Switch.scala 30:36:@4290.4]
  assign _T_22755 = io_inAddr_32 == 6'hd; // @[Switch.scala 30:53:@4292.4]
  assign valid_13_32 = io_inValid_32 & _T_22755; // @[Switch.scala 30:36:@4293.4]
  assign _T_22758 = io_inAddr_33 == 6'hd; // @[Switch.scala 30:53:@4295.4]
  assign valid_13_33 = io_inValid_33 & _T_22758; // @[Switch.scala 30:36:@4296.4]
  assign _T_22761 = io_inAddr_34 == 6'hd; // @[Switch.scala 30:53:@4298.4]
  assign valid_13_34 = io_inValid_34 & _T_22761; // @[Switch.scala 30:36:@4299.4]
  assign _T_22764 = io_inAddr_35 == 6'hd; // @[Switch.scala 30:53:@4301.4]
  assign valid_13_35 = io_inValid_35 & _T_22764; // @[Switch.scala 30:36:@4302.4]
  assign _T_22767 = io_inAddr_36 == 6'hd; // @[Switch.scala 30:53:@4304.4]
  assign valid_13_36 = io_inValid_36 & _T_22767; // @[Switch.scala 30:36:@4305.4]
  assign _T_22770 = io_inAddr_37 == 6'hd; // @[Switch.scala 30:53:@4307.4]
  assign valid_13_37 = io_inValid_37 & _T_22770; // @[Switch.scala 30:36:@4308.4]
  assign _T_22773 = io_inAddr_38 == 6'hd; // @[Switch.scala 30:53:@4310.4]
  assign valid_13_38 = io_inValid_38 & _T_22773; // @[Switch.scala 30:36:@4311.4]
  assign _T_22776 = io_inAddr_39 == 6'hd; // @[Switch.scala 30:53:@4313.4]
  assign valid_13_39 = io_inValid_39 & _T_22776; // @[Switch.scala 30:36:@4314.4]
  assign _T_22779 = io_inAddr_40 == 6'hd; // @[Switch.scala 30:53:@4316.4]
  assign valid_13_40 = io_inValid_40 & _T_22779; // @[Switch.scala 30:36:@4317.4]
  assign _T_22782 = io_inAddr_41 == 6'hd; // @[Switch.scala 30:53:@4319.4]
  assign valid_13_41 = io_inValid_41 & _T_22782; // @[Switch.scala 30:36:@4320.4]
  assign _T_22785 = io_inAddr_42 == 6'hd; // @[Switch.scala 30:53:@4322.4]
  assign valid_13_42 = io_inValid_42 & _T_22785; // @[Switch.scala 30:36:@4323.4]
  assign _T_22788 = io_inAddr_43 == 6'hd; // @[Switch.scala 30:53:@4325.4]
  assign valid_13_43 = io_inValid_43 & _T_22788; // @[Switch.scala 30:36:@4326.4]
  assign _T_22791 = io_inAddr_44 == 6'hd; // @[Switch.scala 30:53:@4328.4]
  assign valid_13_44 = io_inValid_44 & _T_22791; // @[Switch.scala 30:36:@4329.4]
  assign _T_22794 = io_inAddr_45 == 6'hd; // @[Switch.scala 30:53:@4331.4]
  assign valid_13_45 = io_inValid_45 & _T_22794; // @[Switch.scala 30:36:@4332.4]
  assign _T_22797 = io_inAddr_46 == 6'hd; // @[Switch.scala 30:53:@4334.4]
  assign valid_13_46 = io_inValid_46 & _T_22797; // @[Switch.scala 30:36:@4335.4]
  assign _T_22800 = io_inAddr_47 == 6'hd; // @[Switch.scala 30:53:@4337.4]
  assign valid_13_47 = io_inValid_47 & _T_22800; // @[Switch.scala 30:36:@4338.4]
  assign _T_22803 = io_inAddr_48 == 6'hd; // @[Switch.scala 30:53:@4340.4]
  assign valid_13_48 = io_inValid_48 & _T_22803; // @[Switch.scala 30:36:@4341.4]
  assign _T_22806 = io_inAddr_49 == 6'hd; // @[Switch.scala 30:53:@4343.4]
  assign valid_13_49 = io_inValid_49 & _T_22806; // @[Switch.scala 30:36:@4344.4]
  assign _T_22809 = io_inAddr_50 == 6'hd; // @[Switch.scala 30:53:@4346.4]
  assign valid_13_50 = io_inValid_50 & _T_22809; // @[Switch.scala 30:36:@4347.4]
  assign _T_22812 = io_inAddr_51 == 6'hd; // @[Switch.scala 30:53:@4349.4]
  assign valid_13_51 = io_inValid_51 & _T_22812; // @[Switch.scala 30:36:@4350.4]
  assign _T_22815 = io_inAddr_52 == 6'hd; // @[Switch.scala 30:53:@4352.4]
  assign valid_13_52 = io_inValid_52 & _T_22815; // @[Switch.scala 30:36:@4353.4]
  assign _T_22818 = io_inAddr_53 == 6'hd; // @[Switch.scala 30:53:@4355.4]
  assign valid_13_53 = io_inValid_53 & _T_22818; // @[Switch.scala 30:36:@4356.4]
  assign _T_22821 = io_inAddr_54 == 6'hd; // @[Switch.scala 30:53:@4358.4]
  assign valid_13_54 = io_inValid_54 & _T_22821; // @[Switch.scala 30:36:@4359.4]
  assign _T_22824 = io_inAddr_55 == 6'hd; // @[Switch.scala 30:53:@4361.4]
  assign valid_13_55 = io_inValid_55 & _T_22824; // @[Switch.scala 30:36:@4362.4]
  assign _T_22827 = io_inAddr_56 == 6'hd; // @[Switch.scala 30:53:@4364.4]
  assign valid_13_56 = io_inValid_56 & _T_22827; // @[Switch.scala 30:36:@4365.4]
  assign _T_22830 = io_inAddr_57 == 6'hd; // @[Switch.scala 30:53:@4367.4]
  assign valid_13_57 = io_inValid_57 & _T_22830; // @[Switch.scala 30:36:@4368.4]
  assign _T_22833 = io_inAddr_58 == 6'hd; // @[Switch.scala 30:53:@4370.4]
  assign valid_13_58 = io_inValid_58 & _T_22833; // @[Switch.scala 30:36:@4371.4]
  assign _T_22836 = io_inAddr_59 == 6'hd; // @[Switch.scala 30:53:@4373.4]
  assign valid_13_59 = io_inValid_59 & _T_22836; // @[Switch.scala 30:36:@4374.4]
  assign _T_22839 = io_inAddr_60 == 6'hd; // @[Switch.scala 30:53:@4376.4]
  assign valid_13_60 = io_inValid_60 & _T_22839; // @[Switch.scala 30:36:@4377.4]
  assign _T_22842 = io_inAddr_61 == 6'hd; // @[Switch.scala 30:53:@4379.4]
  assign valid_13_61 = io_inValid_61 & _T_22842; // @[Switch.scala 30:36:@4380.4]
  assign _T_22845 = io_inAddr_62 == 6'hd; // @[Switch.scala 30:53:@4382.4]
  assign valid_13_62 = io_inValid_62 & _T_22845; // @[Switch.scala 30:36:@4383.4]
  assign _T_22848 = io_inAddr_63 == 6'hd; // @[Switch.scala 30:53:@4385.4]
  assign valid_13_63 = io_inValid_63 & _T_22848; // @[Switch.scala 30:36:@4386.4]
  assign _T_22914 = valid_13_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@4388.4]
  assign _T_22915 = valid_13_61 ? 6'h3d : _T_22914; // @[Mux.scala 31:69:@4389.4]
  assign _T_22916 = valid_13_60 ? 6'h3c : _T_22915; // @[Mux.scala 31:69:@4390.4]
  assign _T_22917 = valid_13_59 ? 6'h3b : _T_22916; // @[Mux.scala 31:69:@4391.4]
  assign _T_22918 = valid_13_58 ? 6'h3a : _T_22917; // @[Mux.scala 31:69:@4392.4]
  assign _T_22919 = valid_13_57 ? 6'h39 : _T_22918; // @[Mux.scala 31:69:@4393.4]
  assign _T_22920 = valid_13_56 ? 6'h38 : _T_22919; // @[Mux.scala 31:69:@4394.4]
  assign _T_22921 = valid_13_55 ? 6'h37 : _T_22920; // @[Mux.scala 31:69:@4395.4]
  assign _T_22922 = valid_13_54 ? 6'h36 : _T_22921; // @[Mux.scala 31:69:@4396.4]
  assign _T_22923 = valid_13_53 ? 6'h35 : _T_22922; // @[Mux.scala 31:69:@4397.4]
  assign _T_22924 = valid_13_52 ? 6'h34 : _T_22923; // @[Mux.scala 31:69:@4398.4]
  assign _T_22925 = valid_13_51 ? 6'h33 : _T_22924; // @[Mux.scala 31:69:@4399.4]
  assign _T_22926 = valid_13_50 ? 6'h32 : _T_22925; // @[Mux.scala 31:69:@4400.4]
  assign _T_22927 = valid_13_49 ? 6'h31 : _T_22926; // @[Mux.scala 31:69:@4401.4]
  assign _T_22928 = valid_13_48 ? 6'h30 : _T_22927; // @[Mux.scala 31:69:@4402.4]
  assign _T_22929 = valid_13_47 ? 6'h2f : _T_22928; // @[Mux.scala 31:69:@4403.4]
  assign _T_22930 = valid_13_46 ? 6'h2e : _T_22929; // @[Mux.scala 31:69:@4404.4]
  assign _T_22931 = valid_13_45 ? 6'h2d : _T_22930; // @[Mux.scala 31:69:@4405.4]
  assign _T_22932 = valid_13_44 ? 6'h2c : _T_22931; // @[Mux.scala 31:69:@4406.4]
  assign _T_22933 = valid_13_43 ? 6'h2b : _T_22932; // @[Mux.scala 31:69:@4407.4]
  assign _T_22934 = valid_13_42 ? 6'h2a : _T_22933; // @[Mux.scala 31:69:@4408.4]
  assign _T_22935 = valid_13_41 ? 6'h29 : _T_22934; // @[Mux.scala 31:69:@4409.4]
  assign _T_22936 = valid_13_40 ? 6'h28 : _T_22935; // @[Mux.scala 31:69:@4410.4]
  assign _T_22937 = valid_13_39 ? 6'h27 : _T_22936; // @[Mux.scala 31:69:@4411.4]
  assign _T_22938 = valid_13_38 ? 6'h26 : _T_22937; // @[Mux.scala 31:69:@4412.4]
  assign _T_22939 = valid_13_37 ? 6'h25 : _T_22938; // @[Mux.scala 31:69:@4413.4]
  assign _T_22940 = valid_13_36 ? 6'h24 : _T_22939; // @[Mux.scala 31:69:@4414.4]
  assign _T_22941 = valid_13_35 ? 6'h23 : _T_22940; // @[Mux.scala 31:69:@4415.4]
  assign _T_22942 = valid_13_34 ? 6'h22 : _T_22941; // @[Mux.scala 31:69:@4416.4]
  assign _T_22943 = valid_13_33 ? 6'h21 : _T_22942; // @[Mux.scala 31:69:@4417.4]
  assign _T_22944 = valid_13_32 ? 6'h20 : _T_22943; // @[Mux.scala 31:69:@4418.4]
  assign _T_22945 = valid_13_31 ? 6'h1f : _T_22944; // @[Mux.scala 31:69:@4419.4]
  assign _T_22946 = valid_13_30 ? 6'h1e : _T_22945; // @[Mux.scala 31:69:@4420.4]
  assign _T_22947 = valid_13_29 ? 6'h1d : _T_22946; // @[Mux.scala 31:69:@4421.4]
  assign _T_22948 = valid_13_28 ? 6'h1c : _T_22947; // @[Mux.scala 31:69:@4422.4]
  assign _T_22949 = valid_13_27 ? 6'h1b : _T_22948; // @[Mux.scala 31:69:@4423.4]
  assign _T_22950 = valid_13_26 ? 6'h1a : _T_22949; // @[Mux.scala 31:69:@4424.4]
  assign _T_22951 = valid_13_25 ? 6'h19 : _T_22950; // @[Mux.scala 31:69:@4425.4]
  assign _T_22952 = valid_13_24 ? 6'h18 : _T_22951; // @[Mux.scala 31:69:@4426.4]
  assign _T_22953 = valid_13_23 ? 6'h17 : _T_22952; // @[Mux.scala 31:69:@4427.4]
  assign _T_22954 = valid_13_22 ? 6'h16 : _T_22953; // @[Mux.scala 31:69:@4428.4]
  assign _T_22955 = valid_13_21 ? 6'h15 : _T_22954; // @[Mux.scala 31:69:@4429.4]
  assign _T_22956 = valid_13_20 ? 6'h14 : _T_22955; // @[Mux.scala 31:69:@4430.4]
  assign _T_22957 = valid_13_19 ? 6'h13 : _T_22956; // @[Mux.scala 31:69:@4431.4]
  assign _T_22958 = valid_13_18 ? 6'h12 : _T_22957; // @[Mux.scala 31:69:@4432.4]
  assign _T_22959 = valid_13_17 ? 6'h11 : _T_22958; // @[Mux.scala 31:69:@4433.4]
  assign _T_22960 = valid_13_16 ? 6'h10 : _T_22959; // @[Mux.scala 31:69:@4434.4]
  assign _T_22961 = valid_13_15 ? 6'hf : _T_22960; // @[Mux.scala 31:69:@4435.4]
  assign _T_22962 = valid_13_14 ? 6'he : _T_22961; // @[Mux.scala 31:69:@4436.4]
  assign _T_22963 = valid_13_13 ? 6'hd : _T_22962; // @[Mux.scala 31:69:@4437.4]
  assign _T_22964 = valid_13_12 ? 6'hc : _T_22963; // @[Mux.scala 31:69:@4438.4]
  assign _T_22965 = valid_13_11 ? 6'hb : _T_22964; // @[Mux.scala 31:69:@4439.4]
  assign _T_22966 = valid_13_10 ? 6'ha : _T_22965; // @[Mux.scala 31:69:@4440.4]
  assign _T_22967 = valid_13_9 ? 6'h9 : _T_22966; // @[Mux.scala 31:69:@4441.4]
  assign _T_22968 = valid_13_8 ? 6'h8 : _T_22967; // @[Mux.scala 31:69:@4442.4]
  assign _T_22969 = valid_13_7 ? 6'h7 : _T_22968; // @[Mux.scala 31:69:@4443.4]
  assign _T_22970 = valid_13_6 ? 6'h6 : _T_22969; // @[Mux.scala 31:69:@4444.4]
  assign _T_22971 = valid_13_5 ? 6'h5 : _T_22970; // @[Mux.scala 31:69:@4445.4]
  assign _T_22972 = valid_13_4 ? 6'h4 : _T_22971; // @[Mux.scala 31:69:@4446.4]
  assign _T_22973 = valid_13_3 ? 6'h3 : _T_22972; // @[Mux.scala 31:69:@4447.4]
  assign _T_22974 = valid_13_2 ? 6'h2 : _T_22973; // @[Mux.scala 31:69:@4448.4]
  assign _T_22975 = valid_13_1 ? 6'h1 : _T_22974; // @[Mux.scala 31:69:@4449.4]
  assign select_13 = valid_13_0 ? 6'h0 : _T_22975; // @[Mux.scala 31:69:@4450.4]
  assign _GEN_833 = 6'h1 == select_13 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_834 = 6'h2 == select_13 ? io_inData_2 : _GEN_833; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_835 = 6'h3 == select_13 ? io_inData_3 : _GEN_834; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_836 = 6'h4 == select_13 ? io_inData_4 : _GEN_835; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_837 = 6'h5 == select_13 ? io_inData_5 : _GEN_836; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_838 = 6'h6 == select_13 ? io_inData_6 : _GEN_837; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_839 = 6'h7 == select_13 ? io_inData_7 : _GEN_838; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_840 = 6'h8 == select_13 ? io_inData_8 : _GEN_839; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_841 = 6'h9 == select_13 ? io_inData_9 : _GEN_840; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_842 = 6'ha == select_13 ? io_inData_10 : _GEN_841; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_843 = 6'hb == select_13 ? io_inData_11 : _GEN_842; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_844 = 6'hc == select_13 ? io_inData_12 : _GEN_843; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_845 = 6'hd == select_13 ? io_inData_13 : _GEN_844; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_846 = 6'he == select_13 ? io_inData_14 : _GEN_845; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_847 = 6'hf == select_13 ? io_inData_15 : _GEN_846; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_848 = 6'h10 == select_13 ? io_inData_16 : _GEN_847; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_849 = 6'h11 == select_13 ? io_inData_17 : _GEN_848; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_850 = 6'h12 == select_13 ? io_inData_18 : _GEN_849; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_851 = 6'h13 == select_13 ? io_inData_19 : _GEN_850; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_852 = 6'h14 == select_13 ? io_inData_20 : _GEN_851; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_853 = 6'h15 == select_13 ? io_inData_21 : _GEN_852; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_854 = 6'h16 == select_13 ? io_inData_22 : _GEN_853; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_855 = 6'h17 == select_13 ? io_inData_23 : _GEN_854; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_856 = 6'h18 == select_13 ? io_inData_24 : _GEN_855; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_857 = 6'h19 == select_13 ? io_inData_25 : _GEN_856; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_858 = 6'h1a == select_13 ? io_inData_26 : _GEN_857; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_859 = 6'h1b == select_13 ? io_inData_27 : _GEN_858; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_860 = 6'h1c == select_13 ? io_inData_28 : _GEN_859; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_861 = 6'h1d == select_13 ? io_inData_29 : _GEN_860; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_862 = 6'h1e == select_13 ? io_inData_30 : _GEN_861; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_863 = 6'h1f == select_13 ? io_inData_31 : _GEN_862; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_864 = 6'h20 == select_13 ? io_inData_32 : _GEN_863; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_865 = 6'h21 == select_13 ? io_inData_33 : _GEN_864; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_866 = 6'h22 == select_13 ? io_inData_34 : _GEN_865; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_867 = 6'h23 == select_13 ? io_inData_35 : _GEN_866; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_868 = 6'h24 == select_13 ? io_inData_36 : _GEN_867; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_869 = 6'h25 == select_13 ? io_inData_37 : _GEN_868; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_870 = 6'h26 == select_13 ? io_inData_38 : _GEN_869; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_871 = 6'h27 == select_13 ? io_inData_39 : _GEN_870; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_872 = 6'h28 == select_13 ? io_inData_40 : _GEN_871; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_873 = 6'h29 == select_13 ? io_inData_41 : _GEN_872; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_874 = 6'h2a == select_13 ? io_inData_42 : _GEN_873; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_875 = 6'h2b == select_13 ? io_inData_43 : _GEN_874; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_876 = 6'h2c == select_13 ? io_inData_44 : _GEN_875; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_877 = 6'h2d == select_13 ? io_inData_45 : _GEN_876; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_878 = 6'h2e == select_13 ? io_inData_46 : _GEN_877; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_879 = 6'h2f == select_13 ? io_inData_47 : _GEN_878; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_880 = 6'h30 == select_13 ? io_inData_48 : _GEN_879; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_881 = 6'h31 == select_13 ? io_inData_49 : _GEN_880; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_882 = 6'h32 == select_13 ? io_inData_50 : _GEN_881; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_883 = 6'h33 == select_13 ? io_inData_51 : _GEN_882; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_884 = 6'h34 == select_13 ? io_inData_52 : _GEN_883; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_885 = 6'h35 == select_13 ? io_inData_53 : _GEN_884; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_886 = 6'h36 == select_13 ? io_inData_54 : _GEN_885; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_887 = 6'h37 == select_13 ? io_inData_55 : _GEN_886; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_888 = 6'h38 == select_13 ? io_inData_56 : _GEN_887; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_889 = 6'h39 == select_13 ? io_inData_57 : _GEN_888; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_890 = 6'h3a == select_13 ? io_inData_58 : _GEN_889; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_891 = 6'h3b == select_13 ? io_inData_59 : _GEN_890; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_892 = 6'h3c == select_13 ? io_inData_60 : _GEN_891; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_893 = 6'h3d == select_13 ? io_inData_61 : _GEN_892; // @[Switch.scala 33:19:@4452.4]
  assign _GEN_894 = 6'h3e == select_13 ? io_inData_62 : _GEN_893; // @[Switch.scala 33:19:@4452.4]
  assign _T_22984 = {valid_13_7,valid_13_6,valid_13_5,valid_13_4,valid_13_3,valid_13_2,valid_13_1,valid_13_0}; // @[Switch.scala 34:32:@4459.4]
  assign _T_22992 = {valid_13_15,valid_13_14,valid_13_13,valid_13_12,valid_13_11,valid_13_10,valid_13_9,valid_13_8,_T_22984}; // @[Switch.scala 34:32:@4467.4]
  assign _T_22999 = {valid_13_23,valid_13_22,valid_13_21,valid_13_20,valid_13_19,valid_13_18,valid_13_17,valid_13_16}; // @[Switch.scala 34:32:@4474.4]
  assign _T_23008 = {valid_13_31,valid_13_30,valid_13_29,valid_13_28,valid_13_27,valid_13_26,valid_13_25,valid_13_24,_T_22999,_T_22992}; // @[Switch.scala 34:32:@4483.4]
  assign _T_23015 = {valid_13_39,valid_13_38,valid_13_37,valid_13_36,valid_13_35,valid_13_34,valid_13_33,valid_13_32}; // @[Switch.scala 34:32:@4490.4]
  assign _T_23023 = {valid_13_47,valid_13_46,valid_13_45,valid_13_44,valid_13_43,valid_13_42,valid_13_41,valid_13_40,_T_23015}; // @[Switch.scala 34:32:@4498.4]
  assign _T_23030 = {valid_13_55,valid_13_54,valid_13_53,valid_13_52,valid_13_51,valid_13_50,valid_13_49,valid_13_48}; // @[Switch.scala 34:32:@4505.4]
  assign _T_23039 = {valid_13_63,valid_13_62,valid_13_61,valid_13_60,valid_13_59,valid_13_58,valid_13_57,valid_13_56,_T_23030,_T_23023}; // @[Switch.scala 34:32:@4514.4]
  assign _T_23040 = {_T_23039,_T_23008}; // @[Switch.scala 34:32:@4515.4]
  assign _T_23044 = io_inAddr_0 == 6'he; // @[Switch.scala 30:53:@4518.4]
  assign valid_14_0 = io_inValid_0 & _T_23044; // @[Switch.scala 30:36:@4519.4]
  assign _T_23047 = io_inAddr_1 == 6'he; // @[Switch.scala 30:53:@4521.4]
  assign valid_14_1 = io_inValid_1 & _T_23047; // @[Switch.scala 30:36:@4522.4]
  assign _T_23050 = io_inAddr_2 == 6'he; // @[Switch.scala 30:53:@4524.4]
  assign valid_14_2 = io_inValid_2 & _T_23050; // @[Switch.scala 30:36:@4525.4]
  assign _T_23053 = io_inAddr_3 == 6'he; // @[Switch.scala 30:53:@4527.4]
  assign valid_14_3 = io_inValid_3 & _T_23053; // @[Switch.scala 30:36:@4528.4]
  assign _T_23056 = io_inAddr_4 == 6'he; // @[Switch.scala 30:53:@4530.4]
  assign valid_14_4 = io_inValid_4 & _T_23056; // @[Switch.scala 30:36:@4531.4]
  assign _T_23059 = io_inAddr_5 == 6'he; // @[Switch.scala 30:53:@4533.4]
  assign valid_14_5 = io_inValid_5 & _T_23059; // @[Switch.scala 30:36:@4534.4]
  assign _T_23062 = io_inAddr_6 == 6'he; // @[Switch.scala 30:53:@4536.4]
  assign valid_14_6 = io_inValid_6 & _T_23062; // @[Switch.scala 30:36:@4537.4]
  assign _T_23065 = io_inAddr_7 == 6'he; // @[Switch.scala 30:53:@4539.4]
  assign valid_14_7 = io_inValid_7 & _T_23065; // @[Switch.scala 30:36:@4540.4]
  assign _T_23068 = io_inAddr_8 == 6'he; // @[Switch.scala 30:53:@4542.4]
  assign valid_14_8 = io_inValid_8 & _T_23068; // @[Switch.scala 30:36:@4543.4]
  assign _T_23071 = io_inAddr_9 == 6'he; // @[Switch.scala 30:53:@4545.4]
  assign valid_14_9 = io_inValid_9 & _T_23071; // @[Switch.scala 30:36:@4546.4]
  assign _T_23074 = io_inAddr_10 == 6'he; // @[Switch.scala 30:53:@4548.4]
  assign valid_14_10 = io_inValid_10 & _T_23074; // @[Switch.scala 30:36:@4549.4]
  assign _T_23077 = io_inAddr_11 == 6'he; // @[Switch.scala 30:53:@4551.4]
  assign valid_14_11 = io_inValid_11 & _T_23077; // @[Switch.scala 30:36:@4552.4]
  assign _T_23080 = io_inAddr_12 == 6'he; // @[Switch.scala 30:53:@4554.4]
  assign valid_14_12 = io_inValid_12 & _T_23080; // @[Switch.scala 30:36:@4555.4]
  assign _T_23083 = io_inAddr_13 == 6'he; // @[Switch.scala 30:53:@4557.4]
  assign valid_14_13 = io_inValid_13 & _T_23083; // @[Switch.scala 30:36:@4558.4]
  assign _T_23086 = io_inAddr_14 == 6'he; // @[Switch.scala 30:53:@4560.4]
  assign valid_14_14 = io_inValid_14 & _T_23086; // @[Switch.scala 30:36:@4561.4]
  assign _T_23089 = io_inAddr_15 == 6'he; // @[Switch.scala 30:53:@4563.4]
  assign valid_14_15 = io_inValid_15 & _T_23089; // @[Switch.scala 30:36:@4564.4]
  assign _T_23092 = io_inAddr_16 == 6'he; // @[Switch.scala 30:53:@4566.4]
  assign valid_14_16 = io_inValid_16 & _T_23092; // @[Switch.scala 30:36:@4567.4]
  assign _T_23095 = io_inAddr_17 == 6'he; // @[Switch.scala 30:53:@4569.4]
  assign valid_14_17 = io_inValid_17 & _T_23095; // @[Switch.scala 30:36:@4570.4]
  assign _T_23098 = io_inAddr_18 == 6'he; // @[Switch.scala 30:53:@4572.4]
  assign valid_14_18 = io_inValid_18 & _T_23098; // @[Switch.scala 30:36:@4573.4]
  assign _T_23101 = io_inAddr_19 == 6'he; // @[Switch.scala 30:53:@4575.4]
  assign valid_14_19 = io_inValid_19 & _T_23101; // @[Switch.scala 30:36:@4576.4]
  assign _T_23104 = io_inAddr_20 == 6'he; // @[Switch.scala 30:53:@4578.4]
  assign valid_14_20 = io_inValid_20 & _T_23104; // @[Switch.scala 30:36:@4579.4]
  assign _T_23107 = io_inAddr_21 == 6'he; // @[Switch.scala 30:53:@4581.4]
  assign valid_14_21 = io_inValid_21 & _T_23107; // @[Switch.scala 30:36:@4582.4]
  assign _T_23110 = io_inAddr_22 == 6'he; // @[Switch.scala 30:53:@4584.4]
  assign valid_14_22 = io_inValid_22 & _T_23110; // @[Switch.scala 30:36:@4585.4]
  assign _T_23113 = io_inAddr_23 == 6'he; // @[Switch.scala 30:53:@4587.4]
  assign valid_14_23 = io_inValid_23 & _T_23113; // @[Switch.scala 30:36:@4588.4]
  assign _T_23116 = io_inAddr_24 == 6'he; // @[Switch.scala 30:53:@4590.4]
  assign valid_14_24 = io_inValid_24 & _T_23116; // @[Switch.scala 30:36:@4591.4]
  assign _T_23119 = io_inAddr_25 == 6'he; // @[Switch.scala 30:53:@4593.4]
  assign valid_14_25 = io_inValid_25 & _T_23119; // @[Switch.scala 30:36:@4594.4]
  assign _T_23122 = io_inAddr_26 == 6'he; // @[Switch.scala 30:53:@4596.4]
  assign valid_14_26 = io_inValid_26 & _T_23122; // @[Switch.scala 30:36:@4597.4]
  assign _T_23125 = io_inAddr_27 == 6'he; // @[Switch.scala 30:53:@4599.4]
  assign valid_14_27 = io_inValid_27 & _T_23125; // @[Switch.scala 30:36:@4600.4]
  assign _T_23128 = io_inAddr_28 == 6'he; // @[Switch.scala 30:53:@4602.4]
  assign valid_14_28 = io_inValid_28 & _T_23128; // @[Switch.scala 30:36:@4603.4]
  assign _T_23131 = io_inAddr_29 == 6'he; // @[Switch.scala 30:53:@4605.4]
  assign valid_14_29 = io_inValid_29 & _T_23131; // @[Switch.scala 30:36:@4606.4]
  assign _T_23134 = io_inAddr_30 == 6'he; // @[Switch.scala 30:53:@4608.4]
  assign valid_14_30 = io_inValid_30 & _T_23134; // @[Switch.scala 30:36:@4609.4]
  assign _T_23137 = io_inAddr_31 == 6'he; // @[Switch.scala 30:53:@4611.4]
  assign valid_14_31 = io_inValid_31 & _T_23137; // @[Switch.scala 30:36:@4612.4]
  assign _T_23140 = io_inAddr_32 == 6'he; // @[Switch.scala 30:53:@4614.4]
  assign valid_14_32 = io_inValid_32 & _T_23140; // @[Switch.scala 30:36:@4615.4]
  assign _T_23143 = io_inAddr_33 == 6'he; // @[Switch.scala 30:53:@4617.4]
  assign valid_14_33 = io_inValid_33 & _T_23143; // @[Switch.scala 30:36:@4618.4]
  assign _T_23146 = io_inAddr_34 == 6'he; // @[Switch.scala 30:53:@4620.4]
  assign valid_14_34 = io_inValid_34 & _T_23146; // @[Switch.scala 30:36:@4621.4]
  assign _T_23149 = io_inAddr_35 == 6'he; // @[Switch.scala 30:53:@4623.4]
  assign valid_14_35 = io_inValid_35 & _T_23149; // @[Switch.scala 30:36:@4624.4]
  assign _T_23152 = io_inAddr_36 == 6'he; // @[Switch.scala 30:53:@4626.4]
  assign valid_14_36 = io_inValid_36 & _T_23152; // @[Switch.scala 30:36:@4627.4]
  assign _T_23155 = io_inAddr_37 == 6'he; // @[Switch.scala 30:53:@4629.4]
  assign valid_14_37 = io_inValid_37 & _T_23155; // @[Switch.scala 30:36:@4630.4]
  assign _T_23158 = io_inAddr_38 == 6'he; // @[Switch.scala 30:53:@4632.4]
  assign valid_14_38 = io_inValid_38 & _T_23158; // @[Switch.scala 30:36:@4633.4]
  assign _T_23161 = io_inAddr_39 == 6'he; // @[Switch.scala 30:53:@4635.4]
  assign valid_14_39 = io_inValid_39 & _T_23161; // @[Switch.scala 30:36:@4636.4]
  assign _T_23164 = io_inAddr_40 == 6'he; // @[Switch.scala 30:53:@4638.4]
  assign valid_14_40 = io_inValid_40 & _T_23164; // @[Switch.scala 30:36:@4639.4]
  assign _T_23167 = io_inAddr_41 == 6'he; // @[Switch.scala 30:53:@4641.4]
  assign valid_14_41 = io_inValid_41 & _T_23167; // @[Switch.scala 30:36:@4642.4]
  assign _T_23170 = io_inAddr_42 == 6'he; // @[Switch.scala 30:53:@4644.4]
  assign valid_14_42 = io_inValid_42 & _T_23170; // @[Switch.scala 30:36:@4645.4]
  assign _T_23173 = io_inAddr_43 == 6'he; // @[Switch.scala 30:53:@4647.4]
  assign valid_14_43 = io_inValid_43 & _T_23173; // @[Switch.scala 30:36:@4648.4]
  assign _T_23176 = io_inAddr_44 == 6'he; // @[Switch.scala 30:53:@4650.4]
  assign valid_14_44 = io_inValid_44 & _T_23176; // @[Switch.scala 30:36:@4651.4]
  assign _T_23179 = io_inAddr_45 == 6'he; // @[Switch.scala 30:53:@4653.4]
  assign valid_14_45 = io_inValid_45 & _T_23179; // @[Switch.scala 30:36:@4654.4]
  assign _T_23182 = io_inAddr_46 == 6'he; // @[Switch.scala 30:53:@4656.4]
  assign valid_14_46 = io_inValid_46 & _T_23182; // @[Switch.scala 30:36:@4657.4]
  assign _T_23185 = io_inAddr_47 == 6'he; // @[Switch.scala 30:53:@4659.4]
  assign valid_14_47 = io_inValid_47 & _T_23185; // @[Switch.scala 30:36:@4660.4]
  assign _T_23188 = io_inAddr_48 == 6'he; // @[Switch.scala 30:53:@4662.4]
  assign valid_14_48 = io_inValid_48 & _T_23188; // @[Switch.scala 30:36:@4663.4]
  assign _T_23191 = io_inAddr_49 == 6'he; // @[Switch.scala 30:53:@4665.4]
  assign valid_14_49 = io_inValid_49 & _T_23191; // @[Switch.scala 30:36:@4666.4]
  assign _T_23194 = io_inAddr_50 == 6'he; // @[Switch.scala 30:53:@4668.4]
  assign valid_14_50 = io_inValid_50 & _T_23194; // @[Switch.scala 30:36:@4669.4]
  assign _T_23197 = io_inAddr_51 == 6'he; // @[Switch.scala 30:53:@4671.4]
  assign valid_14_51 = io_inValid_51 & _T_23197; // @[Switch.scala 30:36:@4672.4]
  assign _T_23200 = io_inAddr_52 == 6'he; // @[Switch.scala 30:53:@4674.4]
  assign valid_14_52 = io_inValid_52 & _T_23200; // @[Switch.scala 30:36:@4675.4]
  assign _T_23203 = io_inAddr_53 == 6'he; // @[Switch.scala 30:53:@4677.4]
  assign valid_14_53 = io_inValid_53 & _T_23203; // @[Switch.scala 30:36:@4678.4]
  assign _T_23206 = io_inAddr_54 == 6'he; // @[Switch.scala 30:53:@4680.4]
  assign valid_14_54 = io_inValid_54 & _T_23206; // @[Switch.scala 30:36:@4681.4]
  assign _T_23209 = io_inAddr_55 == 6'he; // @[Switch.scala 30:53:@4683.4]
  assign valid_14_55 = io_inValid_55 & _T_23209; // @[Switch.scala 30:36:@4684.4]
  assign _T_23212 = io_inAddr_56 == 6'he; // @[Switch.scala 30:53:@4686.4]
  assign valid_14_56 = io_inValid_56 & _T_23212; // @[Switch.scala 30:36:@4687.4]
  assign _T_23215 = io_inAddr_57 == 6'he; // @[Switch.scala 30:53:@4689.4]
  assign valid_14_57 = io_inValid_57 & _T_23215; // @[Switch.scala 30:36:@4690.4]
  assign _T_23218 = io_inAddr_58 == 6'he; // @[Switch.scala 30:53:@4692.4]
  assign valid_14_58 = io_inValid_58 & _T_23218; // @[Switch.scala 30:36:@4693.4]
  assign _T_23221 = io_inAddr_59 == 6'he; // @[Switch.scala 30:53:@4695.4]
  assign valid_14_59 = io_inValid_59 & _T_23221; // @[Switch.scala 30:36:@4696.4]
  assign _T_23224 = io_inAddr_60 == 6'he; // @[Switch.scala 30:53:@4698.4]
  assign valid_14_60 = io_inValid_60 & _T_23224; // @[Switch.scala 30:36:@4699.4]
  assign _T_23227 = io_inAddr_61 == 6'he; // @[Switch.scala 30:53:@4701.4]
  assign valid_14_61 = io_inValid_61 & _T_23227; // @[Switch.scala 30:36:@4702.4]
  assign _T_23230 = io_inAddr_62 == 6'he; // @[Switch.scala 30:53:@4704.4]
  assign valid_14_62 = io_inValid_62 & _T_23230; // @[Switch.scala 30:36:@4705.4]
  assign _T_23233 = io_inAddr_63 == 6'he; // @[Switch.scala 30:53:@4707.4]
  assign valid_14_63 = io_inValid_63 & _T_23233; // @[Switch.scala 30:36:@4708.4]
  assign _T_23299 = valid_14_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@4710.4]
  assign _T_23300 = valid_14_61 ? 6'h3d : _T_23299; // @[Mux.scala 31:69:@4711.4]
  assign _T_23301 = valid_14_60 ? 6'h3c : _T_23300; // @[Mux.scala 31:69:@4712.4]
  assign _T_23302 = valid_14_59 ? 6'h3b : _T_23301; // @[Mux.scala 31:69:@4713.4]
  assign _T_23303 = valid_14_58 ? 6'h3a : _T_23302; // @[Mux.scala 31:69:@4714.4]
  assign _T_23304 = valid_14_57 ? 6'h39 : _T_23303; // @[Mux.scala 31:69:@4715.4]
  assign _T_23305 = valid_14_56 ? 6'h38 : _T_23304; // @[Mux.scala 31:69:@4716.4]
  assign _T_23306 = valid_14_55 ? 6'h37 : _T_23305; // @[Mux.scala 31:69:@4717.4]
  assign _T_23307 = valid_14_54 ? 6'h36 : _T_23306; // @[Mux.scala 31:69:@4718.4]
  assign _T_23308 = valid_14_53 ? 6'h35 : _T_23307; // @[Mux.scala 31:69:@4719.4]
  assign _T_23309 = valid_14_52 ? 6'h34 : _T_23308; // @[Mux.scala 31:69:@4720.4]
  assign _T_23310 = valid_14_51 ? 6'h33 : _T_23309; // @[Mux.scala 31:69:@4721.4]
  assign _T_23311 = valid_14_50 ? 6'h32 : _T_23310; // @[Mux.scala 31:69:@4722.4]
  assign _T_23312 = valid_14_49 ? 6'h31 : _T_23311; // @[Mux.scala 31:69:@4723.4]
  assign _T_23313 = valid_14_48 ? 6'h30 : _T_23312; // @[Mux.scala 31:69:@4724.4]
  assign _T_23314 = valid_14_47 ? 6'h2f : _T_23313; // @[Mux.scala 31:69:@4725.4]
  assign _T_23315 = valid_14_46 ? 6'h2e : _T_23314; // @[Mux.scala 31:69:@4726.4]
  assign _T_23316 = valid_14_45 ? 6'h2d : _T_23315; // @[Mux.scala 31:69:@4727.4]
  assign _T_23317 = valid_14_44 ? 6'h2c : _T_23316; // @[Mux.scala 31:69:@4728.4]
  assign _T_23318 = valid_14_43 ? 6'h2b : _T_23317; // @[Mux.scala 31:69:@4729.4]
  assign _T_23319 = valid_14_42 ? 6'h2a : _T_23318; // @[Mux.scala 31:69:@4730.4]
  assign _T_23320 = valid_14_41 ? 6'h29 : _T_23319; // @[Mux.scala 31:69:@4731.4]
  assign _T_23321 = valid_14_40 ? 6'h28 : _T_23320; // @[Mux.scala 31:69:@4732.4]
  assign _T_23322 = valid_14_39 ? 6'h27 : _T_23321; // @[Mux.scala 31:69:@4733.4]
  assign _T_23323 = valid_14_38 ? 6'h26 : _T_23322; // @[Mux.scala 31:69:@4734.4]
  assign _T_23324 = valid_14_37 ? 6'h25 : _T_23323; // @[Mux.scala 31:69:@4735.4]
  assign _T_23325 = valid_14_36 ? 6'h24 : _T_23324; // @[Mux.scala 31:69:@4736.4]
  assign _T_23326 = valid_14_35 ? 6'h23 : _T_23325; // @[Mux.scala 31:69:@4737.4]
  assign _T_23327 = valid_14_34 ? 6'h22 : _T_23326; // @[Mux.scala 31:69:@4738.4]
  assign _T_23328 = valid_14_33 ? 6'h21 : _T_23327; // @[Mux.scala 31:69:@4739.4]
  assign _T_23329 = valid_14_32 ? 6'h20 : _T_23328; // @[Mux.scala 31:69:@4740.4]
  assign _T_23330 = valid_14_31 ? 6'h1f : _T_23329; // @[Mux.scala 31:69:@4741.4]
  assign _T_23331 = valid_14_30 ? 6'h1e : _T_23330; // @[Mux.scala 31:69:@4742.4]
  assign _T_23332 = valid_14_29 ? 6'h1d : _T_23331; // @[Mux.scala 31:69:@4743.4]
  assign _T_23333 = valid_14_28 ? 6'h1c : _T_23332; // @[Mux.scala 31:69:@4744.4]
  assign _T_23334 = valid_14_27 ? 6'h1b : _T_23333; // @[Mux.scala 31:69:@4745.4]
  assign _T_23335 = valid_14_26 ? 6'h1a : _T_23334; // @[Mux.scala 31:69:@4746.4]
  assign _T_23336 = valid_14_25 ? 6'h19 : _T_23335; // @[Mux.scala 31:69:@4747.4]
  assign _T_23337 = valid_14_24 ? 6'h18 : _T_23336; // @[Mux.scala 31:69:@4748.4]
  assign _T_23338 = valid_14_23 ? 6'h17 : _T_23337; // @[Mux.scala 31:69:@4749.4]
  assign _T_23339 = valid_14_22 ? 6'h16 : _T_23338; // @[Mux.scala 31:69:@4750.4]
  assign _T_23340 = valid_14_21 ? 6'h15 : _T_23339; // @[Mux.scala 31:69:@4751.4]
  assign _T_23341 = valid_14_20 ? 6'h14 : _T_23340; // @[Mux.scala 31:69:@4752.4]
  assign _T_23342 = valid_14_19 ? 6'h13 : _T_23341; // @[Mux.scala 31:69:@4753.4]
  assign _T_23343 = valid_14_18 ? 6'h12 : _T_23342; // @[Mux.scala 31:69:@4754.4]
  assign _T_23344 = valid_14_17 ? 6'h11 : _T_23343; // @[Mux.scala 31:69:@4755.4]
  assign _T_23345 = valid_14_16 ? 6'h10 : _T_23344; // @[Mux.scala 31:69:@4756.4]
  assign _T_23346 = valid_14_15 ? 6'hf : _T_23345; // @[Mux.scala 31:69:@4757.4]
  assign _T_23347 = valid_14_14 ? 6'he : _T_23346; // @[Mux.scala 31:69:@4758.4]
  assign _T_23348 = valid_14_13 ? 6'hd : _T_23347; // @[Mux.scala 31:69:@4759.4]
  assign _T_23349 = valid_14_12 ? 6'hc : _T_23348; // @[Mux.scala 31:69:@4760.4]
  assign _T_23350 = valid_14_11 ? 6'hb : _T_23349; // @[Mux.scala 31:69:@4761.4]
  assign _T_23351 = valid_14_10 ? 6'ha : _T_23350; // @[Mux.scala 31:69:@4762.4]
  assign _T_23352 = valid_14_9 ? 6'h9 : _T_23351; // @[Mux.scala 31:69:@4763.4]
  assign _T_23353 = valid_14_8 ? 6'h8 : _T_23352; // @[Mux.scala 31:69:@4764.4]
  assign _T_23354 = valid_14_7 ? 6'h7 : _T_23353; // @[Mux.scala 31:69:@4765.4]
  assign _T_23355 = valid_14_6 ? 6'h6 : _T_23354; // @[Mux.scala 31:69:@4766.4]
  assign _T_23356 = valid_14_5 ? 6'h5 : _T_23355; // @[Mux.scala 31:69:@4767.4]
  assign _T_23357 = valid_14_4 ? 6'h4 : _T_23356; // @[Mux.scala 31:69:@4768.4]
  assign _T_23358 = valid_14_3 ? 6'h3 : _T_23357; // @[Mux.scala 31:69:@4769.4]
  assign _T_23359 = valid_14_2 ? 6'h2 : _T_23358; // @[Mux.scala 31:69:@4770.4]
  assign _T_23360 = valid_14_1 ? 6'h1 : _T_23359; // @[Mux.scala 31:69:@4771.4]
  assign select_14 = valid_14_0 ? 6'h0 : _T_23360; // @[Mux.scala 31:69:@4772.4]
  assign _GEN_897 = 6'h1 == select_14 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_898 = 6'h2 == select_14 ? io_inData_2 : _GEN_897; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_899 = 6'h3 == select_14 ? io_inData_3 : _GEN_898; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_900 = 6'h4 == select_14 ? io_inData_4 : _GEN_899; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_901 = 6'h5 == select_14 ? io_inData_5 : _GEN_900; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_902 = 6'h6 == select_14 ? io_inData_6 : _GEN_901; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_903 = 6'h7 == select_14 ? io_inData_7 : _GEN_902; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_904 = 6'h8 == select_14 ? io_inData_8 : _GEN_903; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_905 = 6'h9 == select_14 ? io_inData_9 : _GEN_904; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_906 = 6'ha == select_14 ? io_inData_10 : _GEN_905; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_907 = 6'hb == select_14 ? io_inData_11 : _GEN_906; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_908 = 6'hc == select_14 ? io_inData_12 : _GEN_907; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_909 = 6'hd == select_14 ? io_inData_13 : _GEN_908; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_910 = 6'he == select_14 ? io_inData_14 : _GEN_909; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_911 = 6'hf == select_14 ? io_inData_15 : _GEN_910; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_912 = 6'h10 == select_14 ? io_inData_16 : _GEN_911; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_913 = 6'h11 == select_14 ? io_inData_17 : _GEN_912; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_914 = 6'h12 == select_14 ? io_inData_18 : _GEN_913; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_915 = 6'h13 == select_14 ? io_inData_19 : _GEN_914; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_916 = 6'h14 == select_14 ? io_inData_20 : _GEN_915; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_917 = 6'h15 == select_14 ? io_inData_21 : _GEN_916; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_918 = 6'h16 == select_14 ? io_inData_22 : _GEN_917; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_919 = 6'h17 == select_14 ? io_inData_23 : _GEN_918; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_920 = 6'h18 == select_14 ? io_inData_24 : _GEN_919; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_921 = 6'h19 == select_14 ? io_inData_25 : _GEN_920; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_922 = 6'h1a == select_14 ? io_inData_26 : _GEN_921; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_923 = 6'h1b == select_14 ? io_inData_27 : _GEN_922; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_924 = 6'h1c == select_14 ? io_inData_28 : _GEN_923; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_925 = 6'h1d == select_14 ? io_inData_29 : _GEN_924; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_926 = 6'h1e == select_14 ? io_inData_30 : _GEN_925; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_927 = 6'h1f == select_14 ? io_inData_31 : _GEN_926; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_928 = 6'h20 == select_14 ? io_inData_32 : _GEN_927; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_929 = 6'h21 == select_14 ? io_inData_33 : _GEN_928; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_930 = 6'h22 == select_14 ? io_inData_34 : _GEN_929; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_931 = 6'h23 == select_14 ? io_inData_35 : _GEN_930; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_932 = 6'h24 == select_14 ? io_inData_36 : _GEN_931; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_933 = 6'h25 == select_14 ? io_inData_37 : _GEN_932; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_934 = 6'h26 == select_14 ? io_inData_38 : _GEN_933; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_935 = 6'h27 == select_14 ? io_inData_39 : _GEN_934; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_936 = 6'h28 == select_14 ? io_inData_40 : _GEN_935; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_937 = 6'h29 == select_14 ? io_inData_41 : _GEN_936; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_938 = 6'h2a == select_14 ? io_inData_42 : _GEN_937; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_939 = 6'h2b == select_14 ? io_inData_43 : _GEN_938; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_940 = 6'h2c == select_14 ? io_inData_44 : _GEN_939; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_941 = 6'h2d == select_14 ? io_inData_45 : _GEN_940; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_942 = 6'h2e == select_14 ? io_inData_46 : _GEN_941; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_943 = 6'h2f == select_14 ? io_inData_47 : _GEN_942; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_944 = 6'h30 == select_14 ? io_inData_48 : _GEN_943; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_945 = 6'h31 == select_14 ? io_inData_49 : _GEN_944; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_946 = 6'h32 == select_14 ? io_inData_50 : _GEN_945; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_947 = 6'h33 == select_14 ? io_inData_51 : _GEN_946; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_948 = 6'h34 == select_14 ? io_inData_52 : _GEN_947; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_949 = 6'h35 == select_14 ? io_inData_53 : _GEN_948; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_950 = 6'h36 == select_14 ? io_inData_54 : _GEN_949; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_951 = 6'h37 == select_14 ? io_inData_55 : _GEN_950; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_952 = 6'h38 == select_14 ? io_inData_56 : _GEN_951; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_953 = 6'h39 == select_14 ? io_inData_57 : _GEN_952; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_954 = 6'h3a == select_14 ? io_inData_58 : _GEN_953; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_955 = 6'h3b == select_14 ? io_inData_59 : _GEN_954; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_956 = 6'h3c == select_14 ? io_inData_60 : _GEN_955; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_957 = 6'h3d == select_14 ? io_inData_61 : _GEN_956; // @[Switch.scala 33:19:@4774.4]
  assign _GEN_958 = 6'h3e == select_14 ? io_inData_62 : _GEN_957; // @[Switch.scala 33:19:@4774.4]
  assign _T_23369 = {valid_14_7,valid_14_6,valid_14_5,valid_14_4,valid_14_3,valid_14_2,valid_14_1,valid_14_0}; // @[Switch.scala 34:32:@4781.4]
  assign _T_23377 = {valid_14_15,valid_14_14,valid_14_13,valid_14_12,valid_14_11,valid_14_10,valid_14_9,valid_14_8,_T_23369}; // @[Switch.scala 34:32:@4789.4]
  assign _T_23384 = {valid_14_23,valid_14_22,valid_14_21,valid_14_20,valid_14_19,valid_14_18,valid_14_17,valid_14_16}; // @[Switch.scala 34:32:@4796.4]
  assign _T_23393 = {valid_14_31,valid_14_30,valid_14_29,valid_14_28,valid_14_27,valid_14_26,valid_14_25,valid_14_24,_T_23384,_T_23377}; // @[Switch.scala 34:32:@4805.4]
  assign _T_23400 = {valid_14_39,valid_14_38,valid_14_37,valid_14_36,valid_14_35,valid_14_34,valid_14_33,valid_14_32}; // @[Switch.scala 34:32:@4812.4]
  assign _T_23408 = {valid_14_47,valid_14_46,valid_14_45,valid_14_44,valid_14_43,valid_14_42,valid_14_41,valid_14_40,_T_23400}; // @[Switch.scala 34:32:@4820.4]
  assign _T_23415 = {valid_14_55,valid_14_54,valid_14_53,valid_14_52,valid_14_51,valid_14_50,valid_14_49,valid_14_48}; // @[Switch.scala 34:32:@4827.4]
  assign _T_23424 = {valid_14_63,valid_14_62,valid_14_61,valid_14_60,valid_14_59,valid_14_58,valid_14_57,valid_14_56,_T_23415,_T_23408}; // @[Switch.scala 34:32:@4836.4]
  assign _T_23425 = {_T_23424,_T_23393}; // @[Switch.scala 34:32:@4837.4]
  assign _T_23429 = io_inAddr_0 == 6'hf; // @[Switch.scala 30:53:@4840.4]
  assign valid_15_0 = io_inValid_0 & _T_23429; // @[Switch.scala 30:36:@4841.4]
  assign _T_23432 = io_inAddr_1 == 6'hf; // @[Switch.scala 30:53:@4843.4]
  assign valid_15_1 = io_inValid_1 & _T_23432; // @[Switch.scala 30:36:@4844.4]
  assign _T_23435 = io_inAddr_2 == 6'hf; // @[Switch.scala 30:53:@4846.4]
  assign valid_15_2 = io_inValid_2 & _T_23435; // @[Switch.scala 30:36:@4847.4]
  assign _T_23438 = io_inAddr_3 == 6'hf; // @[Switch.scala 30:53:@4849.4]
  assign valid_15_3 = io_inValid_3 & _T_23438; // @[Switch.scala 30:36:@4850.4]
  assign _T_23441 = io_inAddr_4 == 6'hf; // @[Switch.scala 30:53:@4852.4]
  assign valid_15_4 = io_inValid_4 & _T_23441; // @[Switch.scala 30:36:@4853.4]
  assign _T_23444 = io_inAddr_5 == 6'hf; // @[Switch.scala 30:53:@4855.4]
  assign valid_15_5 = io_inValid_5 & _T_23444; // @[Switch.scala 30:36:@4856.4]
  assign _T_23447 = io_inAddr_6 == 6'hf; // @[Switch.scala 30:53:@4858.4]
  assign valid_15_6 = io_inValid_6 & _T_23447; // @[Switch.scala 30:36:@4859.4]
  assign _T_23450 = io_inAddr_7 == 6'hf; // @[Switch.scala 30:53:@4861.4]
  assign valid_15_7 = io_inValid_7 & _T_23450; // @[Switch.scala 30:36:@4862.4]
  assign _T_23453 = io_inAddr_8 == 6'hf; // @[Switch.scala 30:53:@4864.4]
  assign valid_15_8 = io_inValid_8 & _T_23453; // @[Switch.scala 30:36:@4865.4]
  assign _T_23456 = io_inAddr_9 == 6'hf; // @[Switch.scala 30:53:@4867.4]
  assign valid_15_9 = io_inValid_9 & _T_23456; // @[Switch.scala 30:36:@4868.4]
  assign _T_23459 = io_inAddr_10 == 6'hf; // @[Switch.scala 30:53:@4870.4]
  assign valid_15_10 = io_inValid_10 & _T_23459; // @[Switch.scala 30:36:@4871.4]
  assign _T_23462 = io_inAddr_11 == 6'hf; // @[Switch.scala 30:53:@4873.4]
  assign valid_15_11 = io_inValid_11 & _T_23462; // @[Switch.scala 30:36:@4874.4]
  assign _T_23465 = io_inAddr_12 == 6'hf; // @[Switch.scala 30:53:@4876.4]
  assign valid_15_12 = io_inValid_12 & _T_23465; // @[Switch.scala 30:36:@4877.4]
  assign _T_23468 = io_inAddr_13 == 6'hf; // @[Switch.scala 30:53:@4879.4]
  assign valid_15_13 = io_inValid_13 & _T_23468; // @[Switch.scala 30:36:@4880.4]
  assign _T_23471 = io_inAddr_14 == 6'hf; // @[Switch.scala 30:53:@4882.4]
  assign valid_15_14 = io_inValid_14 & _T_23471; // @[Switch.scala 30:36:@4883.4]
  assign _T_23474 = io_inAddr_15 == 6'hf; // @[Switch.scala 30:53:@4885.4]
  assign valid_15_15 = io_inValid_15 & _T_23474; // @[Switch.scala 30:36:@4886.4]
  assign _T_23477 = io_inAddr_16 == 6'hf; // @[Switch.scala 30:53:@4888.4]
  assign valid_15_16 = io_inValid_16 & _T_23477; // @[Switch.scala 30:36:@4889.4]
  assign _T_23480 = io_inAddr_17 == 6'hf; // @[Switch.scala 30:53:@4891.4]
  assign valid_15_17 = io_inValid_17 & _T_23480; // @[Switch.scala 30:36:@4892.4]
  assign _T_23483 = io_inAddr_18 == 6'hf; // @[Switch.scala 30:53:@4894.4]
  assign valid_15_18 = io_inValid_18 & _T_23483; // @[Switch.scala 30:36:@4895.4]
  assign _T_23486 = io_inAddr_19 == 6'hf; // @[Switch.scala 30:53:@4897.4]
  assign valid_15_19 = io_inValid_19 & _T_23486; // @[Switch.scala 30:36:@4898.4]
  assign _T_23489 = io_inAddr_20 == 6'hf; // @[Switch.scala 30:53:@4900.4]
  assign valid_15_20 = io_inValid_20 & _T_23489; // @[Switch.scala 30:36:@4901.4]
  assign _T_23492 = io_inAddr_21 == 6'hf; // @[Switch.scala 30:53:@4903.4]
  assign valid_15_21 = io_inValid_21 & _T_23492; // @[Switch.scala 30:36:@4904.4]
  assign _T_23495 = io_inAddr_22 == 6'hf; // @[Switch.scala 30:53:@4906.4]
  assign valid_15_22 = io_inValid_22 & _T_23495; // @[Switch.scala 30:36:@4907.4]
  assign _T_23498 = io_inAddr_23 == 6'hf; // @[Switch.scala 30:53:@4909.4]
  assign valid_15_23 = io_inValid_23 & _T_23498; // @[Switch.scala 30:36:@4910.4]
  assign _T_23501 = io_inAddr_24 == 6'hf; // @[Switch.scala 30:53:@4912.4]
  assign valid_15_24 = io_inValid_24 & _T_23501; // @[Switch.scala 30:36:@4913.4]
  assign _T_23504 = io_inAddr_25 == 6'hf; // @[Switch.scala 30:53:@4915.4]
  assign valid_15_25 = io_inValid_25 & _T_23504; // @[Switch.scala 30:36:@4916.4]
  assign _T_23507 = io_inAddr_26 == 6'hf; // @[Switch.scala 30:53:@4918.4]
  assign valid_15_26 = io_inValid_26 & _T_23507; // @[Switch.scala 30:36:@4919.4]
  assign _T_23510 = io_inAddr_27 == 6'hf; // @[Switch.scala 30:53:@4921.4]
  assign valid_15_27 = io_inValid_27 & _T_23510; // @[Switch.scala 30:36:@4922.4]
  assign _T_23513 = io_inAddr_28 == 6'hf; // @[Switch.scala 30:53:@4924.4]
  assign valid_15_28 = io_inValid_28 & _T_23513; // @[Switch.scala 30:36:@4925.4]
  assign _T_23516 = io_inAddr_29 == 6'hf; // @[Switch.scala 30:53:@4927.4]
  assign valid_15_29 = io_inValid_29 & _T_23516; // @[Switch.scala 30:36:@4928.4]
  assign _T_23519 = io_inAddr_30 == 6'hf; // @[Switch.scala 30:53:@4930.4]
  assign valid_15_30 = io_inValid_30 & _T_23519; // @[Switch.scala 30:36:@4931.4]
  assign _T_23522 = io_inAddr_31 == 6'hf; // @[Switch.scala 30:53:@4933.4]
  assign valid_15_31 = io_inValid_31 & _T_23522; // @[Switch.scala 30:36:@4934.4]
  assign _T_23525 = io_inAddr_32 == 6'hf; // @[Switch.scala 30:53:@4936.4]
  assign valid_15_32 = io_inValid_32 & _T_23525; // @[Switch.scala 30:36:@4937.4]
  assign _T_23528 = io_inAddr_33 == 6'hf; // @[Switch.scala 30:53:@4939.4]
  assign valid_15_33 = io_inValid_33 & _T_23528; // @[Switch.scala 30:36:@4940.4]
  assign _T_23531 = io_inAddr_34 == 6'hf; // @[Switch.scala 30:53:@4942.4]
  assign valid_15_34 = io_inValid_34 & _T_23531; // @[Switch.scala 30:36:@4943.4]
  assign _T_23534 = io_inAddr_35 == 6'hf; // @[Switch.scala 30:53:@4945.4]
  assign valid_15_35 = io_inValid_35 & _T_23534; // @[Switch.scala 30:36:@4946.4]
  assign _T_23537 = io_inAddr_36 == 6'hf; // @[Switch.scala 30:53:@4948.4]
  assign valid_15_36 = io_inValid_36 & _T_23537; // @[Switch.scala 30:36:@4949.4]
  assign _T_23540 = io_inAddr_37 == 6'hf; // @[Switch.scala 30:53:@4951.4]
  assign valid_15_37 = io_inValid_37 & _T_23540; // @[Switch.scala 30:36:@4952.4]
  assign _T_23543 = io_inAddr_38 == 6'hf; // @[Switch.scala 30:53:@4954.4]
  assign valid_15_38 = io_inValid_38 & _T_23543; // @[Switch.scala 30:36:@4955.4]
  assign _T_23546 = io_inAddr_39 == 6'hf; // @[Switch.scala 30:53:@4957.4]
  assign valid_15_39 = io_inValid_39 & _T_23546; // @[Switch.scala 30:36:@4958.4]
  assign _T_23549 = io_inAddr_40 == 6'hf; // @[Switch.scala 30:53:@4960.4]
  assign valid_15_40 = io_inValid_40 & _T_23549; // @[Switch.scala 30:36:@4961.4]
  assign _T_23552 = io_inAddr_41 == 6'hf; // @[Switch.scala 30:53:@4963.4]
  assign valid_15_41 = io_inValid_41 & _T_23552; // @[Switch.scala 30:36:@4964.4]
  assign _T_23555 = io_inAddr_42 == 6'hf; // @[Switch.scala 30:53:@4966.4]
  assign valid_15_42 = io_inValid_42 & _T_23555; // @[Switch.scala 30:36:@4967.4]
  assign _T_23558 = io_inAddr_43 == 6'hf; // @[Switch.scala 30:53:@4969.4]
  assign valid_15_43 = io_inValid_43 & _T_23558; // @[Switch.scala 30:36:@4970.4]
  assign _T_23561 = io_inAddr_44 == 6'hf; // @[Switch.scala 30:53:@4972.4]
  assign valid_15_44 = io_inValid_44 & _T_23561; // @[Switch.scala 30:36:@4973.4]
  assign _T_23564 = io_inAddr_45 == 6'hf; // @[Switch.scala 30:53:@4975.4]
  assign valid_15_45 = io_inValid_45 & _T_23564; // @[Switch.scala 30:36:@4976.4]
  assign _T_23567 = io_inAddr_46 == 6'hf; // @[Switch.scala 30:53:@4978.4]
  assign valid_15_46 = io_inValid_46 & _T_23567; // @[Switch.scala 30:36:@4979.4]
  assign _T_23570 = io_inAddr_47 == 6'hf; // @[Switch.scala 30:53:@4981.4]
  assign valid_15_47 = io_inValid_47 & _T_23570; // @[Switch.scala 30:36:@4982.4]
  assign _T_23573 = io_inAddr_48 == 6'hf; // @[Switch.scala 30:53:@4984.4]
  assign valid_15_48 = io_inValid_48 & _T_23573; // @[Switch.scala 30:36:@4985.4]
  assign _T_23576 = io_inAddr_49 == 6'hf; // @[Switch.scala 30:53:@4987.4]
  assign valid_15_49 = io_inValid_49 & _T_23576; // @[Switch.scala 30:36:@4988.4]
  assign _T_23579 = io_inAddr_50 == 6'hf; // @[Switch.scala 30:53:@4990.4]
  assign valid_15_50 = io_inValid_50 & _T_23579; // @[Switch.scala 30:36:@4991.4]
  assign _T_23582 = io_inAddr_51 == 6'hf; // @[Switch.scala 30:53:@4993.4]
  assign valid_15_51 = io_inValid_51 & _T_23582; // @[Switch.scala 30:36:@4994.4]
  assign _T_23585 = io_inAddr_52 == 6'hf; // @[Switch.scala 30:53:@4996.4]
  assign valid_15_52 = io_inValid_52 & _T_23585; // @[Switch.scala 30:36:@4997.4]
  assign _T_23588 = io_inAddr_53 == 6'hf; // @[Switch.scala 30:53:@4999.4]
  assign valid_15_53 = io_inValid_53 & _T_23588; // @[Switch.scala 30:36:@5000.4]
  assign _T_23591 = io_inAddr_54 == 6'hf; // @[Switch.scala 30:53:@5002.4]
  assign valid_15_54 = io_inValid_54 & _T_23591; // @[Switch.scala 30:36:@5003.4]
  assign _T_23594 = io_inAddr_55 == 6'hf; // @[Switch.scala 30:53:@5005.4]
  assign valid_15_55 = io_inValid_55 & _T_23594; // @[Switch.scala 30:36:@5006.4]
  assign _T_23597 = io_inAddr_56 == 6'hf; // @[Switch.scala 30:53:@5008.4]
  assign valid_15_56 = io_inValid_56 & _T_23597; // @[Switch.scala 30:36:@5009.4]
  assign _T_23600 = io_inAddr_57 == 6'hf; // @[Switch.scala 30:53:@5011.4]
  assign valid_15_57 = io_inValid_57 & _T_23600; // @[Switch.scala 30:36:@5012.4]
  assign _T_23603 = io_inAddr_58 == 6'hf; // @[Switch.scala 30:53:@5014.4]
  assign valid_15_58 = io_inValid_58 & _T_23603; // @[Switch.scala 30:36:@5015.4]
  assign _T_23606 = io_inAddr_59 == 6'hf; // @[Switch.scala 30:53:@5017.4]
  assign valid_15_59 = io_inValid_59 & _T_23606; // @[Switch.scala 30:36:@5018.4]
  assign _T_23609 = io_inAddr_60 == 6'hf; // @[Switch.scala 30:53:@5020.4]
  assign valid_15_60 = io_inValid_60 & _T_23609; // @[Switch.scala 30:36:@5021.4]
  assign _T_23612 = io_inAddr_61 == 6'hf; // @[Switch.scala 30:53:@5023.4]
  assign valid_15_61 = io_inValid_61 & _T_23612; // @[Switch.scala 30:36:@5024.4]
  assign _T_23615 = io_inAddr_62 == 6'hf; // @[Switch.scala 30:53:@5026.4]
  assign valid_15_62 = io_inValid_62 & _T_23615; // @[Switch.scala 30:36:@5027.4]
  assign _T_23618 = io_inAddr_63 == 6'hf; // @[Switch.scala 30:53:@5029.4]
  assign valid_15_63 = io_inValid_63 & _T_23618; // @[Switch.scala 30:36:@5030.4]
  assign _T_23684 = valid_15_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@5032.4]
  assign _T_23685 = valid_15_61 ? 6'h3d : _T_23684; // @[Mux.scala 31:69:@5033.4]
  assign _T_23686 = valid_15_60 ? 6'h3c : _T_23685; // @[Mux.scala 31:69:@5034.4]
  assign _T_23687 = valid_15_59 ? 6'h3b : _T_23686; // @[Mux.scala 31:69:@5035.4]
  assign _T_23688 = valid_15_58 ? 6'h3a : _T_23687; // @[Mux.scala 31:69:@5036.4]
  assign _T_23689 = valid_15_57 ? 6'h39 : _T_23688; // @[Mux.scala 31:69:@5037.4]
  assign _T_23690 = valid_15_56 ? 6'h38 : _T_23689; // @[Mux.scala 31:69:@5038.4]
  assign _T_23691 = valid_15_55 ? 6'h37 : _T_23690; // @[Mux.scala 31:69:@5039.4]
  assign _T_23692 = valid_15_54 ? 6'h36 : _T_23691; // @[Mux.scala 31:69:@5040.4]
  assign _T_23693 = valid_15_53 ? 6'h35 : _T_23692; // @[Mux.scala 31:69:@5041.4]
  assign _T_23694 = valid_15_52 ? 6'h34 : _T_23693; // @[Mux.scala 31:69:@5042.4]
  assign _T_23695 = valid_15_51 ? 6'h33 : _T_23694; // @[Mux.scala 31:69:@5043.4]
  assign _T_23696 = valid_15_50 ? 6'h32 : _T_23695; // @[Mux.scala 31:69:@5044.4]
  assign _T_23697 = valid_15_49 ? 6'h31 : _T_23696; // @[Mux.scala 31:69:@5045.4]
  assign _T_23698 = valid_15_48 ? 6'h30 : _T_23697; // @[Mux.scala 31:69:@5046.4]
  assign _T_23699 = valid_15_47 ? 6'h2f : _T_23698; // @[Mux.scala 31:69:@5047.4]
  assign _T_23700 = valid_15_46 ? 6'h2e : _T_23699; // @[Mux.scala 31:69:@5048.4]
  assign _T_23701 = valid_15_45 ? 6'h2d : _T_23700; // @[Mux.scala 31:69:@5049.4]
  assign _T_23702 = valid_15_44 ? 6'h2c : _T_23701; // @[Mux.scala 31:69:@5050.4]
  assign _T_23703 = valid_15_43 ? 6'h2b : _T_23702; // @[Mux.scala 31:69:@5051.4]
  assign _T_23704 = valid_15_42 ? 6'h2a : _T_23703; // @[Mux.scala 31:69:@5052.4]
  assign _T_23705 = valid_15_41 ? 6'h29 : _T_23704; // @[Mux.scala 31:69:@5053.4]
  assign _T_23706 = valid_15_40 ? 6'h28 : _T_23705; // @[Mux.scala 31:69:@5054.4]
  assign _T_23707 = valid_15_39 ? 6'h27 : _T_23706; // @[Mux.scala 31:69:@5055.4]
  assign _T_23708 = valid_15_38 ? 6'h26 : _T_23707; // @[Mux.scala 31:69:@5056.4]
  assign _T_23709 = valid_15_37 ? 6'h25 : _T_23708; // @[Mux.scala 31:69:@5057.4]
  assign _T_23710 = valid_15_36 ? 6'h24 : _T_23709; // @[Mux.scala 31:69:@5058.4]
  assign _T_23711 = valid_15_35 ? 6'h23 : _T_23710; // @[Mux.scala 31:69:@5059.4]
  assign _T_23712 = valid_15_34 ? 6'h22 : _T_23711; // @[Mux.scala 31:69:@5060.4]
  assign _T_23713 = valid_15_33 ? 6'h21 : _T_23712; // @[Mux.scala 31:69:@5061.4]
  assign _T_23714 = valid_15_32 ? 6'h20 : _T_23713; // @[Mux.scala 31:69:@5062.4]
  assign _T_23715 = valid_15_31 ? 6'h1f : _T_23714; // @[Mux.scala 31:69:@5063.4]
  assign _T_23716 = valid_15_30 ? 6'h1e : _T_23715; // @[Mux.scala 31:69:@5064.4]
  assign _T_23717 = valid_15_29 ? 6'h1d : _T_23716; // @[Mux.scala 31:69:@5065.4]
  assign _T_23718 = valid_15_28 ? 6'h1c : _T_23717; // @[Mux.scala 31:69:@5066.4]
  assign _T_23719 = valid_15_27 ? 6'h1b : _T_23718; // @[Mux.scala 31:69:@5067.4]
  assign _T_23720 = valid_15_26 ? 6'h1a : _T_23719; // @[Mux.scala 31:69:@5068.4]
  assign _T_23721 = valid_15_25 ? 6'h19 : _T_23720; // @[Mux.scala 31:69:@5069.4]
  assign _T_23722 = valid_15_24 ? 6'h18 : _T_23721; // @[Mux.scala 31:69:@5070.4]
  assign _T_23723 = valid_15_23 ? 6'h17 : _T_23722; // @[Mux.scala 31:69:@5071.4]
  assign _T_23724 = valid_15_22 ? 6'h16 : _T_23723; // @[Mux.scala 31:69:@5072.4]
  assign _T_23725 = valid_15_21 ? 6'h15 : _T_23724; // @[Mux.scala 31:69:@5073.4]
  assign _T_23726 = valid_15_20 ? 6'h14 : _T_23725; // @[Mux.scala 31:69:@5074.4]
  assign _T_23727 = valid_15_19 ? 6'h13 : _T_23726; // @[Mux.scala 31:69:@5075.4]
  assign _T_23728 = valid_15_18 ? 6'h12 : _T_23727; // @[Mux.scala 31:69:@5076.4]
  assign _T_23729 = valid_15_17 ? 6'h11 : _T_23728; // @[Mux.scala 31:69:@5077.4]
  assign _T_23730 = valid_15_16 ? 6'h10 : _T_23729; // @[Mux.scala 31:69:@5078.4]
  assign _T_23731 = valid_15_15 ? 6'hf : _T_23730; // @[Mux.scala 31:69:@5079.4]
  assign _T_23732 = valid_15_14 ? 6'he : _T_23731; // @[Mux.scala 31:69:@5080.4]
  assign _T_23733 = valid_15_13 ? 6'hd : _T_23732; // @[Mux.scala 31:69:@5081.4]
  assign _T_23734 = valid_15_12 ? 6'hc : _T_23733; // @[Mux.scala 31:69:@5082.4]
  assign _T_23735 = valid_15_11 ? 6'hb : _T_23734; // @[Mux.scala 31:69:@5083.4]
  assign _T_23736 = valid_15_10 ? 6'ha : _T_23735; // @[Mux.scala 31:69:@5084.4]
  assign _T_23737 = valid_15_9 ? 6'h9 : _T_23736; // @[Mux.scala 31:69:@5085.4]
  assign _T_23738 = valid_15_8 ? 6'h8 : _T_23737; // @[Mux.scala 31:69:@5086.4]
  assign _T_23739 = valid_15_7 ? 6'h7 : _T_23738; // @[Mux.scala 31:69:@5087.4]
  assign _T_23740 = valid_15_6 ? 6'h6 : _T_23739; // @[Mux.scala 31:69:@5088.4]
  assign _T_23741 = valid_15_5 ? 6'h5 : _T_23740; // @[Mux.scala 31:69:@5089.4]
  assign _T_23742 = valid_15_4 ? 6'h4 : _T_23741; // @[Mux.scala 31:69:@5090.4]
  assign _T_23743 = valid_15_3 ? 6'h3 : _T_23742; // @[Mux.scala 31:69:@5091.4]
  assign _T_23744 = valid_15_2 ? 6'h2 : _T_23743; // @[Mux.scala 31:69:@5092.4]
  assign _T_23745 = valid_15_1 ? 6'h1 : _T_23744; // @[Mux.scala 31:69:@5093.4]
  assign select_15 = valid_15_0 ? 6'h0 : _T_23745; // @[Mux.scala 31:69:@5094.4]
  assign _GEN_961 = 6'h1 == select_15 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_962 = 6'h2 == select_15 ? io_inData_2 : _GEN_961; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_963 = 6'h3 == select_15 ? io_inData_3 : _GEN_962; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_964 = 6'h4 == select_15 ? io_inData_4 : _GEN_963; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_965 = 6'h5 == select_15 ? io_inData_5 : _GEN_964; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_966 = 6'h6 == select_15 ? io_inData_6 : _GEN_965; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_967 = 6'h7 == select_15 ? io_inData_7 : _GEN_966; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_968 = 6'h8 == select_15 ? io_inData_8 : _GEN_967; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_969 = 6'h9 == select_15 ? io_inData_9 : _GEN_968; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_970 = 6'ha == select_15 ? io_inData_10 : _GEN_969; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_971 = 6'hb == select_15 ? io_inData_11 : _GEN_970; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_972 = 6'hc == select_15 ? io_inData_12 : _GEN_971; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_973 = 6'hd == select_15 ? io_inData_13 : _GEN_972; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_974 = 6'he == select_15 ? io_inData_14 : _GEN_973; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_975 = 6'hf == select_15 ? io_inData_15 : _GEN_974; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_976 = 6'h10 == select_15 ? io_inData_16 : _GEN_975; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_977 = 6'h11 == select_15 ? io_inData_17 : _GEN_976; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_978 = 6'h12 == select_15 ? io_inData_18 : _GEN_977; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_979 = 6'h13 == select_15 ? io_inData_19 : _GEN_978; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_980 = 6'h14 == select_15 ? io_inData_20 : _GEN_979; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_981 = 6'h15 == select_15 ? io_inData_21 : _GEN_980; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_982 = 6'h16 == select_15 ? io_inData_22 : _GEN_981; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_983 = 6'h17 == select_15 ? io_inData_23 : _GEN_982; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_984 = 6'h18 == select_15 ? io_inData_24 : _GEN_983; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_985 = 6'h19 == select_15 ? io_inData_25 : _GEN_984; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_986 = 6'h1a == select_15 ? io_inData_26 : _GEN_985; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_987 = 6'h1b == select_15 ? io_inData_27 : _GEN_986; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_988 = 6'h1c == select_15 ? io_inData_28 : _GEN_987; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_989 = 6'h1d == select_15 ? io_inData_29 : _GEN_988; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_990 = 6'h1e == select_15 ? io_inData_30 : _GEN_989; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_991 = 6'h1f == select_15 ? io_inData_31 : _GEN_990; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_992 = 6'h20 == select_15 ? io_inData_32 : _GEN_991; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_993 = 6'h21 == select_15 ? io_inData_33 : _GEN_992; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_994 = 6'h22 == select_15 ? io_inData_34 : _GEN_993; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_995 = 6'h23 == select_15 ? io_inData_35 : _GEN_994; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_996 = 6'h24 == select_15 ? io_inData_36 : _GEN_995; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_997 = 6'h25 == select_15 ? io_inData_37 : _GEN_996; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_998 = 6'h26 == select_15 ? io_inData_38 : _GEN_997; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_999 = 6'h27 == select_15 ? io_inData_39 : _GEN_998; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_1000 = 6'h28 == select_15 ? io_inData_40 : _GEN_999; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_1001 = 6'h29 == select_15 ? io_inData_41 : _GEN_1000; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_1002 = 6'h2a == select_15 ? io_inData_42 : _GEN_1001; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_1003 = 6'h2b == select_15 ? io_inData_43 : _GEN_1002; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_1004 = 6'h2c == select_15 ? io_inData_44 : _GEN_1003; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_1005 = 6'h2d == select_15 ? io_inData_45 : _GEN_1004; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_1006 = 6'h2e == select_15 ? io_inData_46 : _GEN_1005; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_1007 = 6'h2f == select_15 ? io_inData_47 : _GEN_1006; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_1008 = 6'h30 == select_15 ? io_inData_48 : _GEN_1007; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_1009 = 6'h31 == select_15 ? io_inData_49 : _GEN_1008; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_1010 = 6'h32 == select_15 ? io_inData_50 : _GEN_1009; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_1011 = 6'h33 == select_15 ? io_inData_51 : _GEN_1010; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_1012 = 6'h34 == select_15 ? io_inData_52 : _GEN_1011; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_1013 = 6'h35 == select_15 ? io_inData_53 : _GEN_1012; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_1014 = 6'h36 == select_15 ? io_inData_54 : _GEN_1013; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_1015 = 6'h37 == select_15 ? io_inData_55 : _GEN_1014; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_1016 = 6'h38 == select_15 ? io_inData_56 : _GEN_1015; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_1017 = 6'h39 == select_15 ? io_inData_57 : _GEN_1016; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_1018 = 6'h3a == select_15 ? io_inData_58 : _GEN_1017; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_1019 = 6'h3b == select_15 ? io_inData_59 : _GEN_1018; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_1020 = 6'h3c == select_15 ? io_inData_60 : _GEN_1019; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_1021 = 6'h3d == select_15 ? io_inData_61 : _GEN_1020; // @[Switch.scala 33:19:@5096.4]
  assign _GEN_1022 = 6'h3e == select_15 ? io_inData_62 : _GEN_1021; // @[Switch.scala 33:19:@5096.4]
  assign _T_23754 = {valid_15_7,valid_15_6,valid_15_5,valid_15_4,valid_15_3,valid_15_2,valid_15_1,valid_15_0}; // @[Switch.scala 34:32:@5103.4]
  assign _T_23762 = {valid_15_15,valid_15_14,valid_15_13,valid_15_12,valid_15_11,valid_15_10,valid_15_9,valid_15_8,_T_23754}; // @[Switch.scala 34:32:@5111.4]
  assign _T_23769 = {valid_15_23,valid_15_22,valid_15_21,valid_15_20,valid_15_19,valid_15_18,valid_15_17,valid_15_16}; // @[Switch.scala 34:32:@5118.4]
  assign _T_23778 = {valid_15_31,valid_15_30,valid_15_29,valid_15_28,valid_15_27,valid_15_26,valid_15_25,valid_15_24,_T_23769,_T_23762}; // @[Switch.scala 34:32:@5127.4]
  assign _T_23785 = {valid_15_39,valid_15_38,valid_15_37,valid_15_36,valid_15_35,valid_15_34,valid_15_33,valid_15_32}; // @[Switch.scala 34:32:@5134.4]
  assign _T_23793 = {valid_15_47,valid_15_46,valid_15_45,valid_15_44,valid_15_43,valid_15_42,valid_15_41,valid_15_40,_T_23785}; // @[Switch.scala 34:32:@5142.4]
  assign _T_23800 = {valid_15_55,valid_15_54,valid_15_53,valid_15_52,valid_15_51,valid_15_50,valid_15_49,valid_15_48}; // @[Switch.scala 34:32:@5149.4]
  assign _T_23809 = {valid_15_63,valid_15_62,valid_15_61,valid_15_60,valid_15_59,valid_15_58,valid_15_57,valid_15_56,_T_23800,_T_23793}; // @[Switch.scala 34:32:@5158.4]
  assign _T_23810 = {_T_23809,_T_23778}; // @[Switch.scala 34:32:@5159.4]
  assign _T_23814 = io_inAddr_0 == 6'h10; // @[Switch.scala 30:53:@5162.4]
  assign valid_16_0 = io_inValid_0 & _T_23814; // @[Switch.scala 30:36:@5163.4]
  assign _T_23817 = io_inAddr_1 == 6'h10; // @[Switch.scala 30:53:@5165.4]
  assign valid_16_1 = io_inValid_1 & _T_23817; // @[Switch.scala 30:36:@5166.4]
  assign _T_23820 = io_inAddr_2 == 6'h10; // @[Switch.scala 30:53:@5168.4]
  assign valid_16_2 = io_inValid_2 & _T_23820; // @[Switch.scala 30:36:@5169.4]
  assign _T_23823 = io_inAddr_3 == 6'h10; // @[Switch.scala 30:53:@5171.4]
  assign valid_16_3 = io_inValid_3 & _T_23823; // @[Switch.scala 30:36:@5172.4]
  assign _T_23826 = io_inAddr_4 == 6'h10; // @[Switch.scala 30:53:@5174.4]
  assign valid_16_4 = io_inValid_4 & _T_23826; // @[Switch.scala 30:36:@5175.4]
  assign _T_23829 = io_inAddr_5 == 6'h10; // @[Switch.scala 30:53:@5177.4]
  assign valid_16_5 = io_inValid_5 & _T_23829; // @[Switch.scala 30:36:@5178.4]
  assign _T_23832 = io_inAddr_6 == 6'h10; // @[Switch.scala 30:53:@5180.4]
  assign valid_16_6 = io_inValid_6 & _T_23832; // @[Switch.scala 30:36:@5181.4]
  assign _T_23835 = io_inAddr_7 == 6'h10; // @[Switch.scala 30:53:@5183.4]
  assign valid_16_7 = io_inValid_7 & _T_23835; // @[Switch.scala 30:36:@5184.4]
  assign _T_23838 = io_inAddr_8 == 6'h10; // @[Switch.scala 30:53:@5186.4]
  assign valid_16_8 = io_inValid_8 & _T_23838; // @[Switch.scala 30:36:@5187.4]
  assign _T_23841 = io_inAddr_9 == 6'h10; // @[Switch.scala 30:53:@5189.4]
  assign valid_16_9 = io_inValid_9 & _T_23841; // @[Switch.scala 30:36:@5190.4]
  assign _T_23844 = io_inAddr_10 == 6'h10; // @[Switch.scala 30:53:@5192.4]
  assign valid_16_10 = io_inValid_10 & _T_23844; // @[Switch.scala 30:36:@5193.4]
  assign _T_23847 = io_inAddr_11 == 6'h10; // @[Switch.scala 30:53:@5195.4]
  assign valid_16_11 = io_inValid_11 & _T_23847; // @[Switch.scala 30:36:@5196.4]
  assign _T_23850 = io_inAddr_12 == 6'h10; // @[Switch.scala 30:53:@5198.4]
  assign valid_16_12 = io_inValid_12 & _T_23850; // @[Switch.scala 30:36:@5199.4]
  assign _T_23853 = io_inAddr_13 == 6'h10; // @[Switch.scala 30:53:@5201.4]
  assign valid_16_13 = io_inValid_13 & _T_23853; // @[Switch.scala 30:36:@5202.4]
  assign _T_23856 = io_inAddr_14 == 6'h10; // @[Switch.scala 30:53:@5204.4]
  assign valid_16_14 = io_inValid_14 & _T_23856; // @[Switch.scala 30:36:@5205.4]
  assign _T_23859 = io_inAddr_15 == 6'h10; // @[Switch.scala 30:53:@5207.4]
  assign valid_16_15 = io_inValid_15 & _T_23859; // @[Switch.scala 30:36:@5208.4]
  assign _T_23862 = io_inAddr_16 == 6'h10; // @[Switch.scala 30:53:@5210.4]
  assign valid_16_16 = io_inValid_16 & _T_23862; // @[Switch.scala 30:36:@5211.4]
  assign _T_23865 = io_inAddr_17 == 6'h10; // @[Switch.scala 30:53:@5213.4]
  assign valid_16_17 = io_inValid_17 & _T_23865; // @[Switch.scala 30:36:@5214.4]
  assign _T_23868 = io_inAddr_18 == 6'h10; // @[Switch.scala 30:53:@5216.4]
  assign valid_16_18 = io_inValid_18 & _T_23868; // @[Switch.scala 30:36:@5217.4]
  assign _T_23871 = io_inAddr_19 == 6'h10; // @[Switch.scala 30:53:@5219.4]
  assign valid_16_19 = io_inValid_19 & _T_23871; // @[Switch.scala 30:36:@5220.4]
  assign _T_23874 = io_inAddr_20 == 6'h10; // @[Switch.scala 30:53:@5222.4]
  assign valid_16_20 = io_inValid_20 & _T_23874; // @[Switch.scala 30:36:@5223.4]
  assign _T_23877 = io_inAddr_21 == 6'h10; // @[Switch.scala 30:53:@5225.4]
  assign valid_16_21 = io_inValid_21 & _T_23877; // @[Switch.scala 30:36:@5226.4]
  assign _T_23880 = io_inAddr_22 == 6'h10; // @[Switch.scala 30:53:@5228.4]
  assign valid_16_22 = io_inValid_22 & _T_23880; // @[Switch.scala 30:36:@5229.4]
  assign _T_23883 = io_inAddr_23 == 6'h10; // @[Switch.scala 30:53:@5231.4]
  assign valid_16_23 = io_inValid_23 & _T_23883; // @[Switch.scala 30:36:@5232.4]
  assign _T_23886 = io_inAddr_24 == 6'h10; // @[Switch.scala 30:53:@5234.4]
  assign valid_16_24 = io_inValid_24 & _T_23886; // @[Switch.scala 30:36:@5235.4]
  assign _T_23889 = io_inAddr_25 == 6'h10; // @[Switch.scala 30:53:@5237.4]
  assign valid_16_25 = io_inValid_25 & _T_23889; // @[Switch.scala 30:36:@5238.4]
  assign _T_23892 = io_inAddr_26 == 6'h10; // @[Switch.scala 30:53:@5240.4]
  assign valid_16_26 = io_inValid_26 & _T_23892; // @[Switch.scala 30:36:@5241.4]
  assign _T_23895 = io_inAddr_27 == 6'h10; // @[Switch.scala 30:53:@5243.4]
  assign valid_16_27 = io_inValid_27 & _T_23895; // @[Switch.scala 30:36:@5244.4]
  assign _T_23898 = io_inAddr_28 == 6'h10; // @[Switch.scala 30:53:@5246.4]
  assign valid_16_28 = io_inValid_28 & _T_23898; // @[Switch.scala 30:36:@5247.4]
  assign _T_23901 = io_inAddr_29 == 6'h10; // @[Switch.scala 30:53:@5249.4]
  assign valid_16_29 = io_inValid_29 & _T_23901; // @[Switch.scala 30:36:@5250.4]
  assign _T_23904 = io_inAddr_30 == 6'h10; // @[Switch.scala 30:53:@5252.4]
  assign valid_16_30 = io_inValid_30 & _T_23904; // @[Switch.scala 30:36:@5253.4]
  assign _T_23907 = io_inAddr_31 == 6'h10; // @[Switch.scala 30:53:@5255.4]
  assign valid_16_31 = io_inValid_31 & _T_23907; // @[Switch.scala 30:36:@5256.4]
  assign _T_23910 = io_inAddr_32 == 6'h10; // @[Switch.scala 30:53:@5258.4]
  assign valid_16_32 = io_inValid_32 & _T_23910; // @[Switch.scala 30:36:@5259.4]
  assign _T_23913 = io_inAddr_33 == 6'h10; // @[Switch.scala 30:53:@5261.4]
  assign valid_16_33 = io_inValid_33 & _T_23913; // @[Switch.scala 30:36:@5262.4]
  assign _T_23916 = io_inAddr_34 == 6'h10; // @[Switch.scala 30:53:@5264.4]
  assign valid_16_34 = io_inValid_34 & _T_23916; // @[Switch.scala 30:36:@5265.4]
  assign _T_23919 = io_inAddr_35 == 6'h10; // @[Switch.scala 30:53:@5267.4]
  assign valid_16_35 = io_inValid_35 & _T_23919; // @[Switch.scala 30:36:@5268.4]
  assign _T_23922 = io_inAddr_36 == 6'h10; // @[Switch.scala 30:53:@5270.4]
  assign valid_16_36 = io_inValid_36 & _T_23922; // @[Switch.scala 30:36:@5271.4]
  assign _T_23925 = io_inAddr_37 == 6'h10; // @[Switch.scala 30:53:@5273.4]
  assign valid_16_37 = io_inValid_37 & _T_23925; // @[Switch.scala 30:36:@5274.4]
  assign _T_23928 = io_inAddr_38 == 6'h10; // @[Switch.scala 30:53:@5276.4]
  assign valid_16_38 = io_inValid_38 & _T_23928; // @[Switch.scala 30:36:@5277.4]
  assign _T_23931 = io_inAddr_39 == 6'h10; // @[Switch.scala 30:53:@5279.4]
  assign valid_16_39 = io_inValid_39 & _T_23931; // @[Switch.scala 30:36:@5280.4]
  assign _T_23934 = io_inAddr_40 == 6'h10; // @[Switch.scala 30:53:@5282.4]
  assign valid_16_40 = io_inValid_40 & _T_23934; // @[Switch.scala 30:36:@5283.4]
  assign _T_23937 = io_inAddr_41 == 6'h10; // @[Switch.scala 30:53:@5285.4]
  assign valid_16_41 = io_inValid_41 & _T_23937; // @[Switch.scala 30:36:@5286.4]
  assign _T_23940 = io_inAddr_42 == 6'h10; // @[Switch.scala 30:53:@5288.4]
  assign valid_16_42 = io_inValid_42 & _T_23940; // @[Switch.scala 30:36:@5289.4]
  assign _T_23943 = io_inAddr_43 == 6'h10; // @[Switch.scala 30:53:@5291.4]
  assign valid_16_43 = io_inValid_43 & _T_23943; // @[Switch.scala 30:36:@5292.4]
  assign _T_23946 = io_inAddr_44 == 6'h10; // @[Switch.scala 30:53:@5294.4]
  assign valid_16_44 = io_inValid_44 & _T_23946; // @[Switch.scala 30:36:@5295.4]
  assign _T_23949 = io_inAddr_45 == 6'h10; // @[Switch.scala 30:53:@5297.4]
  assign valid_16_45 = io_inValid_45 & _T_23949; // @[Switch.scala 30:36:@5298.4]
  assign _T_23952 = io_inAddr_46 == 6'h10; // @[Switch.scala 30:53:@5300.4]
  assign valid_16_46 = io_inValid_46 & _T_23952; // @[Switch.scala 30:36:@5301.4]
  assign _T_23955 = io_inAddr_47 == 6'h10; // @[Switch.scala 30:53:@5303.4]
  assign valid_16_47 = io_inValid_47 & _T_23955; // @[Switch.scala 30:36:@5304.4]
  assign _T_23958 = io_inAddr_48 == 6'h10; // @[Switch.scala 30:53:@5306.4]
  assign valid_16_48 = io_inValid_48 & _T_23958; // @[Switch.scala 30:36:@5307.4]
  assign _T_23961 = io_inAddr_49 == 6'h10; // @[Switch.scala 30:53:@5309.4]
  assign valid_16_49 = io_inValid_49 & _T_23961; // @[Switch.scala 30:36:@5310.4]
  assign _T_23964 = io_inAddr_50 == 6'h10; // @[Switch.scala 30:53:@5312.4]
  assign valid_16_50 = io_inValid_50 & _T_23964; // @[Switch.scala 30:36:@5313.4]
  assign _T_23967 = io_inAddr_51 == 6'h10; // @[Switch.scala 30:53:@5315.4]
  assign valid_16_51 = io_inValid_51 & _T_23967; // @[Switch.scala 30:36:@5316.4]
  assign _T_23970 = io_inAddr_52 == 6'h10; // @[Switch.scala 30:53:@5318.4]
  assign valid_16_52 = io_inValid_52 & _T_23970; // @[Switch.scala 30:36:@5319.4]
  assign _T_23973 = io_inAddr_53 == 6'h10; // @[Switch.scala 30:53:@5321.4]
  assign valid_16_53 = io_inValid_53 & _T_23973; // @[Switch.scala 30:36:@5322.4]
  assign _T_23976 = io_inAddr_54 == 6'h10; // @[Switch.scala 30:53:@5324.4]
  assign valid_16_54 = io_inValid_54 & _T_23976; // @[Switch.scala 30:36:@5325.4]
  assign _T_23979 = io_inAddr_55 == 6'h10; // @[Switch.scala 30:53:@5327.4]
  assign valid_16_55 = io_inValid_55 & _T_23979; // @[Switch.scala 30:36:@5328.4]
  assign _T_23982 = io_inAddr_56 == 6'h10; // @[Switch.scala 30:53:@5330.4]
  assign valid_16_56 = io_inValid_56 & _T_23982; // @[Switch.scala 30:36:@5331.4]
  assign _T_23985 = io_inAddr_57 == 6'h10; // @[Switch.scala 30:53:@5333.4]
  assign valid_16_57 = io_inValid_57 & _T_23985; // @[Switch.scala 30:36:@5334.4]
  assign _T_23988 = io_inAddr_58 == 6'h10; // @[Switch.scala 30:53:@5336.4]
  assign valid_16_58 = io_inValid_58 & _T_23988; // @[Switch.scala 30:36:@5337.4]
  assign _T_23991 = io_inAddr_59 == 6'h10; // @[Switch.scala 30:53:@5339.4]
  assign valid_16_59 = io_inValid_59 & _T_23991; // @[Switch.scala 30:36:@5340.4]
  assign _T_23994 = io_inAddr_60 == 6'h10; // @[Switch.scala 30:53:@5342.4]
  assign valid_16_60 = io_inValid_60 & _T_23994; // @[Switch.scala 30:36:@5343.4]
  assign _T_23997 = io_inAddr_61 == 6'h10; // @[Switch.scala 30:53:@5345.4]
  assign valid_16_61 = io_inValid_61 & _T_23997; // @[Switch.scala 30:36:@5346.4]
  assign _T_24000 = io_inAddr_62 == 6'h10; // @[Switch.scala 30:53:@5348.4]
  assign valid_16_62 = io_inValid_62 & _T_24000; // @[Switch.scala 30:36:@5349.4]
  assign _T_24003 = io_inAddr_63 == 6'h10; // @[Switch.scala 30:53:@5351.4]
  assign valid_16_63 = io_inValid_63 & _T_24003; // @[Switch.scala 30:36:@5352.4]
  assign _T_24069 = valid_16_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@5354.4]
  assign _T_24070 = valid_16_61 ? 6'h3d : _T_24069; // @[Mux.scala 31:69:@5355.4]
  assign _T_24071 = valid_16_60 ? 6'h3c : _T_24070; // @[Mux.scala 31:69:@5356.4]
  assign _T_24072 = valid_16_59 ? 6'h3b : _T_24071; // @[Mux.scala 31:69:@5357.4]
  assign _T_24073 = valid_16_58 ? 6'h3a : _T_24072; // @[Mux.scala 31:69:@5358.4]
  assign _T_24074 = valid_16_57 ? 6'h39 : _T_24073; // @[Mux.scala 31:69:@5359.4]
  assign _T_24075 = valid_16_56 ? 6'h38 : _T_24074; // @[Mux.scala 31:69:@5360.4]
  assign _T_24076 = valid_16_55 ? 6'h37 : _T_24075; // @[Mux.scala 31:69:@5361.4]
  assign _T_24077 = valid_16_54 ? 6'h36 : _T_24076; // @[Mux.scala 31:69:@5362.4]
  assign _T_24078 = valid_16_53 ? 6'h35 : _T_24077; // @[Mux.scala 31:69:@5363.4]
  assign _T_24079 = valid_16_52 ? 6'h34 : _T_24078; // @[Mux.scala 31:69:@5364.4]
  assign _T_24080 = valid_16_51 ? 6'h33 : _T_24079; // @[Mux.scala 31:69:@5365.4]
  assign _T_24081 = valid_16_50 ? 6'h32 : _T_24080; // @[Mux.scala 31:69:@5366.4]
  assign _T_24082 = valid_16_49 ? 6'h31 : _T_24081; // @[Mux.scala 31:69:@5367.4]
  assign _T_24083 = valid_16_48 ? 6'h30 : _T_24082; // @[Mux.scala 31:69:@5368.4]
  assign _T_24084 = valid_16_47 ? 6'h2f : _T_24083; // @[Mux.scala 31:69:@5369.4]
  assign _T_24085 = valid_16_46 ? 6'h2e : _T_24084; // @[Mux.scala 31:69:@5370.4]
  assign _T_24086 = valid_16_45 ? 6'h2d : _T_24085; // @[Mux.scala 31:69:@5371.4]
  assign _T_24087 = valid_16_44 ? 6'h2c : _T_24086; // @[Mux.scala 31:69:@5372.4]
  assign _T_24088 = valid_16_43 ? 6'h2b : _T_24087; // @[Mux.scala 31:69:@5373.4]
  assign _T_24089 = valid_16_42 ? 6'h2a : _T_24088; // @[Mux.scala 31:69:@5374.4]
  assign _T_24090 = valid_16_41 ? 6'h29 : _T_24089; // @[Mux.scala 31:69:@5375.4]
  assign _T_24091 = valid_16_40 ? 6'h28 : _T_24090; // @[Mux.scala 31:69:@5376.4]
  assign _T_24092 = valid_16_39 ? 6'h27 : _T_24091; // @[Mux.scala 31:69:@5377.4]
  assign _T_24093 = valid_16_38 ? 6'h26 : _T_24092; // @[Mux.scala 31:69:@5378.4]
  assign _T_24094 = valid_16_37 ? 6'h25 : _T_24093; // @[Mux.scala 31:69:@5379.4]
  assign _T_24095 = valid_16_36 ? 6'h24 : _T_24094; // @[Mux.scala 31:69:@5380.4]
  assign _T_24096 = valid_16_35 ? 6'h23 : _T_24095; // @[Mux.scala 31:69:@5381.4]
  assign _T_24097 = valid_16_34 ? 6'h22 : _T_24096; // @[Mux.scala 31:69:@5382.4]
  assign _T_24098 = valid_16_33 ? 6'h21 : _T_24097; // @[Mux.scala 31:69:@5383.4]
  assign _T_24099 = valid_16_32 ? 6'h20 : _T_24098; // @[Mux.scala 31:69:@5384.4]
  assign _T_24100 = valid_16_31 ? 6'h1f : _T_24099; // @[Mux.scala 31:69:@5385.4]
  assign _T_24101 = valid_16_30 ? 6'h1e : _T_24100; // @[Mux.scala 31:69:@5386.4]
  assign _T_24102 = valid_16_29 ? 6'h1d : _T_24101; // @[Mux.scala 31:69:@5387.4]
  assign _T_24103 = valid_16_28 ? 6'h1c : _T_24102; // @[Mux.scala 31:69:@5388.4]
  assign _T_24104 = valid_16_27 ? 6'h1b : _T_24103; // @[Mux.scala 31:69:@5389.4]
  assign _T_24105 = valid_16_26 ? 6'h1a : _T_24104; // @[Mux.scala 31:69:@5390.4]
  assign _T_24106 = valid_16_25 ? 6'h19 : _T_24105; // @[Mux.scala 31:69:@5391.4]
  assign _T_24107 = valid_16_24 ? 6'h18 : _T_24106; // @[Mux.scala 31:69:@5392.4]
  assign _T_24108 = valid_16_23 ? 6'h17 : _T_24107; // @[Mux.scala 31:69:@5393.4]
  assign _T_24109 = valid_16_22 ? 6'h16 : _T_24108; // @[Mux.scala 31:69:@5394.4]
  assign _T_24110 = valid_16_21 ? 6'h15 : _T_24109; // @[Mux.scala 31:69:@5395.4]
  assign _T_24111 = valid_16_20 ? 6'h14 : _T_24110; // @[Mux.scala 31:69:@5396.4]
  assign _T_24112 = valid_16_19 ? 6'h13 : _T_24111; // @[Mux.scala 31:69:@5397.4]
  assign _T_24113 = valid_16_18 ? 6'h12 : _T_24112; // @[Mux.scala 31:69:@5398.4]
  assign _T_24114 = valid_16_17 ? 6'h11 : _T_24113; // @[Mux.scala 31:69:@5399.4]
  assign _T_24115 = valid_16_16 ? 6'h10 : _T_24114; // @[Mux.scala 31:69:@5400.4]
  assign _T_24116 = valid_16_15 ? 6'hf : _T_24115; // @[Mux.scala 31:69:@5401.4]
  assign _T_24117 = valid_16_14 ? 6'he : _T_24116; // @[Mux.scala 31:69:@5402.4]
  assign _T_24118 = valid_16_13 ? 6'hd : _T_24117; // @[Mux.scala 31:69:@5403.4]
  assign _T_24119 = valid_16_12 ? 6'hc : _T_24118; // @[Mux.scala 31:69:@5404.4]
  assign _T_24120 = valid_16_11 ? 6'hb : _T_24119; // @[Mux.scala 31:69:@5405.4]
  assign _T_24121 = valid_16_10 ? 6'ha : _T_24120; // @[Mux.scala 31:69:@5406.4]
  assign _T_24122 = valid_16_9 ? 6'h9 : _T_24121; // @[Mux.scala 31:69:@5407.4]
  assign _T_24123 = valid_16_8 ? 6'h8 : _T_24122; // @[Mux.scala 31:69:@5408.4]
  assign _T_24124 = valid_16_7 ? 6'h7 : _T_24123; // @[Mux.scala 31:69:@5409.4]
  assign _T_24125 = valid_16_6 ? 6'h6 : _T_24124; // @[Mux.scala 31:69:@5410.4]
  assign _T_24126 = valid_16_5 ? 6'h5 : _T_24125; // @[Mux.scala 31:69:@5411.4]
  assign _T_24127 = valid_16_4 ? 6'h4 : _T_24126; // @[Mux.scala 31:69:@5412.4]
  assign _T_24128 = valid_16_3 ? 6'h3 : _T_24127; // @[Mux.scala 31:69:@5413.4]
  assign _T_24129 = valid_16_2 ? 6'h2 : _T_24128; // @[Mux.scala 31:69:@5414.4]
  assign _T_24130 = valid_16_1 ? 6'h1 : _T_24129; // @[Mux.scala 31:69:@5415.4]
  assign select_16 = valid_16_0 ? 6'h0 : _T_24130; // @[Mux.scala 31:69:@5416.4]
  assign _GEN_1025 = 6'h1 == select_16 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1026 = 6'h2 == select_16 ? io_inData_2 : _GEN_1025; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1027 = 6'h3 == select_16 ? io_inData_3 : _GEN_1026; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1028 = 6'h4 == select_16 ? io_inData_4 : _GEN_1027; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1029 = 6'h5 == select_16 ? io_inData_5 : _GEN_1028; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1030 = 6'h6 == select_16 ? io_inData_6 : _GEN_1029; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1031 = 6'h7 == select_16 ? io_inData_7 : _GEN_1030; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1032 = 6'h8 == select_16 ? io_inData_8 : _GEN_1031; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1033 = 6'h9 == select_16 ? io_inData_9 : _GEN_1032; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1034 = 6'ha == select_16 ? io_inData_10 : _GEN_1033; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1035 = 6'hb == select_16 ? io_inData_11 : _GEN_1034; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1036 = 6'hc == select_16 ? io_inData_12 : _GEN_1035; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1037 = 6'hd == select_16 ? io_inData_13 : _GEN_1036; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1038 = 6'he == select_16 ? io_inData_14 : _GEN_1037; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1039 = 6'hf == select_16 ? io_inData_15 : _GEN_1038; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1040 = 6'h10 == select_16 ? io_inData_16 : _GEN_1039; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1041 = 6'h11 == select_16 ? io_inData_17 : _GEN_1040; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1042 = 6'h12 == select_16 ? io_inData_18 : _GEN_1041; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1043 = 6'h13 == select_16 ? io_inData_19 : _GEN_1042; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1044 = 6'h14 == select_16 ? io_inData_20 : _GEN_1043; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1045 = 6'h15 == select_16 ? io_inData_21 : _GEN_1044; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1046 = 6'h16 == select_16 ? io_inData_22 : _GEN_1045; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1047 = 6'h17 == select_16 ? io_inData_23 : _GEN_1046; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1048 = 6'h18 == select_16 ? io_inData_24 : _GEN_1047; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1049 = 6'h19 == select_16 ? io_inData_25 : _GEN_1048; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1050 = 6'h1a == select_16 ? io_inData_26 : _GEN_1049; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1051 = 6'h1b == select_16 ? io_inData_27 : _GEN_1050; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1052 = 6'h1c == select_16 ? io_inData_28 : _GEN_1051; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1053 = 6'h1d == select_16 ? io_inData_29 : _GEN_1052; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1054 = 6'h1e == select_16 ? io_inData_30 : _GEN_1053; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1055 = 6'h1f == select_16 ? io_inData_31 : _GEN_1054; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1056 = 6'h20 == select_16 ? io_inData_32 : _GEN_1055; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1057 = 6'h21 == select_16 ? io_inData_33 : _GEN_1056; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1058 = 6'h22 == select_16 ? io_inData_34 : _GEN_1057; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1059 = 6'h23 == select_16 ? io_inData_35 : _GEN_1058; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1060 = 6'h24 == select_16 ? io_inData_36 : _GEN_1059; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1061 = 6'h25 == select_16 ? io_inData_37 : _GEN_1060; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1062 = 6'h26 == select_16 ? io_inData_38 : _GEN_1061; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1063 = 6'h27 == select_16 ? io_inData_39 : _GEN_1062; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1064 = 6'h28 == select_16 ? io_inData_40 : _GEN_1063; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1065 = 6'h29 == select_16 ? io_inData_41 : _GEN_1064; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1066 = 6'h2a == select_16 ? io_inData_42 : _GEN_1065; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1067 = 6'h2b == select_16 ? io_inData_43 : _GEN_1066; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1068 = 6'h2c == select_16 ? io_inData_44 : _GEN_1067; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1069 = 6'h2d == select_16 ? io_inData_45 : _GEN_1068; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1070 = 6'h2e == select_16 ? io_inData_46 : _GEN_1069; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1071 = 6'h2f == select_16 ? io_inData_47 : _GEN_1070; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1072 = 6'h30 == select_16 ? io_inData_48 : _GEN_1071; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1073 = 6'h31 == select_16 ? io_inData_49 : _GEN_1072; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1074 = 6'h32 == select_16 ? io_inData_50 : _GEN_1073; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1075 = 6'h33 == select_16 ? io_inData_51 : _GEN_1074; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1076 = 6'h34 == select_16 ? io_inData_52 : _GEN_1075; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1077 = 6'h35 == select_16 ? io_inData_53 : _GEN_1076; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1078 = 6'h36 == select_16 ? io_inData_54 : _GEN_1077; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1079 = 6'h37 == select_16 ? io_inData_55 : _GEN_1078; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1080 = 6'h38 == select_16 ? io_inData_56 : _GEN_1079; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1081 = 6'h39 == select_16 ? io_inData_57 : _GEN_1080; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1082 = 6'h3a == select_16 ? io_inData_58 : _GEN_1081; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1083 = 6'h3b == select_16 ? io_inData_59 : _GEN_1082; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1084 = 6'h3c == select_16 ? io_inData_60 : _GEN_1083; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1085 = 6'h3d == select_16 ? io_inData_61 : _GEN_1084; // @[Switch.scala 33:19:@5418.4]
  assign _GEN_1086 = 6'h3e == select_16 ? io_inData_62 : _GEN_1085; // @[Switch.scala 33:19:@5418.4]
  assign _T_24139 = {valid_16_7,valid_16_6,valid_16_5,valid_16_4,valid_16_3,valid_16_2,valid_16_1,valid_16_0}; // @[Switch.scala 34:32:@5425.4]
  assign _T_24147 = {valid_16_15,valid_16_14,valid_16_13,valid_16_12,valid_16_11,valid_16_10,valid_16_9,valid_16_8,_T_24139}; // @[Switch.scala 34:32:@5433.4]
  assign _T_24154 = {valid_16_23,valid_16_22,valid_16_21,valid_16_20,valid_16_19,valid_16_18,valid_16_17,valid_16_16}; // @[Switch.scala 34:32:@5440.4]
  assign _T_24163 = {valid_16_31,valid_16_30,valid_16_29,valid_16_28,valid_16_27,valid_16_26,valid_16_25,valid_16_24,_T_24154,_T_24147}; // @[Switch.scala 34:32:@5449.4]
  assign _T_24170 = {valid_16_39,valid_16_38,valid_16_37,valid_16_36,valid_16_35,valid_16_34,valid_16_33,valid_16_32}; // @[Switch.scala 34:32:@5456.4]
  assign _T_24178 = {valid_16_47,valid_16_46,valid_16_45,valid_16_44,valid_16_43,valid_16_42,valid_16_41,valid_16_40,_T_24170}; // @[Switch.scala 34:32:@5464.4]
  assign _T_24185 = {valid_16_55,valid_16_54,valid_16_53,valid_16_52,valid_16_51,valid_16_50,valid_16_49,valid_16_48}; // @[Switch.scala 34:32:@5471.4]
  assign _T_24194 = {valid_16_63,valid_16_62,valid_16_61,valid_16_60,valid_16_59,valid_16_58,valid_16_57,valid_16_56,_T_24185,_T_24178}; // @[Switch.scala 34:32:@5480.4]
  assign _T_24195 = {_T_24194,_T_24163}; // @[Switch.scala 34:32:@5481.4]
  assign _T_24199 = io_inAddr_0 == 6'h11; // @[Switch.scala 30:53:@5484.4]
  assign valid_17_0 = io_inValid_0 & _T_24199; // @[Switch.scala 30:36:@5485.4]
  assign _T_24202 = io_inAddr_1 == 6'h11; // @[Switch.scala 30:53:@5487.4]
  assign valid_17_1 = io_inValid_1 & _T_24202; // @[Switch.scala 30:36:@5488.4]
  assign _T_24205 = io_inAddr_2 == 6'h11; // @[Switch.scala 30:53:@5490.4]
  assign valid_17_2 = io_inValid_2 & _T_24205; // @[Switch.scala 30:36:@5491.4]
  assign _T_24208 = io_inAddr_3 == 6'h11; // @[Switch.scala 30:53:@5493.4]
  assign valid_17_3 = io_inValid_3 & _T_24208; // @[Switch.scala 30:36:@5494.4]
  assign _T_24211 = io_inAddr_4 == 6'h11; // @[Switch.scala 30:53:@5496.4]
  assign valid_17_4 = io_inValid_4 & _T_24211; // @[Switch.scala 30:36:@5497.4]
  assign _T_24214 = io_inAddr_5 == 6'h11; // @[Switch.scala 30:53:@5499.4]
  assign valid_17_5 = io_inValid_5 & _T_24214; // @[Switch.scala 30:36:@5500.4]
  assign _T_24217 = io_inAddr_6 == 6'h11; // @[Switch.scala 30:53:@5502.4]
  assign valid_17_6 = io_inValid_6 & _T_24217; // @[Switch.scala 30:36:@5503.4]
  assign _T_24220 = io_inAddr_7 == 6'h11; // @[Switch.scala 30:53:@5505.4]
  assign valid_17_7 = io_inValid_7 & _T_24220; // @[Switch.scala 30:36:@5506.4]
  assign _T_24223 = io_inAddr_8 == 6'h11; // @[Switch.scala 30:53:@5508.4]
  assign valid_17_8 = io_inValid_8 & _T_24223; // @[Switch.scala 30:36:@5509.4]
  assign _T_24226 = io_inAddr_9 == 6'h11; // @[Switch.scala 30:53:@5511.4]
  assign valid_17_9 = io_inValid_9 & _T_24226; // @[Switch.scala 30:36:@5512.4]
  assign _T_24229 = io_inAddr_10 == 6'h11; // @[Switch.scala 30:53:@5514.4]
  assign valid_17_10 = io_inValid_10 & _T_24229; // @[Switch.scala 30:36:@5515.4]
  assign _T_24232 = io_inAddr_11 == 6'h11; // @[Switch.scala 30:53:@5517.4]
  assign valid_17_11 = io_inValid_11 & _T_24232; // @[Switch.scala 30:36:@5518.4]
  assign _T_24235 = io_inAddr_12 == 6'h11; // @[Switch.scala 30:53:@5520.4]
  assign valid_17_12 = io_inValid_12 & _T_24235; // @[Switch.scala 30:36:@5521.4]
  assign _T_24238 = io_inAddr_13 == 6'h11; // @[Switch.scala 30:53:@5523.4]
  assign valid_17_13 = io_inValid_13 & _T_24238; // @[Switch.scala 30:36:@5524.4]
  assign _T_24241 = io_inAddr_14 == 6'h11; // @[Switch.scala 30:53:@5526.4]
  assign valid_17_14 = io_inValid_14 & _T_24241; // @[Switch.scala 30:36:@5527.4]
  assign _T_24244 = io_inAddr_15 == 6'h11; // @[Switch.scala 30:53:@5529.4]
  assign valid_17_15 = io_inValid_15 & _T_24244; // @[Switch.scala 30:36:@5530.4]
  assign _T_24247 = io_inAddr_16 == 6'h11; // @[Switch.scala 30:53:@5532.4]
  assign valid_17_16 = io_inValid_16 & _T_24247; // @[Switch.scala 30:36:@5533.4]
  assign _T_24250 = io_inAddr_17 == 6'h11; // @[Switch.scala 30:53:@5535.4]
  assign valid_17_17 = io_inValid_17 & _T_24250; // @[Switch.scala 30:36:@5536.4]
  assign _T_24253 = io_inAddr_18 == 6'h11; // @[Switch.scala 30:53:@5538.4]
  assign valid_17_18 = io_inValid_18 & _T_24253; // @[Switch.scala 30:36:@5539.4]
  assign _T_24256 = io_inAddr_19 == 6'h11; // @[Switch.scala 30:53:@5541.4]
  assign valid_17_19 = io_inValid_19 & _T_24256; // @[Switch.scala 30:36:@5542.4]
  assign _T_24259 = io_inAddr_20 == 6'h11; // @[Switch.scala 30:53:@5544.4]
  assign valid_17_20 = io_inValid_20 & _T_24259; // @[Switch.scala 30:36:@5545.4]
  assign _T_24262 = io_inAddr_21 == 6'h11; // @[Switch.scala 30:53:@5547.4]
  assign valid_17_21 = io_inValid_21 & _T_24262; // @[Switch.scala 30:36:@5548.4]
  assign _T_24265 = io_inAddr_22 == 6'h11; // @[Switch.scala 30:53:@5550.4]
  assign valid_17_22 = io_inValid_22 & _T_24265; // @[Switch.scala 30:36:@5551.4]
  assign _T_24268 = io_inAddr_23 == 6'h11; // @[Switch.scala 30:53:@5553.4]
  assign valid_17_23 = io_inValid_23 & _T_24268; // @[Switch.scala 30:36:@5554.4]
  assign _T_24271 = io_inAddr_24 == 6'h11; // @[Switch.scala 30:53:@5556.4]
  assign valid_17_24 = io_inValid_24 & _T_24271; // @[Switch.scala 30:36:@5557.4]
  assign _T_24274 = io_inAddr_25 == 6'h11; // @[Switch.scala 30:53:@5559.4]
  assign valid_17_25 = io_inValid_25 & _T_24274; // @[Switch.scala 30:36:@5560.4]
  assign _T_24277 = io_inAddr_26 == 6'h11; // @[Switch.scala 30:53:@5562.4]
  assign valid_17_26 = io_inValid_26 & _T_24277; // @[Switch.scala 30:36:@5563.4]
  assign _T_24280 = io_inAddr_27 == 6'h11; // @[Switch.scala 30:53:@5565.4]
  assign valid_17_27 = io_inValid_27 & _T_24280; // @[Switch.scala 30:36:@5566.4]
  assign _T_24283 = io_inAddr_28 == 6'h11; // @[Switch.scala 30:53:@5568.4]
  assign valid_17_28 = io_inValid_28 & _T_24283; // @[Switch.scala 30:36:@5569.4]
  assign _T_24286 = io_inAddr_29 == 6'h11; // @[Switch.scala 30:53:@5571.4]
  assign valid_17_29 = io_inValid_29 & _T_24286; // @[Switch.scala 30:36:@5572.4]
  assign _T_24289 = io_inAddr_30 == 6'h11; // @[Switch.scala 30:53:@5574.4]
  assign valid_17_30 = io_inValid_30 & _T_24289; // @[Switch.scala 30:36:@5575.4]
  assign _T_24292 = io_inAddr_31 == 6'h11; // @[Switch.scala 30:53:@5577.4]
  assign valid_17_31 = io_inValid_31 & _T_24292; // @[Switch.scala 30:36:@5578.4]
  assign _T_24295 = io_inAddr_32 == 6'h11; // @[Switch.scala 30:53:@5580.4]
  assign valid_17_32 = io_inValid_32 & _T_24295; // @[Switch.scala 30:36:@5581.4]
  assign _T_24298 = io_inAddr_33 == 6'h11; // @[Switch.scala 30:53:@5583.4]
  assign valid_17_33 = io_inValid_33 & _T_24298; // @[Switch.scala 30:36:@5584.4]
  assign _T_24301 = io_inAddr_34 == 6'h11; // @[Switch.scala 30:53:@5586.4]
  assign valid_17_34 = io_inValid_34 & _T_24301; // @[Switch.scala 30:36:@5587.4]
  assign _T_24304 = io_inAddr_35 == 6'h11; // @[Switch.scala 30:53:@5589.4]
  assign valid_17_35 = io_inValid_35 & _T_24304; // @[Switch.scala 30:36:@5590.4]
  assign _T_24307 = io_inAddr_36 == 6'h11; // @[Switch.scala 30:53:@5592.4]
  assign valid_17_36 = io_inValid_36 & _T_24307; // @[Switch.scala 30:36:@5593.4]
  assign _T_24310 = io_inAddr_37 == 6'h11; // @[Switch.scala 30:53:@5595.4]
  assign valid_17_37 = io_inValid_37 & _T_24310; // @[Switch.scala 30:36:@5596.4]
  assign _T_24313 = io_inAddr_38 == 6'h11; // @[Switch.scala 30:53:@5598.4]
  assign valid_17_38 = io_inValid_38 & _T_24313; // @[Switch.scala 30:36:@5599.4]
  assign _T_24316 = io_inAddr_39 == 6'h11; // @[Switch.scala 30:53:@5601.4]
  assign valid_17_39 = io_inValid_39 & _T_24316; // @[Switch.scala 30:36:@5602.4]
  assign _T_24319 = io_inAddr_40 == 6'h11; // @[Switch.scala 30:53:@5604.4]
  assign valid_17_40 = io_inValid_40 & _T_24319; // @[Switch.scala 30:36:@5605.4]
  assign _T_24322 = io_inAddr_41 == 6'h11; // @[Switch.scala 30:53:@5607.4]
  assign valid_17_41 = io_inValid_41 & _T_24322; // @[Switch.scala 30:36:@5608.4]
  assign _T_24325 = io_inAddr_42 == 6'h11; // @[Switch.scala 30:53:@5610.4]
  assign valid_17_42 = io_inValid_42 & _T_24325; // @[Switch.scala 30:36:@5611.4]
  assign _T_24328 = io_inAddr_43 == 6'h11; // @[Switch.scala 30:53:@5613.4]
  assign valid_17_43 = io_inValid_43 & _T_24328; // @[Switch.scala 30:36:@5614.4]
  assign _T_24331 = io_inAddr_44 == 6'h11; // @[Switch.scala 30:53:@5616.4]
  assign valid_17_44 = io_inValid_44 & _T_24331; // @[Switch.scala 30:36:@5617.4]
  assign _T_24334 = io_inAddr_45 == 6'h11; // @[Switch.scala 30:53:@5619.4]
  assign valid_17_45 = io_inValid_45 & _T_24334; // @[Switch.scala 30:36:@5620.4]
  assign _T_24337 = io_inAddr_46 == 6'h11; // @[Switch.scala 30:53:@5622.4]
  assign valid_17_46 = io_inValid_46 & _T_24337; // @[Switch.scala 30:36:@5623.4]
  assign _T_24340 = io_inAddr_47 == 6'h11; // @[Switch.scala 30:53:@5625.4]
  assign valid_17_47 = io_inValid_47 & _T_24340; // @[Switch.scala 30:36:@5626.4]
  assign _T_24343 = io_inAddr_48 == 6'h11; // @[Switch.scala 30:53:@5628.4]
  assign valid_17_48 = io_inValid_48 & _T_24343; // @[Switch.scala 30:36:@5629.4]
  assign _T_24346 = io_inAddr_49 == 6'h11; // @[Switch.scala 30:53:@5631.4]
  assign valid_17_49 = io_inValid_49 & _T_24346; // @[Switch.scala 30:36:@5632.4]
  assign _T_24349 = io_inAddr_50 == 6'h11; // @[Switch.scala 30:53:@5634.4]
  assign valid_17_50 = io_inValid_50 & _T_24349; // @[Switch.scala 30:36:@5635.4]
  assign _T_24352 = io_inAddr_51 == 6'h11; // @[Switch.scala 30:53:@5637.4]
  assign valid_17_51 = io_inValid_51 & _T_24352; // @[Switch.scala 30:36:@5638.4]
  assign _T_24355 = io_inAddr_52 == 6'h11; // @[Switch.scala 30:53:@5640.4]
  assign valid_17_52 = io_inValid_52 & _T_24355; // @[Switch.scala 30:36:@5641.4]
  assign _T_24358 = io_inAddr_53 == 6'h11; // @[Switch.scala 30:53:@5643.4]
  assign valid_17_53 = io_inValid_53 & _T_24358; // @[Switch.scala 30:36:@5644.4]
  assign _T_24361 = io_inAddr_54 == 6'h11; // @[Switch.scala 30:53:@5646.4]
  assign valid_17_54 = io_inValid_54 & _T_24361; // @[Switch.scala 30:36:@5647.4]
  assign _T_24364 = io_inAddr_55 == 6'h11; // @[Switch.scala 30:53:@5649.4]
  assign valid_17_55 = io_inValid_55 & _T_24364; // @[Switch.scala 30:36:@5650.4]
  assign _T_24367 = io_inAddr_56 == 6'h11; // @[Switch.scala 30:53:@5652.4]
  assign valid_17_56 = io_inValid_56 & _T_24367; // @[Switch.scala 30:36:@5653.4]
  assign _T_24370 = io_inAddr_57 == 6'h11; // @[Switch.scala 30:53:@5655.4]
  assign valid_17_57 = io_inValid_57 & _T_24370; // @[Switch.scala 30:36:@5656.4]
  assign _T_24373 = io_inAddr_58 == 6'h11; // @[Switch.scala 30:53:@5658.4]
  assign valid_17_58 = io_inValid_58 & _T_24373; // @[Switch.scala 30:36:@5659.4]
  assign _T_24376 = io_inAddr_59 == 6'h11; // @[Switch.scala 30:53:@5661.4]
  assign valid_17_59 = io_inValid_59 & _T_24376; // @[Switch.scala 30:36:@5662.4]
  assign _T_24379 = io_inAddr_60 == 6'h11; // @[Switch.scala 30:53:@5664.4]
  assign valid_17_60 = io_inValid_60 & _T_24379; // @[Switch.scala 30:36:@5665.4]
  assign _T_24382 = io_inAddr_61 == 6'h11; // @[Switch.scala 30:53:@5667.4]
  assign valid_17_61 = io_inValid_61 & _T_24382; // @[Switch.scala 30:36:@5668.4]
  assign _T_24385 = io_inAddr_62 == 6'h11; // @[Switch.scala 30:53:@5670.4]
  assign valid_17_62 = io_inValid_62 & _T_24385; // @[Switch.scala 30:36:@5671.4]
  assign _T_24388 = io_inAddr_63 == 6'h11; // @[Switch.scala 30:53:@5673.4]
  assign valid_17_63 = io_inValid_63 & _T_24388; // @[Switch.scala 30:36:@5674.4]
  assign _T_24454 = valid_17_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@5676.4]
  assign _T_24455 = valid_17_61 ? 6'h3d : _T_24454; // @[Mux.scala 31:69:@5677.4]
  assign _T_24456 = valid_17_60 ? 6'h3c : _T_24455; // @[Mux.scala 31:69:@5678.4]
  assign _T_24457 = valid_17_59 ? 6'h3b : _T_24456; // @[Mux.scala 31:69:@5679.4]
  assign _T_24458 = valid_17_58 ? 6'h3a : _T_24457; // @[Mux.scala 31:69:@5680.4]
  assign _T_24459 = valid_17_57 ? 6'h39 : _T_24458; // @[Mux.scala 31:69:@5681.4]
  assign _T_24460 = valid_17_56 ? 6'h38 : _T_24459; // @[Mux.scala 31:69:@5682.4]
  assign _T_24461 = valid_17_55 ? 6'h37 : _T_24460; // @[Mux.scala 31:69:@5683.4]
  assign _T_24462 = valid_17_54 ? 6'h36 : _T_24461; // @[Mux.scala 31:69:@5684.4]
  assign _T_24463 = valid_17_53 ? 6'h35 : _T_24462; // @[Mux.scala 31:69:@5685.4]
  assign _T_24464 = valid_17_52 ? 6'h34 : _T_24463; // @[Mux.scala 31:69:@5686.4]
  assign _T_24465 = valid_17_51 ? 6'h33 : _T_24464; // @[Mux.scala 31:69:@5687.4]
  assign _T_24466 = valid_17_50 ? 6'h32 : _T_24465; // @[Mux.scala 31:69:@5688.4]
  assign _T_24467 = valid_17_49 ? 6'h31 : _T_24466; // @[Mux.scala 31:69:@5689.4]
  assign _T_24468 = valid_17_48 ? 6'h30 : _T_24467; // @[Mux.scala 31:69:@5690.4]
  assign _T_24469 = valid_17_47 ? 6'h2f : _T_24468; // @[Mux.scala 31:69:@5691.4]
  assign _T_24470 = valid_17_46 ? 6'h2e : _T_24469; // @[Mux.scala 31:69:@5692.4]
  assign _T_24471 = valid_17_45 ? 6'h2d : _T_24470; // @[Mux.scala 31:69:@5693.4]
  assign _T_24472 = valid_17_44 ? 6'h2c : _T_24471; // @[Mux.scala 31:69:@5694.4]
  assign _T_24473 = valid_17_43 ? 6'h2b : _T_24472; // @[Mux.scala 31:69:@5695.4]
  assign _T_24474 = valid_17_42 ? 6'h2a : _T_24473; // @[Mux.scala 31:69:@5696.4]
  assign _T_24475 = valid_17_41 ? 6'h29 : _T_24474; // @[Mux.scala 31:69:@5697.4]
  assign _T_24476 = valid_17_40 ? 6'h28 : _T_24475; // @[Mux.scala 31:69:@5698.4]
  assign _T_24477 = valid_17_39 ? 6'h27 : _T_24476; // @[Mux.scala 31:69:@5699.4]
  assign _T_24478 = valid_17_38 ? 6'h26 : _T_24477; // @[Mux.scala 31:69:@5700.4]
  assign _T_24479 = valid_17_37 ? 6'h25 : _T_24478; // @[Mux.scala 31:69:@5701.4]
  assign _T_24480 = valid_17_36 ? 6'h24 : _T_24479; // @[Mux.scala 31:69:@5702.4]
  assign _T_24481 = valid_17_35 ? 6'h23 : _T_24480; // @[Mux.scala 31:69:@5703.4]
  assign _T_24482 = valid_17_34 ? 6'h22 : _T_24481; // @[Mux.scala 31:69:@5704.4]
  assign _T_24483 = valid_17_33 ? 6'h21 : _T_24482; // @[Mux.scala 31:69:@5705.4]
  assign _T_24484 = valid_17_32 ? 6'h20 : _T_24483; // @[Mux.scala 31:69:@5706.4]
  assign _T_24485 = valid_17_31 ? 6'h1f : _T_24484; // @[Mux.scala 31:69:@5707.4]
  assign _T_24486 = valid_17_30 ? 6'h1e : _T_24485; // @[Mux.scala 31:69:@5708.4]
  assign _T_24487 = valid_17_29 ? 6'h1d : _T_24486; // @[Mux.scala 31:69:@5709.4]
  assign _T_24488 = valid_17_28 ? 6'h1c : _T_24487; // @[Mux.scala 31:69:@5710.4]
  assign _T_24489 = valid_17_27 ? 6'h1b : _T_24488; // @[Mux.scala 31:69:@5711.4]
  assign _T_24490 = valid_17_26 ? 6'h1a : _T_24489; // @[Mux.scala 31:69:@5712.4]
  assign _T_24491 = valid_17_25 ? 6'h19 : _T_24490; // @[Mux.scala 31:69:@5713.4]
  assign _T_24492 = valid_17_24 ? 6'h18 : _T_24491; // @[Mux.scala 31:69:@5714.4]
  assign _T_24493 = valid_17_23 ? 6'h17 : _T_24492; // @[Mux.scala 31:69:@5715.4]
  assign _T_24494 = valid_17_22 ? 6'h16 : _T_24493; // @[Mux.scala 31:69:@5716.4]
  assign _T_24495 = valid_17_21 ? 6'h15 : _T_24494; // @[Mux.scala 31:69:@5717.4]
  assign _T_24496 = valid_17_20 ? 6'h14 : _T_24495; // @[Mux.scala 31:69:@5718.4]
  assign _T_24497 = valid_17_19 ? 6'h13 : _T_24496; // @[Mux.scala 31:69:@5719.4]
  assign _T_24498 = valid_17_18 ? 6'h12 : _T_24497; // @[Mux.scala 31:69:@5720.4]
  assign _T_24499 = valid_17_17 ? 6'h11 : _T_24498; // @[Mux.scala 31:69:@5721.4]
  assign _T_24500 = valid_17_16 ? 6'h10 : _T_24499; // @[Mux.scala 31:69:@5722.4]
  assign _T_24501 = valid_17_15 ? 6'hf : _T_24500; // @[Mux.scala 31:69:@5723.4]
  assign _T_24502 = valid_17_14 ? 6'he : _T_24501; // @[Mux.scala 31:69:@5724.4]
  assign _T_24503 = valid_17_13 ? 6'hd : _T_24502; // @[Mux.scala 31:69:@5725.4]
  assign _T_24504 = valid_17_12 ? 6'hc : _T_24503; // @[Mux.scala 31:69:@5726.4]
  assign _T_24505 = valid_17_11 ? 6'hb : _T_24504; // @[Mux.scala 31:69:@5727.4]
  assign _T_24506 = valid_17_10 ? 6'ha : _T_24505; // @[Mux.scala 31:69:@5728.4]
  assign _T_24507 = valid_17_9 ? 6'h9 : _T_24506; // @[Mux.scala 31:69:@5729.4]
  assign _T_24508 = valid_17_8 ? 6'h8 : _T_24507; // @[Mux.scala 31:69:@5730.4]
  assign _T_24509 = valid_17_7 ? 6'h7 : _T_24508; // @[Mux.scala 31:69:@5731.4]
  assign _T_24510 = valid_17_6 ? 6'h6 : _T_24509; // @[Mux.scala 31:69:@5732.4]
  assign _T_24511 = valid_17_5 ? 6'h5 : _T_24510; // @[Mux.scala 31:69:@5733.4]
  assign _T_24512 = valid_17_4 ? 6'h4 : _T_24511; // @[Mux.scala 31:69:@5734.4]
  assign _T_24513 = valid_17_3 ? 6'h3 : _T_24512; // @[Mux.scala 31:69:@5735.4]
  assign _T_24514 = valid_17_2 ? 6'h2 : _T_24513; // @[Mux.scala 31:69:@5736.4]
  assign _T_24515 = valid_17_1 ? 6'h1 : _T_24514; // @[Mux.scala 31:69:@5737.4]
  assign select_17 = valid_17_0 ? 6'h0 : _T_24515; // @[Mux.scala 31:69:@5738.4]
  assign _GEN_1089 = 6'h1 == select_17 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1090 = 6'h2 == select_17 ? io_inData_2 : _GEN_1089; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1091 = 6'h3 == select_17 ? io_inData_3 : _GEN_1090; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1092 = 6'h4 == select_17 ? io_inData_4 : _GEN_1091; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1093 = 6'h5 == select_17 ? io_inData_5 : _GEN_1092; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1094 = 6'h6 == select_17 ? io_inData_6 : _GEN_1093; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1095 = 6'h7 == select_17 ? io_inData_7 : _GEN_1094; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1096 = 6'h8 == select_17 ? io_inData_8 : _GEN_1095; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1097 = 6'h9 == select_17 ? io_inData_9 : _GEN_1096; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1098 = 6'ha == select_17 ? io_inData_10 : _GEN_1097; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1099 = 6'hb == select_17 ? io_inData_11 : _GEN_1098; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1100 = 6'hc == select_17 ? io_inData_12 : _GEN_1099; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1101 = 6'hd == select_17 ? io_inData_13 : _GEN_1100; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1102 = 6'he == select_17 ? io_inData_14 : _GEN_1101; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1103 = 6'hf == select_17 ? io_inData_15 : _GEN_1102; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1104 = 6'h10 == select_17 ? io_inData_16 : _GEN_1103; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1105 = 6'h11 == select_17 ? io_inData_17 : _GEN_1104; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1106 = 6'h12 == select_17 ? io_inData_18 : _GEN_1105; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1107 = 6'h13 == select_17 ? io_inData_19 : _GEN_1106; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1108 = 6'h14 == select_17 ? io_inData_20 : _GEN_1107; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1109 = 6'h15 == select_17 ? io_inData_21 : _GEN_1108; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1110 = 6'h16 == select_17 ? io_inData_22 : _GEN_1109; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1111 = 6'h17 == select_17 ? io_inData_23 : _GEN_1110; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1112 = 6'h18 == select_17 ? io_inData_24 : _GEN_1111; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1113 = 6'h19 == select_17 ? io_inData_25 : _GEN_1112; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1114 = 6'h1a == select_17 ? io_inData_26 : _GEN_1113; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1115 = 6'h1b == select_17 ? io_inData_27 : _GEN_1114; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1116 = 6'h1c == select_17 ? io_inData_28 : _GEN_1115; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1117 = 6'h1d == select_17 ? io_inData_29 : _GEN_1116; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1118 = 6'h1e == select_17 ? io_inData_30 : _GEN_1117; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1119 = 6'h1f == select_17 ? io_inData_31 : _GEN_1118; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1120 = 6'h20 == select_17 ? io_inData_32 : _GEN_1119; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1121 = 6'h21 == select_17 ? io_inData_33 : _GEN_1120; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1122 = 6'h22 == select_17 ? io_inData_34 : _GEN_1121; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1123 = 6'h23 == select_17 ? io_inData_35 : _GEN_1122; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1124 = 6'h24 == select_17 ? io_inData_36 : _GEN_1123; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1125 = 6'h25 == select_17 ? io_inData_37 : _GEN_1124; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1126 = 6'h26 == select_17 ? io_inData_38 : _GEN_1125; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1127 = 6'h27 == select_17 ? io_inData_39 : _GEN_1126; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1128 = 6'h28 == select_17 ? io_inData_40 : _GEN_1127; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1129 = 6'h29 == select_17 ? io_inData_41 : _GEN_1128; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1130 = 6'h2a == select_17 ? io_inData_42 : _GEN_1129; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1131 = 6'h2b == select_17 ? io_inData_43 : _GEN_1130; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1132 = 6'h2c == select_17 ? io_inData_44 : _GEN_1131; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1133 = 6'h2d == select_17 ? io_inData_45 : _GEN_1132; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1134 = 6'h2e == select_17 ? io_inData_46 : _GEN_1133; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1135 = 6'h2f == select_17 ? io_inData_47 : _GEN_1134; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1136 = 6'h30 == select_17 ? io_inData_48 : _GEN_1135; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1137 = 6'h31 == select_17 ? io_inData_49 : _GEN_1136; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1138 = 6'h32 == select_17 ? io_inData_50 : _GEN_1137; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1139 = 6'h33 == select_17 ? io_inData_51 : _GEN_1138; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1140 = 6'h34 == select_17 ? io_inData_52 : _GEN_1139; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1141 = 6'h35 == select_17 ? io_inData_53 : _GEN_1140; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1142 = 6'h36 == select_17 ? io_inData_54 : _GEN_1141; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1143 = 6'h37 == select_17 ? io_inData_55 : _GEN_1142; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1144 = 6'h38 == select_17 ? io_inData_56 : _GEN_1143; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1145 = 6'h39 == select_17 ? io_inData_57 : _GEN_1144; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1146 = 6'h3a == select_17 ? io_inData_58 : _GEN_1145; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1147 = 6'h3b == select_17 ? io_inData_59 : _GEN_1146; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1148 = 6'h3c == select_17 ? io_inData_60 : _GEN_1147; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1149 = 6'h3d == select_17 ? io_inData_61 : _GEN_1148; // @[Switch.scala 33:19:@5740.4]
  assign _GEN_1150 = 6'h3e == select_17 ? io_inData_62 : _GEN_1149; // @[Switch.scala 33:19:@5740.4]
  assign _T_24524 = {valid_17_7,valid_17_6,valid_17_5,valid_17_4,valid_17_3,valid_17_2,valid_17_1,valid_17_0}; // @[Switch.scala 34:32:@5747.4]
  assign _T_24532 = {valid_17_15,valid_17_14,valid_17_13,valid_17_12,valid_17_11,valid_17_10,valid_17_9,valid_17_8,_T_24524}; // @[Switch.scala 34:32:@5755.4]
  assign _T_24539 = {valid_17_23,valid_17_22,valid_17_21,valid_17_20,valid_17_19,valid_17_18,valid_17_17,valid_17_16}; // @[Switch.scala 34:32:@5762.4]
  assign _T_24548 = {valid_17_31,valid_17_30,valid_17_29,valid_17_28,valid_17_27,valid_17_26,valid_17_25,valid_17_24,_T_24539,_T_24532}; // @[Switch.scala 34:32:@5771.4]
  assign _T_24555 = {valid_17_39,valid_17_38,valid_17_37,valid_17_36,valid_17_35,valid_17_34,valid_17_33,valid_17_32}; // @[Switch.scala 34:32:@5778.4]
  assign _T_24563 = {valid_17_47,valid_17_46,valid_17_45,valid_17_44,valid_17_43,valid_17_42,valid_17_41,valid_17_40,_T_24555}; // @[Switch.scala 34:32:@5786.4]
  assign _T_24570 = {valid_17_55,valid_17_54,valid_17_53,valid_17_52,valid_17_51,valid_17_50,valid_17_49,valid_17_48}; // @[Switch.scala 34:32:@5793.4]
  assign _T_24579 = {valid_17_63,valid_17_62,valid_17_61,valid_17_60,valid_17_59,valid_17_58,valid_17_57,valid_17_56,_T_24570,_T_24563}; // @[Switch.scala 34:32:@5802.4]
  assign _T_24580 = {_T_24579,_T_24548}; // @[Switch.scala 34:32:@5803.4]
  assign _T_24584 = io_inAddr_0 == 6'h12; // @[Switch.scala 30:53:@5806.4]
  assign valid_18_0 = io_inValid_0 & _T_24584; // @[Switch.scala 30:36:@5807.4]
  assign _T_24587 = io_inAddr_1 == 6'h12; // @[Switch.scala 30:53:@5809.4]
  assign valid_18_1 = io_inValid_1 & _T_24587; // @[Switch.scala 30:36:@5810.4]
  assign _T_24590 = io_inAddr_2 == 6'h12; // @[Switch.scala 30:53:@5812.4]
  assign valid_18_2 = io_inValid_2 & _T_24590; // @[Switch.scala 30:36:@5813.4]
  assign _T_24593 = io_inAddr_3 == 6'h12; // @[Switch.scala 30:53:@5815.4]
  assign valid_18_3 = io_inValid_3 & _T_24593; // @[Switch.scala 30:36:@5816.4]
  assign _T_24596 = io_inAddr_4 == 6'h12; // @[Switch.scala 30:53:@5818.4]
  assign valid_18_4 = io_inValid_4 & _T_24596; // @[Switch.scala 30:36:@5819.4]
  assign _T_24599 = io_inAddr_5 == 6'h12; // @[Switch.scala 30:53:@5821.4]
  assign valid_18_5 = io_inValid_5 & _T_24599; // @[Switch.scala 30:36:@5822.4]
  assign _T_24602 = io_inAddr_6 == 6'h12; // @[Switch.scala 30:53:@5824.4]
  assign valid_18_6 = io_inValid_6 & _T_24602; // @[Switch.scala 30:36:@5825.4]
  assign _T_24605 = io_inAddr_7 == 6'h12; // @[Switch.scala 30:53:@5827.4]
  assign valid_18_7 = io_inValid_7 & _T_24605; // @[Switch.scala 30:36:@5828.4]
  assign _T_24608 = io_inAddr_8 == 6'h12; // @[Switch.scala 30:53:@5830.4]
  assign valid_18_8 = io_inValid_8 & _T_24608; // @[Switch.scala 30:36:@5831.4]
  assign _T_24611 = io_inAddr_9 == 6'h12; // @[Switch.scala 30:53:@5833.4]
  assign valid_18_9 = io_inValid_9 & _T_24611; // @[Switch.scala 30:36:@5834.4]
  assign _T_24614 = io_inAddr_10 == 6'h12; // @[Switch.scala 30:53:@5836.4]
  assign valid_18_10 = io_inValid_10 & _T_24614; // @[Switch.scala 30:36:@5837.4]
  assign _T_24617 = io_inAddr_11 == 6'h12; // @[Switch.scala 30:53:@5839.4]
  assign valid_18_11 = io_inValid_11 & _T_24617; // @[Switch.scala 30:36:@5840.4]
  assign _T_24620 = io_inAddr_12 == 6'h12; // @[Switch.scala 30:53:@5842.4]
  assign valid_18_12 = io_inValid_12 & _T_24620; // @[Switch.scala 30:36:@5843.4]
  assign _T_24623 = io_inAddr_13 == 6'h12; // @[Switch.scala 30:53:@5845.4]
  assign valid_18_13 = io_inValid_13 & _T_24623; // @[Switch.scala 30:36:@5846.4]
  assign _T_24626 = io_inAddr_14 == 6'h12; // @[Switch.scala 30:53:@5848.4]
  assign valid_18_14 = io_inValid_14 & _T_24626; // @[Switch.scala 30:36:@5849.4]
  assign _T_24629 = io_inAddr_15 == 6'h12; // @[Switch.scala 30:53:@5851.4]
  assign valid_18_15 = io_inValid_15 & _T_24629; // @[Switch.scala 30:36:@5852.4]
  assign _T_24632 = io_inAddr_16 == 6'h12; // @[Switch.scala 30:53:@5854.4]
  assign valid_18_16 = io_inValid_16 & _T_24632; // @[Switch.scala 30:36:@5855.4]
  assign _T_24635 = io_inAddr_17 == 6'h12; // @[Switch.scala 30:53:@5857.4]
  assign valid_18_17 = io_inValid_17 & _T_24635; // @[Switch.scala 30:36:@5858.4]
  assign _T_24638 = io_inAddr_18 == 6'h12; // @[Switch.scala 30:53:@5860.4]
  assign valid_18_18 = io_inValid_18 & _T_24638; // @[Switch.scala 30:36:@5861.4]
  assign _T_24641 = io_inAddr_19 == 6'h12; // @[Switch.scala 30:53:@5863.4]
  assign valid_18_19 = io_inValid_19 & _T_24641; // @[Switch.scala 30:36:@5864.4]
  assign _T_24644 = io_inAddr_20 == 6'h12; // @[Switch.scala 30:53:@5866.4]
  assign valid_18_20 = io_inValid_20 & _T_24644; // @[Switch.scala 30:36:@5867.4]
  assign _T_24647 = io_inAddr_21 == 6'h12; // @[Switch.scala 30:53:@5869.4]
  assign valid_18_21 = io_inValid_21 & _T_24647; // @[Switch.scala 30:36:@5870.4]
  assign _T_24650 = io_inAddr_22 == 6'h12; // @[Switch.scala 30:53:@5872.4]
  assign valid_18_22 = io_inValid_22 & _T_24650; // @[Switch.scala 30:36:@5873.4]
  assign _T_24653 = io_inAddr_23 == 6'h12; // @[Switch.scala 30:53:@5875.4]
  assign valid_18_23 = io_inValid_23 & _T_24653; // @[Switch.scala 30:36:@5876.4]
  assign _T_24656 = io_inAddr_24 == 6'h12; // @[Switch.scala 30:53:@5878.4]
  assign valid_18_24 = io_inValid_24 & _T_24656; // @[Switch.scala 30:36:@5879.4]
  assign _T_24659 = io_inAddr_25 == 6'h12; // @[Switch.scala 30:53:@5881.4]
  assign valid_18_25 = io_inValid_25 & _T_24659; // @[Switch.scala 30:36:@5882.4]
  assign _T_24662 = io_inAddr_26 == 6'h12; // @[Switch.scala 30:53:@5884.4]
  assign valid_18_26 = io_inValid_26 & _T_24662; // @[Switch.scala 30:36:@5885.4]
  assign _T_24665 = io_inAddr_27 == 6'h12; // @[Switch.scala 30:53:@5887.4]
  assign valid_18_27 = io_inValid_27 & _T_24665; // @[Switch.scala 30:36:@5888.4]
  assign _T_24668 = io_inAddr_28 == 6'h12; // @[Switch.scala 30:53:@5890.4]
  assign valid_18_28 = io_inValid_28 & _T_24668; // @[Switch.scala 30:36:@5891.4]
  assign _T_24671 = io_inAddr_29 == 6'h12; // @[Switch.scala 30:53:@5893.4]
  assign valid_18_29 = io_inValid_29 & _T_24671; // @[Switch.scala 30:36:@5894.4]
  assign _T_24674 = io_inAddr_30 == 6'h12; // @[Switch.scala 30:53:@5896.4]
  assign valid_18_30 = io_inValid_30 & _T_24674; // @[Switch.scala 30:36:@5897.4]
  assign _T_24677 = io_inAddr_31 == 6'h12; // @[Switch.scala 30:53:@5899.4]
  assign valid_18_31 = io_inValid_31 & _T_24677; // @[Switch.scala 30:36:@5900.4]
  assign _T_24680 = io_inAddr_32 == 6'h12; // @[Switch.scala 30:53:@5902.4]
  assign valid_18_32 = io_inValid_32 & _T_24680; // @[Switch.scala 30:36:@5903.4]
  assign _T_24683 = io_inAddr_33 == 6'h12; // @[Switch.scala 30:53:@5905.4]
  assign valid_18_33 = io_inValid_33 & _T_24683; // @[Switch.scala 30:36:@5906.4]
  assign _T_24686 = io_inAddr_34 == 6'h12; // @[Switch.scala 30:53:@5908.4]
  assign valid_18_34 = io_inValid_34 & _T_24686; // @[Switch.scala 30:36:@5909.4]
  assign _T_24689 = io_inAddr_35 == 6'h12; // @[Switch.scala 30:53:@5911.4]
  assign valid_18_35 = io_inValid_35 & _T_24689; // @[Switch.scala 30:36:@5912.4]
  assign _T_24692 = io_inAddr_36 == 6'h12; // @[Switch.scala 30:53:@5914.4]
  assign valid_18_36 = io_inValid_36 & _T_24692; // @[Switch.scala 30:36:@5915.4]
  assign _T_24695 = io_inAddr_37 == 6'h12; // @[Switch.scala 30:53:@5917.4]
  assign valid_18_37 = io_inValid_37 & _T_24695; // @[Switch.scala 30:36:@5918.4]
  assign _T_24698 = io_inAddr_38 == 6'h12; // @[Switch.scala 30:53:@5920.4]
  assign valid_18_38 = io_inValid_38 & _T_24698; // @[Switch.scala 30:36:@5921.4]
  assign _T_24701 = io_inAddr_39 == 6'h12; // @[Switch.scala 30:53:@5923.4]
  assign valid_18_39 = io_inValid_39 & _T_24701; // @[Switch.scala 30:36:@5924.4]
  assign _T_24704 = io_inAddr_40 == 6'h12; // @[Switch.scala 30:53:@5926.4]
  assign valid_18_40 = io_inValid_40 & _T_24704; // @[Switch.scala 30:36:@5927.4]
  assign _T_24707 = io_inAddr_41 == 6'h12; // @[Switch.scala 30:53:@5929.4]
  assign valid_18_41 = io_inValid_41 & _T_24707; // @[Switch.scala 30:36:@5930.4]
  assign _T_24710 = io_inAddr_42 == 6'h12; // @[Switch.scala 30:53:@5932.4]
  assign valid_18_42 = io_inValid_42 & _T_24710; // @[Switch.scala 30:36:@5933.4]
  assign _T_24713 = io_inAddr_43 == 6'h12; // @[Switch.scala 30:53:@5935.4]
  assign valid_18_43 = io_inValid_43 & _T_24713; // @[Switch.scala 30:36:@5936.4]
  assign _T_24716 = io_inAddr_44 == 6'h12; // @[Switch.scala 30:53:@5938.4]
  assign valid_18_44 = io_inValid_44 & _T_24716; // @[Switch.scala 30:36:@5939.4]
  assign _T_24719 = io_inAddr_45 == 6'h12; // @[Switch.scala 30:53:@5941.4]
  assign valid_18_45 = io_inValid_45 & _T_24719; // @[Switch.scala 30:36:@5942.4]
  assign _T_24722 = io_inAddr_46 == 6'h12; // @[Switch.scala 30:53:@5944.4]
  assign valid_18_46 = io_inValid_46 & _T_24722; // @[Switch.scala 30:36:@5945.4]
  assign _T_24725 = io_inAddr_47 == 6'h12; // @[Switch.scala 30:53:@5947.4]
  assign valid_18_47 = io_inValid_47 & _T_24725; // @[Switch.scala 30:36:@5948.4]
  assign _T_24728 = io_inAddr_48 == 6'h12; // @[Switch.scala 30:53:@5950.4]
  assign valid_18_48 = io_inValid_48 & _T_24728; // @[Switch.scala 30:36:@5951.4]
  assign _T_24731 = io_inAddr_49 == 6'h12; // @[Switch.scala 30:53:@5953.4]
  assign valid_18_49 = io_inValid_49 & _T_24731; // @[Switch.scala 30:36:@5954.4]
  assign _T_24734 = io_inAddr_50 == 6'h12; // @[Switch.scala 30:53:@5956.4]
  assign valid_18_50 = io_inValid_50 & _T_24734; // @[Switch.scala 30:36:@5957.4]
  assign _T_24737 = io_inAddr_51 == 6'h12; // @[Switch.scala 30:53:@5959.4]
  assign valid_18_51 = io_inValid_51 & _T_24737; // @[Switch.scala 30:36:@5960.4]
  assign _T_24740 = io_inAddr_52 == 6'h12; // @[Switch.scala 30:53:@5962.4]
  assign valid_18_52 = io_inValid_52 & _T_24740; // @[Switch.scala 30:36:@5963.4]
  assign _T_24743 = io_inAddr_53 == 6'h12; // @[Switch.scala 30:53:@5965.4]
  assign valid_18_53 = io_inValid_53 & _T_24743; // @[Switch.scala 30:36:@5966.4]
  assign _T_24746 = io_inAddr_54 == 6'h12; // @[Switch.scala 30:53:@5968.4]
  assign valid_18_54 = io_inValid_54 & _T_24746; // @[Switch.scala 30:36:@5969.4]
  assign _T_24749 = io_inAddr_55 == 6'h12; // @[Switch.scala 30:53:@5971.4]
  assign valid_18_55 = io_inValid_55 & _T_24749; // @[Switch.scala 30:36:@5972.4]
  assign _T_24752 = io_inAddr_56 == 6'h12; // @[Switch.scala 30:53:@5974.4]
  assign valid_18_56 = io_inValid_56 & _T_24752; // @[Switch.scala 30:36:@5975.4]
  assign _T_24755 = io_inAddr_57 == 6'h12; // @[Switch.scala 30:53:@5977.4]
  assign valid_18_57 = io_inValid_57 & _T_24755; // @[Switch.scala 30:36:@5978.4]
  assign _T_24758 = io_inAddr_58 == 6'h12; // @[Switch.scala 30:53:@5980.4]
  assign valid_18_58 = io_inValid_58 & _T_24758; // @[Switch.scala 30:36:@5981.4]
  assign _T_24761 = io_inAddr_59 == 6'h12; // @[Switch.scala 30:53:@5983.4]
  assign valid_18_59 = io_inValid_59 & _T_24761; // @[Switch.scala 30:36:@5984.4]
  assign _T_24764 = io_inAddr_60 == 6'h12; // @[Switch.scala 30:53:@5986.4]
  assign valid_18_60 = io_inValid_60 & _T_24764; // @[Switch.scala 30:36:@5987.4]
  assign _T_24767 = io_inAddr_61 == 6'h12; // @[Switch.scala 30:53:@5989.4]
  assign valid_18_61 = io_inValid_61 & _T_24767; // @[Switch.scala 30:36:@5990.4]
  assign _T_24770 = io_inAddr_62 == 6'h12; // @[Switch.scala 30:53:@5992.4]
  assign valid_18_62 = io_inValid_62 & _T_24770; // @[Switch.scala 30:36:@5993.4]
  assign _T_24773 = io_inAddr_63 == 6'h12; // @[Switch.scala 30:53:@5995.4]
  assign valid_18_63 = io_inValid_63 & _T_24773; // @[Switch.scala 30:36:@5996.4]
  assign _T_24839 = valid_18_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@5998.4]
  assign _T_24840 = valid_18_61 ? 6'h3d : _T_24839; // @[Mux.scala 31:69:@5999.4]
  assign _T_24841 = valid_18_60 ? 6'h3c : _T_24840; // @[Mux.scala 31:69:@6000.4]
  assign _T_24842 = valid_18_59 ? 6'h3b : _T_24841; // @[Mux.scala 31:69:@6001.4]
  assign _T_24843 = valid_18_58 ? 6'h3a : _T_24842; // @[Mux.scala 31:69:@6002.4]
  assign _T_24844 = valid_18_57 ? 6'h39 : _T_24843; // @[Mux.scala 31:69:@6003.4]
  assign _T_24845 = valid_18_56 ? 6'h38 : _T_24844; // @[Mux.scala 31:69:@6004.4]
  assign _T_24846 = valid_18_55 ? 6'h37 : _T_24845; // @[Mux.scala 31:69:@6005.4]
  assign _T_24847 = valid_18_54 ? 6'h36 : _T_24846; // @[Mux.scala 31:69:@6006.4]
  assign _T_24848 = valid_18_53 ? 6'h35 : _T_24847; // @[Mux.scala 31:69:@6007.4]
  assign _T_24849 = valid_18_52 ? 6'h34 : _T_24848; // @[Mux.scala 31:69:@6008.4]
  assign _T_24850 = valid_18_51 ? 6'h33 : _T_24849; // @[Mux.scala 31:69:@6009.4]
  assign _T_24851 = valid_18_50 ? 6'h32 : _T_24850; // @[Mux.scala 31:69:@6010.4]
  assign _T_24852 = valid_18_49 ? 6'h31 : _T_24851; // @[Mux.scala 31:69:@6011.4]
  assign _T_24853 = valid_18_48 ? 6'h30 : _T_24852; // @[Mux.scala 31:69:@6012.4]
  assign _T_24854 = valid_18_47 ? 6'h2f : _T_24853; // @[Mux.scala 31:69:@6013.4]
  assign _T_24855 = valid_18_46 ? 6'h2e : _T_24854; // @[Mux.scala 31:69:@6014.4]
  assign _T_24856 = valid_18_45 ? 6'h2d : _T_24855; // @[Mux.scala 31:69:@6015.4]
  assign _T_24857 = valid_18_44 ? 6'h2c : _T_24856; // @[Mux.scala 31:69:@6016.4]
  assign _T_24858 = valid_18_43 ? 6'h2b : _T_24857; // @[Mux.scala 31:69:@6017.4]
  assign _T_24859 = valid_18_42 ? 6'h2a : _T_24858; // @[Mux.scala 31:69:@6018.4]
  assign _T_24860 = valid_18_41 ? 6'h29 : _T_24859; // @[Mux.scala 31:69:@6019.4]
  assign _T_24861 = valid_18_40 ? 6'h28 : _T_24860; // @[Mux.scala 31:69:@6020.4]
  assign _T_24862 = valid_18_39 ? 6'h27 : _T_24861; // @[Mux.scala 31:69:@6021.4]
  assign _T_24863 = valid_18_38 ? 6'h26 : _T_24862; // @[Mux.scala 31:69:@6022.4]
  assign _T_24864 = valid_18_37 ? 6'h25 : _T_24863; // @[Mux.scala 31:69:@6023.4]
  assign _T_24865 = valid_18_36 ? 6'h24 : _T_24864; // @[Mux.scala 31:69:@6024.4]
  assign _T_24866 = valid_18_35 ? 6'h23 : _T_24865; // @[Mux.scala 31:69:@6025.4]
  assign _T_24867 = valid_18_34 ? 6'h22 : _T_24866; // @[Mux.scala 31:69:@6026.4]
  assign _T_24868 = valid_18_33 ? 6'h21 : _T_24867; // @[Mux.scala 31:69:@6027.4]
  assign _T_24869 = valid_18_32 ? 6'h20 : _T_24868; // @[Mux.scala 31:69:@6028.4]
  assign _T_24870 = valid_18_31 ? 6'h1f : _T_24869; // @[Mux.scala 31:69:@6029.4]
  assign _T_24871 = valid_18_30 ? 6'h1e : _T_24870; // @[Mux.scala 31:69:@6030.4]
  assign _T_24872 = valid_18_29 ? 6'h1d : _T_24871; // @[Mux.scala 31:69:@6031.4]
  assign _T_24873 = valid_18_28 ? 6'h1c : _T_24872; // @[Mux.scala 31:69:@6032.4]
  assign _T_24874 = valid_18_27 ? 6'h1b : _T_24873; // @[Mux.scala 31:69:@6033.4]
  assign _T_24875 = valid_18_26 ? 6'h1a : _T_24874; // @[Mux.scala 31:69:@6034.4]
  assign _T_24876 = valid_18_25 ? 6'h19 : _T_24875; // @[Mux.scala 31:69:@6035.4]
  assign _T_24877 = valid_18_24 ? 6'h18 : _T_24876; // @[Mux.scala 31:69:@6036.4]
  assign _T_24878 = valid_18_23 ? 6'h17 : _T_24877; // @[Mux.scala 31:69:@6037.4]
  assign _T_24879 = valid_18_22 ? 6'h16 : _T_24878; // @[Mux.scala 31:69:@6038.4]
  assign _T_24880 = valid_18_21 ? 6'h15 : _T_24879; // @[Mux.scala 31:69:@6039.4]
  assign _T_24881 = valid_18_20 ? 6'h14 : _T_24880; // @[Mux.scala 31:69:@6040.4]
  assign _T_24882 = valid_18_19 ? 6'h13 : _T_24881; // @[Mux.scala 31:69:@6041.4]
  assign _T_24883 = valid_18_18 ? 6'h12 : _T_24882; // @[Mux.scala 31:69:@6042.4]
  assign _T_24884 = valid_18_17 ? 6'h11 : _T_24883; // @[Mux.scala 31:69:@6043.4]
  assign _T_24885 = valid_18_16 ? 6'h10 : _T_24884; // @[Mux.scala 31:69:@6044.4]
  assign _T_24886 = valid_18_15 ? 6'hf : _T_24885; // @[Mux.scala 31:69:@6045.4]
  assign _T_24887 = valid_18_14 ? 6'he : _T_24886; // @[Mux.scala 31:69:@6046.4]
  assign _T_24888 = valid_18_13 ? 6'hd : _T_24887; // @[Mux.scala 31:69:@6047.4]
  assign _T_24889 = valid_18_12 ? 6'hc : _T_24888; // @[Mux.scala 31:69:@6048.4]
  assign _T_24890 = valid_18_11 ? 6'hb : _T_24889; // @[Mux.scala 31:69:@6049.4]
  assign _T_24891 = valid_18_10 ? 6'ha : _T_24890; // @[Mux.scala 31:69:@6050.4]
  assign _T_24892 = valid_18_9 ? 6'h9 : _T_24891; // @[Mux.scala 31:69:@6051.4]
  assign _T_24893 = valid_18_8 ? 6'h8 : _T_24892; // @[Mux.scala 31:69:@6052.4]
  assign _T_24894 = valid_18_7 ? 6'h7 : _T_24893; // @[Mux.scala 31:69:@6053.4]
  assign _T_24895 = valid_18_6 ? 6'h6 : _T_24894; // @[Mux.scala 31:69:@6054.4]
  assign _T_24896 = valid_18_5 ? 6'h5 : _T_24895; // @[Mux.scala 31:69:@6055.4]
  assign _T_24897 = valid_18_4 ? 6'h4 : _T_24896; // @[Mux.scala 31:69:@6056.4]
  assign _T_24898 = valid_18_3 ? 6'h3 : _T_24897; // @[Mux.scala 31:69:@6057.4]
  assign _T_24899 = valid_18_2 ? 6'h2 : _T_24898; // @[Mux.scala 31:69:@6058.4]
  assign _T_24900 = valid_18_1 ? 6'h1 : _T_24899; // @[Mux.scala 31:69:@6059.4]
  assign select_18 = valid_18_0 ? 6'h0 : _T_24900; // @[Mux.scala 31:69:@6060.4]
  assign _GEN_1153 = 6'h1 == select_18 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1154 = 6'h2 == select_18 ? io_inData_2 : _GEN_1153; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1155 = 6'h3 == select_18 ? io_inData_3 : _GEN_1154; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1156 = 6'h4 == select_18 ? io_inData_4 : _GEN_1155; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1157 = 6'h5 == select_18 ? io_inData_5 : _GEN_1156; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1158 = 6'h6 == select_18 ? io_inData_6 : _GEN_1157; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1159 = 6'h7 == select_18 ? io_inData_7 : _GEN_1158; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1160 = 6'h8 == select_18 ? io_inData_8 : _GEN_1159; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1161 = 6'h9 == select_18 ? io_inData_9 : _GEN_1160; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1162 = 6'ha == select_18 ? io_inData_10 : _GEN_1161; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1163 = 6'hb == select_18 ? io_inData_11 : _GEN_1162; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1164 = 6'hc == select_18 ? io_inData_12 : _GEN_1163; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1165 = 6'hd == select_18 ? io_inData_13 : _GEN_1164; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1166 = 6'he == select_18 ? io_inData_14 : _GEN_1165; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1167 = 6'hf == select_18 ? io_inData_15 : _GEN_1166; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1168 = 6'h10 == select_18 ? io_inData_16 : _GEN_1167; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1169 = 6'h11 == select_18 ? io_inData_17 : _GEN_1168; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1170 = 6'h12 == select_18 ? io_inData_18 : _GEN_1169; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1171 = 6'h13 == select_18 ? io_inData_19 : _GEN_1170; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1172 = 6'h14 == select_18 ? io_inData_20 : _GEN_1171; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1173 = 6'h15 == select_18 ? io_inData_21 : _GEN_1172; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1174 = 6'h16 == select_18 ? io_inData_22 : _GEN_1173; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1175 = 6'h17 == select_18 ? io_inData_23 : _GEN_1174; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1176 = 6'h18 == select_18 ? io_inData_24 : _GEN_1175; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1177 = 6'h19 == select_18 ? io_inData_25 : _GEN_1176; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1178 = 6'h1a == select_18 ? io_inData_26 : _GEN_1177; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1179 = 6'h1b == select_18 ? io_inData_27 : _GEN_1178; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1180 = 6'h1c == select_18 ? io_inData_28 : _GEN_1179; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1181 = 6'h1d == select_18 ? io_inData_29 : _GEN_1180; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1182 = 6'h1e == select_18 ? io_inData_30 : _GEN_1181; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1183 = 6'h1f == select_18 ? io_inData_31 : _GEN_1182; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1184 = 6'h20 == select_18 ? io_inData_32 : _GEN_1183; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1185 = 6'h21 == select_18 ? io_inData_33 : _GEN_1184; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1186 = 6'h22 == select_18 ? io_inData_34 : _GEN_1185; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1187 = 6'h23 == select_18 ? io_inData_35 : _GEN_1186; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1188 = 6'h24 == select_18 ? io_inData_36 : _GEN_1187; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1189 = 6'h25 == select_18 ? io_inData_37 : _GEN_1188; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1190 = 6'h26 == select_18 ? io_inData_38 : _GEN_1189; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1191 = 6'h27 == select_18 ? io_inData_39 : _GEN_1190; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1192 = 6'h28 == select_18 ? io_inData_40 : _GEN_1191; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1193 = 6'h29 == select_18 ? io_inData_41 : _GEN_1192; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1194 = 6'h2a == select_18 ? io_inData_42 : _GEN_1193; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1195 = 6'h2b == select_18 ? io_inData_43 : _GEN_1194; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1196 = 6'h2c == select_18 ? io_inData_44 : _GEN_1195; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1197 = 6'h2d == select_18 ? io_inData_45 : _GEN_1196; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1198 = 6'h2e == select_18 ? io_inData_46 : _GEN_1197; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1199 = 6'h2f == select_18 ? io_inData_47 : _GEN_1198; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1200 = 6'h30 == select_18 ? io_inData_48 : _GEN_1199; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1201 = 6'h31 == select_18 ? io_inData_49 : _GEN_1200; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1202 = 6'h32 == select_18 ? io_inData_50 : _GEN_1201; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1203 = 6'h33 == select_18 ? io_inData_51 : _GEN_1202; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1204 = 6'h34 == select_18 ? io_inData_52 : _GEN_1203; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1205 = 6'h35 == select_18 ? io_inData_53 : _GEN_1204; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1206 = 6'h36 == select_18 ? io_inData_54 : _GEN_1205; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1207 = 6'h37 == select_18 ? io_inData_55 : _GEN_1206; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1208 = 6'h38 == select_18 ? io_inData_56 : _GEN_1207; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1209 = 6'h39 == select_18 ? io_inData_57 : _GEN_1208; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1210 = 6'h3a == select_18 ? io_inData_58 : _GEN_1209; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1211 = 6'h3b == select_18 ? io_inData_59 : _GEN_1210; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1212 = 6'h3c == select_18 ? io_inData_60 : _GEN_1211; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1213 = 6'h3d == select_18 ? io_inData_61 : _GEN_1212; // @[Switch.scala 33:19:@6062.4]
  assign _GEN_1214 = 6'h3e == select_18 ? io_inData_62 : _GEN_1213; // @[Switch.scala 33:19:@6062.4]
  assign _T_24909 = {valid_18_7,valid_18_6,valid_18_5,valid_18_4,valid_18_3,valid_18_2,valid_18_1,valid_18_0}; // @[Switch.scala 34:32:@6069.4]
  assign _T_24917 = {valid_18_15,valid_18_14,valid_18_13,valid_18_12,valid_18_11,valid_18_10,valid_18_9,valid_18_8,_T_24909}; // @[Switch.scala 34:32:@6077.4]
  assign _T_24924 = {valid_18_23,valid_18_22,valid_18_21,valid_18_20,valid_18_19,valid_18_18,valid_18_17,valid_18_16}; // @[Switch.scala 34:32:@6084.4]
  assign _T_24933 = {valid_18_31,valid_18_30,valid_18_29,valid_18_28,valid_18_27,valid_18_26,valid_18_25,valid_18_24,_T_24924,_T_24917}; // @[Switch.scala 34:32:@6093.4]
  assign _T_24940 = {valid_18_39,valid_18_38,valid_18_37,valid_18_36,valid_18_35,valid_18_34,valid_18_33,valid_18_32}; // @[Switch.scala 34:32:@6100.4]
  assign _T_24948 = {valid_18_47,valid_18_46,valid_18_45,valid_18_44,valid_18_43,valid_18_42,valid_18_41,valid_18_40,_T_24940}; // @[Switch.scala 34:32:@6108.4]
  assign _T_24955 = {valid_18_55,valid_18_54,valid_18_53,valid_18_52,valid_18_51,valid_18_50,valid_18_49,valid_18_48}; // @[Switch.scala 34:32:@6115.4]
  assign _T_24964 = {valid_18_63,valid_18_62,valid_18_61,valid_18_60,valid_18_59,valid_18_58,valid_18_57,valid_18_56,_T_24955,_T_24948}; // @[Switch.scala 34:32:@6124.4]
  assign _T_24965 = {_T_24964,_T_24933}; // @[Switch.scala 34:32:@6125.4]
  assign _T_24969 = io_inAddr_0 == 6'h13; // @[Switch.scala 30:53:@6128.4]
  assign valid_19_0 = io_inValid_0 & _T_24969; // @[Switch.scala 30:36:@6129.4]
  assign _T_24972 = io_inAddr_1 == 6'h13; // @[Switch.scala 30:53:@6131.4]
  assign valid_19_1 = io_inValid_1 & _T_24972; // @[Switch.scala 30:36:@6132.4]
  assign _T_24975 = io_inAddr_2 == 6'h13; // @[Switch.scala 30:53:@6134.4]
  assign valid_19_2 = io_inValid_2 & _T_24975; // @[Switch.scala 30:36:@6135.4]
  assign _T_24978 = io_inAddr_3 == 6'h13; // @[Switch.scala 30:53:@6137.4]
  assign valid_19_3 = io_inValid_3 & _T_24978; // @[Switch.scala 30:36:@6138.4]
  assign _T_24981 = io_inAddr_4 == 6'h13; // @[Switch.scala 30:53:@6140.4]
  assign valid_19_4 = io_inValid_4 & _T_24981; // @[Switch.scala 30:36:@6141.4]
  assign _T_24984 = io_inAddr_5 == 6'h13; // @[Switch.scala 30:53:@6143.4]
  assign valid_19_5 = io_inValid_5 & _T_24984; // @[Switch.scala 30:36:@6144.4]
  assign _T_24987 = io_inAddr_6 == 6'h13; // @[Switch.scala 30:53:@6146.4]
  assign valid_19_6 = io_inValid_6 & _T_24987; // @[Switch.scala 30:36:@6147.4]
  assign _T_24990 = io_inAddr_7 == 6'h13; // @[Switch.scala 30:53:@6149.4]
  assign valid_19_7 = io_inValid_7 & _T_24990; // @[Switch.scala 30:36:@6150.4]
  assign _T_24993 = io_inAddr_8 == 6'h13; // @[Switch.scala 30:53:@6152.4]
  assign valid_19_8 = io_inValid_8 & _T_24993; // @[Switch.scala 30:36:@6153.4]
  assign _T_24996 = io_inAddr_9 == 6'h13; // @[Switch.scala 30:53:@6155.4]
  assign valid_19_9 = io_inValid_9 & _T_24996; // @[Switch.scala 30:36:@6156.4]
  assign _T_24999 = io_inAddr_10 == 6'h13; // @[Switch.scala 30:53:@6158.4]
  assign valid_19_10 = io_inValid_10 & _T_24999; // @[Switch.scala 30:36:@6159.4]
  assign _T_25002 = io_inAddr_11 == 6'h13; // @[Switch.scala 30:53:@6161.4]
  assign valid_19_11 = io_inValid_11 & _T_25002; // @[Switch.scala 30:36:@6162.4]
  assign _T_25005 = io_inAddr_12 == 6'h13; // @[Switch.scala 30:53:@6164.4]
  assign valid_19_12 = io_inValid_12 & _T_25005; // @[Switch.scala 30:36:@6165.4]
  assign _T_25008 = io_inAddr_13 == 6'h13; // @[Switch.scala 30:53:@6167.4]
  assign valid_19_13 = io_inValid_13 & _T_25008; // @[Switch.scala 30:36:@6168.4]
  assign _T_25011 = io_inAddr_14 == 6'h13; // @[Switch.scala 30:53:@6170.4]
  assign valid_19_14 = io_inValid_14 & _T_25011; // @[Switch.scala 30:36:@6171.4]
  assign _T_25014 = io_inAddr_15 == 6'h13; // @[Switch.scala 30:53:@6173.4]
  assign valid_19_15 = io_inValid_15 & _T_25014; // @[Switch.scala 30:36:@6174.4]
  assign _T_25017 = io_inAddr_16 == 6'h13; // @[Switch.scala 30:53:@6176.4]
  assign valid_19_16 = io_inValid_16 & _T_25017; // @[Switch.scala 30:36:@6177.4]
  assign _T_25020 = io_inAddr_17 == 6'h13; // @[Switch.scala 30:53:@6179.4]
  assign valid_19_17 = io_inValid_17 & _T_25020; // @[Switch.scala 30:36:@6180.4]
  assign _T_25023 = io_inAddr_18 == 6'h13; // @[Switch.scala 30:53:@6182.4]
  assign valid_19_18 = io_inValid_18 & _T_25023; // @[Switch.scala 30:36:@6183.4]
  assign _T_25026 = io_inAddr_19 == 6'h13; // @[Switch.scala 30:53:@6185.4]
  assign valid_19_19 = io_inValid_19 & _T_25026; // @[Switch.scala 30:36:@6186.4]
  assign _T_25029 = io_inAddr_20 == 6'h13; // @[Switch.scala 30:53:@6188.4]
  assign valid_19_20 = io_inValid_20 & _T_25029; // @[Switch.scala 30:36:@6189.4]
  assign _T_25032 = io_inAddr_21 == 6'h13; // @[Switch.scala 30:53:@6191.4]
  assign valid_19_21 = io_inValid_21 & _T_25032; // @[Switch.scala 30:36:@6192.4]
  assign _T_25035 = io_inAddr_22 == 6'h13; // @[Switch.scala 30:53:@6194.4]
  assign valid_19_22 = io_inValid_22 & _T_25035; // @[Switch.scala 30:36:@6195.4]
  assign _T_25038 = io_inAddr_23 == 6'h13; // @[Switch.scala 30:53:@6197.4]
  assign valid_19_23 = io_inValid_23 & _T_25038; // @[Switch.scala 30:36:@6198.4]
  assign _T_25041 = io_inAddr_24 == 6'h13; // @[Switch.scala 30:53:@6200.4]
  assign valid_19_24 = io_inValid_24 & _T_25041; // @[Switch.scala 30:36:@6201.4]
  assign _T_25044 = io_inAddr_25 == 6'h13; // @[Switch.scala 30:53:@6203.4]
  assign valid_19_25 = io_inValid_25 & _T_25044; // @[Switch.scala 30:36:@6204.4]
  assign _T_25047 = io_inAddr_26 == 6'h13; // @[Switch.scala 30:53:@6206.4]
  assign valid_19_26 = io_inValid_26 & _T_25047; // @[Switch.scala 30:36:@6207.4]
  assign _T_25050 = io_inAddr_27 == 6'h13; // @[Switch.scala 30:53:@6209.4]
  assign valid_19_27 = io_inValid_27 & _T_25050; // @[Switch.scala 30:36:@6210.4]
  assign _T_25053 = io_inAddr_28 == 6'h13; // @[Switch.scala 30:53:@6212.4]
  assign valid_19_28 = io_inValid_28 & _T_25053; // @[Switch.scala 30:36:@6213.4]
  assign _T_25056 = io_inAddr_29 == 6'h13; // @[Switch.scala 30:53:@6215.4]
  assign valid_19_29 = io_inValid_29 & _T_25056; // @[Switch.scala 30:36:@6216.4]
  assign _T_25059 = io_inAddr_30 == 6'h13; // @[Switch.scala 30:53:@6218.4]
  assign valid_19_30 = io_inValid_30 & _T_25059; // @[Switch.scala 30:36:@6219.4]
  assign _T_25062 = io_inAddr_31 == 6'h13; // @[Switch.scala 30:53:@6221.4]
  assign valid_19_31 = io_inValid_31 & _T_25062; // @[Switch.scala 30:36:@6222.4]
  assign _T_25065 = io_inAddr_32 == 6'h13; // @[Switch.scala 30:53:@6224.4]
  assign valid_19_32 = io_inValid_32 & _T_25065; // @[Switch.scala 30:36:@6225.4]
  assign _T_25068 = io_inAddr_33 == 6'h13; // @[Switch.scala 30:53:@6227.4]
  assign valid_19_33 = io_inValid_33 & _T_25068; // @[Switch.scala 30:36:@6228.4]
  assign _T_25071 = io_inAddr_34 == 6'h13; // @[Switch.scala 30:53:@6230.4]
  assign valid_19_34 = io_inValid_34 & _T_25071; // @[Switch.scala 30:36:@6231.4]
  assign _T_25074 = io_inAddr_35 == 6'h13; // @[Switch.scala 30:53:@6233.4]
  assign valid_19_35 = io_inValid_35 & _T_25074; // @[Switch.scala 30:36:@6234.4]
  assign _T_25077 = io_inAddr_36 == 6'h13; // @[Switch.scala 30:53:@6236.4]
  assign valid_19_36 = io_inValid_36 & _T_25077; // @[Switch.scala 30:36:@6237.4]
  assign _T_25080 = io_inAddr_37 == 6'h13; // @[Switch.scala 30:53:@6239.4]
  assign valid_19_37 = io_inValid_37 & _T_25080; // @[Switch.scala 30:36:@6240.4]
  assign _T_25083 = io_inAddr_38 == 6'h13; // @[Switch.scala 30:53:@6242.4]
  assign valid_19_38 = io_inValid_38 & _T_25083; // @[Switch.scala 30:36:@6243.4]
  assign _T_25086 = io_inAddr_39 == 6'h13; // @[Switch.scala 30:53:@6245.4]
  assign valid_19_39 = io_inValid_39 & _T_25086; // @[Switch.scala 30:36:@6246.4]
  assign _T_25089 = io_inAddr_40 == 6'h13; // @[Switch.scala 30:53:@6248.4]
  assign valid_19_40 = io_inValid_40 & _T_25089; // @[Switch.scala 30:36:@6249.4]
  assign _T_25092 = io_inAddr_41 == 6'h13; // @[Switch.scala 30:53:@6251.4]
  assign valid_19_41 = io_inValid_41 & _T_25092; // @[Switch.scala 30:36:@6252.4]
  assign _T_25095 = io_inAddr_42 == 6'h13; // @[Switch.scala 30:53:@6254.4]
  assign valid_19_42 = io_inValid_42 & _T_25095; // @[Switch.scala 30:36:@6255.4]
  assign _T_25098 = io_inAddr_43 == 6'h13; // @[Switch.scala 30:53:@6257.4]
  assign valid_19_43 = io_inValid_43 & _T_25098; // @[Switch.scala 30:36:@6258.4]
  assign _T_25101 = io_inAddr_44 == 6'h13; // @[Switch.scala 30:53:@6260.4]
  assign valid_19_44 = io_inValid_44 & _T_25101; // @[Switch.scala 30:36:@6261.4]
  assign _T_25104 = io_inAddr_45 == 6'h13; // @[Switch.scala 30:53:@6263.4]
  assign valid_19_45 = io_inValid_45 & _T_25104; // @[Switch.scala 30:36:@6264.4]
  assign _T_25107 = io_inAddr_46 == 6'h13; // @[Switch.scala 30:53:@6266.4]
  assign valid_19_46 = io_inValid_46 & _T_25107; // @[Switch.scala 30:36:@6267.4]
  assign _T_25110 = io_inAddr_47 == 6'h13; // @[Switch.scala 30:53:@6269.4]
  assign valid_19_47 = io_inValid_47 & _T_25110; // @[Switch.scala 30:36:@6270.4]
  assign _T_25113 = io_inAddr_48 == 6'h13; // @[Switch.scala 30:53:@6272.4]
  assign valid_19_48 = io_inValid_48 & _T_25113; // @[Switch.scala 30:36:@6273.4]
  assign _T_25116 = io_inAddr_49 == 6'h13; // @[Switch.scala 30:53:@6275.4]
  assign valid_19_49 = io_inValid_49 & _T_25116; // @[Switch.scala 30:36:@6276.4]
  assign _T_25119 = io_inAddr_50 == 6'h13; // @[Switch.scala 30:53:@6278.4]
  assign valid_19_50 = io_inValid_50 & _T_25119; // @[Switch.scala 30:36:@6279.4]
  assign _T_25122 = io_inAddr_51 == 6'h13; // @[Switch.scala 30:53:@6281.4]
  assign valid_19_51 = io_inValid_51 & _T_25122; // @[Switch.scala 30:36:@6282.4]
  assign _T_25125 = io_inAddr_52 == 6'h13; // @[Switch.scala 30:53:@6284.4]
  assign valid_19_52 = io_inValid_52 & _T_25125; // @[Switch.scala 30:36:@6285.4]
  assign _T_25128 = io_inAddr_53 == 6'h13; // @[Switch.scala 30:53:@6287.4]
  assign valid_19_53 = io_inValid_53 & _T_25128; // @[Switch.scala 30:36:@6288.4]
  assign _T_25131 = io_inAddr_54 == 6'h13; // @[Switch.scala 30:53:@6290.4]
  assign valid_19_54 = io_inValid_54 & _T_25131; // @[Switch.scala 30:36:@6291.4]
  assign _T_25134 = io_inAddr_55 == 6'h13; // @[Switch.scala 30:53:@6293.4]
  assign valid_19_55 = io_inValid_55 & _T_25134; // @[Switch.scala 30:36:@6294.4]
  assign _T_25137 = io_inAddr_56 == 6'h13; // @[Switch.scala 30:53:@6296.4]
  assign valid_19_56 = io_inValid_56 & _T_25137; // @[Switch.scala 30:36:@6297.4]
  assign _T_25140 = io_inAddr_57 == 6'h13; // @[Switch.scala 30:53:@6299.4]
  assign valid_19_57 = io_inValid_57 & _T_25140; // @[Switch.scala 30:36:@6300.4]
  assign _T_25143 = io_inAddr_58 == 6'h13; // @[Switch.scala 30:53:@6302.4]
  assign valid_19_58 = io_inValid_58 & _T_25143; // @[Switch.scala 30:36:@6303.4]
  assign _T_25146 = io_inAddr_59 == 6'h13; // @[Switch.scala 30:53:@6305.4]
  assign valid_19_59 = io_inValid_59 & _T_25146; // @[Switch.scala 30:36:@6306.4]
  assign _T_25149 = io_inAddr_60 == 6'h13; // @[Switch.scala 30:53:@6308.4]
  assign valid_19_60 = io_inValid_60 & _T_25149; // @[Switch.scala 30:36:@6309.4]
  assign _T_25152 = io_inAddr_61 == 6'h13; // @[Switch.scala 30:53:@6311.4]
  assign valid_19_61 = io_inValid_61 & _T_25152; // @[Switch.scala 30:36:@6312.4]
  assign _T_25155 = io_inAddr_62 == 6'h13; // @[Switch.scala 30:53:@6314.4]
  assign valid_19_62 = io_inValid_62 & _T_25155; // @[Switch.scala 30:36:@6315.4]
  assign _T_25158 = io_inAddr_63 == 6'h13; // @[Switch.scala 30:53:@6317.4]
  assign valid_19_63 = io_inValid_63 & _T_25158; // @[Switch.scala 30:36:@6318.4]
  assign _T_25224 = valid_19_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@6320.4]
  assign _T_25225 = valid_19_61 ? 6'h3d : _T_25224; // @[Mux.scala 31:69:@6321.4]
  assign _T_25226 = valid_19_60 ? 6'h3c : _T_25225; // @[Mux.scala 31:69:@6322.4]
  assign _T_25227 = valid_19_59 ? 6'h3b : _T_25226; // @[Mux.scala 31:69:@6323.4]
  assign _T_25228 = valid_19_58 ? 6'h3a : _T_25227; // @[Mux.scala 31:69:@6324.4]
  assign _T_25229 = valid_19_57 ? 6'h39 : _T_25228; // @[Mux.scala 31:69:@6325.4]
  assign _T_25230 = valid_19_56 ? 6'h38 : _T_25229; // @[Mux.scala 31:69:@6326.4]
  assign _T_25231 = valid_19_55 ? 6'h37 : _T_25230; // @[Mux.scala 31:69:@6327.4]
  assign _T_25232 = valid_19_54 ? 6'h36 : _T_25231; // @[Mux.scala 31:69:@6328.4]
  assign _T_25233 = valid_19_53 ? 6'h35 : _T_25232; // @[Mux.scala 31:69:@6329.4]
  assign _T_25234 = valid_19_52 ? 6'h34 : _T_25233; // @[Mux.scala 31:69:@6330.4]
  assign _T_25235 = valid_19_51 ? 6'h33 : _T_25234; // @[Mux.scala 31:69:@6331.4]
  assign _T_25236 = valid_19_50 ? 6'h32 : _T_25235; // @[Mux.scala 31:69:@6332.4]
  assign _T_25237 = valid_19_49 ? 6'h31 : _T_25236; // @[Mux.scala 31:69:@6333.4]
  assign _T_25238 = valid_19_48 ? 6'h30 : _T_25237; // @[Mux.scala 31:69:@6334.4]
  assign _T_25239 = valid_19_47 ? 6'h2f : _T_25238; // @[Mux.scala 31:69:@6335.4]
  assign _T_25240 = valid_19_46 ? 6'h2e : _T_25239; // @[Mux.scala 31:69:@6336.4]
  assign _T_25241 = valid_19_45 ? 6'h2d : _T_25240; // @[Mux.scala 31:69:@6337.4]
  assign _T_25242 = valid_19_44 ? 6'h2c : _T_25241; // @[Mux.scala 31:69:@6338.4]
  assign _T_25243 = valid_19_43 ? 6'h2b : _T_25242; // @[Mux.scala 31:69:@6339.4]
  assign _T_25244 = valid_19_42 ? 6'h2a : _T_25243; // @[Mux.scala 31:69:@6340.4]
  assign _T_25245 = valid_19_41 ? 6'h29 : _T_25244; // @[Mux.scala 31:69:@6341.4]
  assign _T_25246 = valid_19_40 ? 6'h28 : _T_25245; // @[Mux.scala 31:69:@6342.4]
  assign _T_25247 = valid_19_39 ? 6'h27 : _T_25246; // @[Mux.scala 31:69:@6343.4]
  assign _T_25248 = valid_19_38 ? 6'h26 : _T_25247; // @[Mux.scala 31:69:@6344.4]
  assign _T_25249 = valid_19_37 ? 6'h25 : _T_25248; // @[Mux.scala 31:69:@6345.4]
  assign _T_25250 = valid_19_36 ? 6'h24 : _T_25249; // @[Mux.scala 31:69:@6346.4]
  assign _T_25251 = valid_19_35 ? 6'h23 : _T_25250; // @[Mux.scala 31:69:@6347.4]
  assign _T_25252 = valid_19_34 ? 6'h22 : _T_25251; // @[Mux.scala 31:69:@6348.4]
  assign _T_25253 = valid_19_33 ? 6'h21 : _T_25252; // @[Mux.scala 31:69:@6349.4]
  assign _T_25254 = valid_19_32 ? 6'h20 : _T_25253; // @[Mux.scala 31:69:@6350.4]
  assign _T_25255 = valid_19_31 ? 6'h1f : _T_25254; // @[Mux.scala 31:69:@6351.4]
  assign _T_25256 = valid_19_30 ? 6'h1e : _T_25255; // @[Mux.scala 31:69:@6352.4]
  assign _T_25257 = valid_19_29 ? 6'h1d : _T_25256; // @[Mux.scala 31:69:@6353.4]
  assign _T_25258 = valid_19_28 ? 6'h1c : _T_25257; // @[Mux.scala 31:69:@6354.4]
  assign _T_25259 = valid_19_27 ? 6'h1b : _T_25258; // @[Mux.scala 31:69:@6355.4]
  assign _T_25260 = valid_19_26 ? 6'h1a : _T_25259; // @[Mux.scala 31:69:@6356.4]
  assign _T_25261 = valid_19_25 ? 6'h19 : _T_25260; // @[Mux.scala 31:69:@6357.4]
  assign _T_25262 = valid_19_24 ? 6'h18 : _T_25261; // @[Mux.scala 31:69:@6358.4]
  assign _T_25263 = valid_19_23 ? 6'h17 : _T_25262; // @[Mux.scala 31:69:@6359.4]
  assign _T_25264 = valid_19_22 ? 6'h16 : _T_25263; // @[Mux.scala 31:69:@6360.4]
  assign _T_25265 = valid_19_21 ? 6'h15 : _T_25264; // @[Mux.scala 31:69:@6361.4]
  assign _T_25266 = valid_19_20 ? 6'h14 : _T_25265; // @[Mux.scala 31:69:@6362.4]
  assign _T_25267 = valid_19_19 ? 6'h13 : _T_25266; // @[Mux.scala 31:69:@6363.4]
  assign _T_25268 = valid_19_18 ? 6'h12 : _T_25267; // @[Mux.scala 31:69:@6364.4]
  assign _T_25269 = valid_19_17 ? 6'h11 : _T_25268; // @[Mux.scala 31:69:@6365.4]
  assign _T_25270 = valid_19_16 ? 6'h10 : _T_25269; // @[Mux.scala 31:69:@6366.4]
  assign _T_25271 = valid_19_15 ? 6'hf : _T_25270; // @[Mux.scala 31:69:@6367.4]
  assign _T_25272 = valid_19_14 ? 6'he : _T_25271; // @[Mux.scala 31:69:@6368.4]
  assign _T_25273 = valid_19_13 ? 6'hd : _T_25272; // @[Mux.scala 31:69:@6369.4]
  assign _T_25274 = valid_19_12 ? 6'hc : _T_25273; // @[Mux.scala 31:69:@6370.4]
  assign _T_25275 = valid_19_11 ? 6'hb : _T_25274; // @[Mux.scala 31:69:@6371.4]
  assign _T_25276 = valid_19_10 ? 6'ha : _T_25275; // @[Mux.scala 31:69:@6372.4]
  assign _T_25277 = valid_19_9 ? 6'h9 : _T_25276; // @[Mux.scala 31:69:@6373.4]
  assign _T_25278 = valid_19_8 ? 6'h8 : _T_25277; // @[Mux.scala 31:69:@6374.4]
  assign _T_25279 = valid_19_7 ? 6'h7 : _T_25278; // @[Mux.scala 31:69:@6375.4]
  assign _T_25280 = valid_19_6 ? 6'h6 : _T_25279; // @[Mux.scala 31:69:@6376.4]
  assign _T_25281 = valid_19_5 ? 6'h5 : _T_25280; // @[Mux.scala 31:69:@6377.4]
  assign _T_25282 = valid_19_4 ? 6'h4 : _T_25281; // @[Mux.scala 31:69:@6378.4]
  assign _T_25283 = valid_19_3 ? 6'h3 : _T_25282; // @[Mux.scala 31:69:@6379.4]
  assign _T_25284 = valid_19_2 ? 6'h2 : _T_25283; // @[Mux.scala 31:69:@6380.4]
  assign _T_25285 = valid_19_1 ? 6'h1 : _T_25284; // @[Mux.scala 31:69:@6381.4]
  assign select_19 = valid_19_0 ? 6'h0 : _T_25285; // @[Mux.scala 31:69:@6382.4]
  assign _GEN_1217 = 6'h1 == select_19 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1218 = 6'h2 == select_19 ? io_inData_2 : _GEN_1217; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1219 = 6'h3 == select_19 ? io_inData_3 : _GEN_1218; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1220 = 6'h4 == select_19 ? io_inData_4 : _GEN_1219; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1221 = 6'h5 == select_19 ? io_inData_5 : _GEN_1220; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1222 = 6'h6 == select_19 ? io_inData_6 : _GEN_1221; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1223 = 6'h7 == select_19 ? io_inData_7 : _GEN_1222; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1224 = 6'h8 == select_19 ? io_inData_8 : _GEN_1223; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1225 = 6'h9 == select_19 ? io_inData_9 : _GEN_1224; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1226 = 6'ha == select_19 ? io_inData_10 : _GEN_1225; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1227 = 6'hb == select_19 ? io_inData_11 : _GEN_1226; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1228 = 6'hc == select_19 ? io_inData_12 : _GEN_1227; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1229 = 6'hd == select_19 ? io_inData_13 : _GEN_1228; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1230 = 6'he == select_19 ? io_inData_14 : _GEN_1229; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1231 = 6'hf == select_19 ? io_inData_15 : _GEN_1230; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1232 = 6'h10 == select_19 ? io_inData_16 : _GEN_1231; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1233 = 6'h11 == select_19 ? io_inData_17 : _GEN_1232; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1234 = 6'h12 == select_19 ? io_inData_18 : _GEN_1233; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1235 = 6'h13 == select_19 ? io_inData_19 : _GEN_1234; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1236 = 6'h14 == select_19 ? io_inData_20 : _GEN_1235; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1237 = 6'h15 == select_19 ? io_inData_21 : _GEN_1236; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1238 = 6'h16 == select_19 ? io_inData_22 : _GEN_1237; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1239 = 6'h17 == select_19 ? io_inData_23 : _GEN_1238; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1240 = 6'h18 == select_19 ? io_inData_24 : _GEN_1239; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1241 = 6'h19 == select_19 ? io_inData_25 : _GEN_1240; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1242 = 6'h1a == select_19 ? io_inData_26 : _GEN_1241; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1243 = 6'h1b == select_19 ? io_inData_27 : _GEN_1242; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1244 = 6'h1c == select_19 ? io_inData_28 : _GEN_1243; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1245 = 6'h1d == select_19 ? io_inData_29 : _GEN_1244; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1246 = 6'h1e == select_19 ? io_inData_30 : _GEN_1245; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1247 = 6'h1f == select_19 ? io_inData_31 : _GEN_1246; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1248 = 6'h20 == select_19 ? io_inData_32 : _GEN_1247; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1249 = 6'h21 == select_19 ? io_inData_33 : _GEN_1248; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1250 = 6'h22 == select_19 ? io_inData_34 : _GEN_1249; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1251 = 6'h23 == select_19 ? io_inData_35 : _GEN_1250; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1252 = 6'h24 == select_19 ? io_inData_36 : _GEN_1251; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1253 = 6'h25 == select_19 ? io_inData_37 : _GEN_1252; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1254 = 6'h26 == select_19 ? io_inData_38 : _GEN_1253; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1255 = 6'h27 == select_19 ? io_inData_39 : _GEN_1254; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1256 = 6'h28 == select_19 ? io_inData_40 : _GEN_1255; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1257 = 6'h29 == select_19 ? io_inData_41 : _GEN_1256; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1258 = 6'h2a == select_19 ? io_inData_42 : _GEN_1257; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1259 = 6'h2b == select_19 ? io_inData_43 : _GEN_1258; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1260 = 6'h2c == select_19 ? io_inData_44 : _GEN_1259; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1261 = 6'h2d == select_19 ? io_inData_45 : _GEN_1260; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1262 = 6'h2e == select_19 ? io_inData_46 : _GEN_1261; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1263 = 6'h2f == select_19 ? io_inData_47 : _GEN_1262; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1264 = 6'h30 == select_19 ? io_inData_48 : _GEN_1263; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1265 = 6'h31 == select_19 ? io_inData_49 : _GEN_1264; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1266 = 6'h32 == select_19 ? io_inData_50 : _GEN_1265; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1267 = 6'h33 == select_19 ? io_inData_51 : _GEN_1266; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1268 = 6'h34 == select_19 ? io_inData_52 : _GEN_1267; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1269 = 6'h35 == select_19 ? io_inData_53 : _GEN_1268; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1270 = 6'h36 == select_19 ? io_inData_54 : _GEN_1269; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1271 = 6'h37 == select_19 ? io_inData_55 : _GEN_1270; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1272 = 6'h38 == select_19 ? io_inData_56 : _GEN_1271; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1273 = 6'h39 == select_19 ? io_inData_57 : _GEN_1272; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1274 = 6'h3a == select_19 ? io_inData_58 : _GEN_1273; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1275 = 6'h3b == select_19 ? io_inData_59 : _GEN_1274; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1276 = 6'h3c == select_19 ? io_inData_60 : _GEN_1275; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1277 = 6'h3d == select_19 ? io_inData_61 : _GEN_1276; // @[Switch.scala 33:19:@6384.4]
  assign _GEN_1278 = 6'h3e == select_19 ? io_inData_62 : _GEN_1277; // @[Switch.scala 33:19:@6384.4]
  assign _T_25294 = {valid_19_7,valid_19_6,valid_19_5,valid_19_4,valid_19_3,valid_19_2,valid_19_1,valid_19_0}; // @[Switch.scala 34:32:@6391.4]
  assign _T_25302 = {valid_19_15,valid_19_14,valid_19_13,valid_19_12,valid_19_11,valid_19_10,valid_19_9,valid_19_8,_T_25294}; // @[Switch.scala 34:32:@6399.4]
  assign _T_25309 = {valid_19_23,valid_19_22,valid_19_21,valid_19_20,valid_19_19,valid_19_18,valid_19_17,valid_19_16}; // @[Switch.scala 34:32:@6406.4]
  assign _T_25318 = {valid_19_31,valid_19_30,valid_19_29,valid_19_28,valid_19_27,valid_19_26,valid_19_25,valid_19_24,_T_25309,_T_25302}; // @[Switch.scala 34:32:@6415.4]
  assign _T_25325 = {valid_19_39,valid_19_38,valid_19_37,valid_19_36,valid_19_35,valid_19_34,valid_19_33,valid_19_32}; // @[Switch.scala 34:32:@6422.4]
  assign _T_25333 = {valid_19_47,valid_19_46,valid_19_45,valid_19_44,valid_19_43,valid_19_42,valid_19_41,valid_19_40,_T_25325}; // @[Switch.scala 34:32:@6430.4]
  assign _T_25340 = {valid_19_55,valid_19_54,valid_19_53,valid_19_52,valid_19_51,valid_19_50,valid_19_49,valid_19_48}; // @[Switch.scala 34:32:@6437.4]
  assign _T_25349 = {valid_19_63,valid_19_62,valid_19_61,valid_19_60,valid_19_59,valid_19_58,valid_19_57,valid_19_56,_T_25340,_T_25333}; // @[Switch.scala 34:32:@6446.4]
  assign _T_25350 = {_T_25349,_T_25318}; // @[Switch.scala 34:32:@6447.4]
  assign _T_25354 = io_inAddr_0 == 6'h14; // @[Switch.scala 30:53:@6450.4]
  assign valid_20_0 = io_inValid_0 & _T_25354; // @[Switch.scala 30:36:@6451.4]
  assign _T_25357 = io_inAddr_1 == 6'h14; // @[Switch.scala 30:53:@6453.4]
  assign valid_20_1 = io_inValid_1 & _T_25357; // @[Switch.scala 30:36:@6454.4]
  assign _T_25360 = io_inAddr_2 == 6'h14; // @[Switch.scala 30:53:@6456.4]
  assign valid_20_2 = io_inValid_2 & _T_25360; // @[Switch.scala 30:36:@6457.4]
  assign _T_25363 = io_inAddr_3 == 6'h14; // @[Switch.scala 30:53:@6459.4]
  assign valid_20_3 = io_inValid_3 & _T_25363; // @[Switch.scala 30:36:@6460.4]
  assign _T_25366 = io_inAddr_4 == 6'h14; // @[Switch.scala 30:53:@6462.4]
  assign valid_20_4 = io_inValid_4 & _T_25366; // @[Switch.scala 30:36:@6463.4]
  assign _T_25369 = io_inAddr_5 == 6'h14; // @[Switch.scala 30:53:@6465.4]
  assign valid_20_5 = io_inValid_5 & _T_25369; // @[Switch.scala 30:36:@6466.4]
  assign _T_25372 = io_inAddr_6 == 6'h14; // @[Switch.scala 30:53:@6468.4]
  assign valid_20_6 = io_inValid_6 & _T_25372; // @[Switch.scala 30:36:@6469.4]
  assign _T_25375 = io_inAddr_7 == 6'h14; // @[Switch.scala 30:53:@6471.4]
  assign valid_20_7 = io_inValid_7 & _T_25375; // @[Switch.scala 30:36:@6472.4]
  assign _T_25378 = io_inAddr_8 == 6'h14; // @[Switch.scala 30:53:@6474.4]
  assign valid_20_8 = io_inValid_8 & _T_25378; // @[Switch.scala 30:36:@6475.4]
  assign _T_25381 = io_inAddr_9 == 6'h14; // @[Switch.scala 30:53:@6477.4]
  assign valid_20_9 = io_inValid_9 & _T_25381; // @[Switch.scala 30:36:@6478.4]
  assign _T_25384 = io_inAddr_10 == 6'h14; // @[Switch.scala 30:53:@6480.4]
  assign valid_20_10 = io_inValid_10 & _T_25384; // @[Switch.scala 30:36:@6481.4]
  assign _T_25387 = io_inAddr_11 == 6'h14; // @[Switch.scala 30:53:@6483.4]
  assign valid_20_11 = io_inValid_11 & _T_25387; // @[Switch.scala 30:36:@6484.4]
  assign _T_25390 = io_inAddr_12 == 6'h14; // @[Switch.scala 30:53:@6486.4]
  assign valid_20_12 = io_inValid_12 & _T_25390; // @[Switch.scala 30:36:@6487.4]
  assign _T_25393 = io_inAddr_13 == 6'h14; // @[Switch.scala 30:53:@6489.4]
  assign valid_20_13 = io_inValid_13 & _T_25393; // @[Switch.scala 30:36:@6490.4]
  assign _T_25396 = io_inAddr_14 == 6'h14; // @[Switch.scala 30:53:@6492.4]
  assign valid_20_14 = io_inValid_14 & _T_25396; // @[Switch.scala 30:36:@6493.4]
  assign _T_25399 = io_inAddr_15 == 6'h14; // @[Switch.scala 30:53:@6495.4]
  assign valid_20_15 = io_inValid_15 & _T_25399; // @[Switch.scala 30:36:@6496.4]
  assign _T_25402 = io_inAddr_16 == 6'h14; // @[Switch.scala 30:53:@6498.4]
  assign valid_20_16 = io_inValid_16 & _T_25402; // @[Switch.scala 30:36:@6499.4]
  assign _T_25405 = io_inAddr_17 == 6'h14; // @[Switch.scala 30:53:@6501.4]
  assign valid_20_17 = io_inValid_17 & _T_25405; // @[Switch.scala 30:36:@6502.4]
  assign _T_25408 = io_inAddr_18 == 6'h14; // @[Switch.scala 30:53:@6504.4]
  assign valid_20_18 = io_inValid_18 & _T_25408; // @[Switch.scala 30:36:@6505.4]
  assign _T_25411 = io_inAddr_19 == 6'h14; // @[Switch.scala 30:53:@6507.4]
  assign valid_20_19 = io_inValid_19 & _T_25411; // @[Switch.scala 30:36:@6508.4]
  assign _T_25414 = io_inAddr_20 == 6'h14; // @[Switch.scala 30:53:@6510.4]
  assign valid_20_20 = io_inValid_20 & _T_25414; // @[Switch.scala 30:36:@6511.4]
  assign _T_25417 = io_inAddr_21 == 6'h14; // @[Switch.scala 30:53:@6513.4]
  assign valid_20_21 = io_inValid_21 & _T_25417; // @[Switch.scala 30:36:@6514.4]
  assign _T_25420 = io_inAddr_22 == 6'h14; // @[Switch.scala 30:53:@6516.4]
  assign valid_20_22 = io_inValid_22 & _T_25420; // @[Switch.scala 30:36:@6517.4]
  assign _T_25423 = io_inAddr_23 == 6'h14; // @[Switch.scala 30:53:@6519.4]
  assign valid_20_23 = io_inValid_23 & _T_25423; // @[Switch.scala 30:36:@6520.4]
  assign _T_25426 = io_inAddr_24 == 6'h14; // @[Switch.scala 30:53:@6522.4]
  assign valid_20_24 = io_inValid_24 & _T_25426; // @[Switch.scala 30:36:@6523.4]
  assign _T_25429 = io_inAddr_25 == 6'h14; // @[Switch.scala 30:53:@6525.4]
  assign valid_20_25 = io_inValid_25 & _T_25429; // @[Switch.scala 30:36:@6526.4]
  assign _T_25432 = io_inAddr_26 == 6'h14; // @[Switch.scala 30:53:@6528.4]
  assign valid_20_26 = io_inValid_26 & _T_25432; // @[Switch.scala 30:36:@6529.4]
  assign _T_25435 = io_inAddr_27 == 6'h14; // @[Switch.scala 30:53:@6531.4]
  assign valid_20_27 = io_inValid_27 & _T_25435; // @[Switch.scala 30:36:@6532.4]
  assign _T_25438 = io_inAddr_28 == 6'h14; // @[Switch.scala 30:53:@6534.4]
  assign valid_20_28 = io_inValid_28 & _T_25438; // @[Switch.scala 30:36:@6535.4]
  assign _T_25441 = io_inAddr_29 == 6'h14; // @[Switch.scala 30:53:@6537.4]
  assign valid_20_29 = io_inValid_29 & _T_25441; // @[Switch.scala 30:36:@6538.4]
  assign _T_25444 = io_inAddr_30 == 6'h14; // @[Switch.scala 30:53:@6540.4]
  assign valid_20_30 = io_inValid_30 & _T_25444; // @[Switch.scala 30:36:@6541.4]
  assign _T_25447 = io_inAddr_31 == 6'h14; // @[Switch.scala 30:53:@6543.4]
  assign valid_20_31 = io_inValid_31 & _T_25447; // @[Switch.scala 30:36:@6544.4]
  assign _T_25450 = io_inAddr_32 == 6'h14; // @[Switch.scala 30:53:@6546.4]
  assign valid_20_32 = io_inValid_32 & _T_25450; // @[Switch.scala 30:36:@6547.4]
  assign _T_25453 = io_inAddr_33 == 6'h14; // @[Switch.scala 30:53:@6549.4]
  assign valid_20_33 = io_inValid_33 & _T_25453; // @[Switch.scala 30:36:@6550.4]
  assign _T_25456 = io_inAddr_34 == 6'h14; // @[Switch.scala 30:53:@6552.4]
  assign valid_20_34 = io_inValid_34 & _T_25456; // @[Switch.scala 30:36:@6553.4]
  assign _T_25459 = io_inAddr_35 == 6'h14; // @[Switch.scala 30:53:@6555.4]
  assign valid_20_35 = io_inValid_35 & _T_25459; // @[Switch.scala 30:36:@6556.4]
  assign _T_25462 = io_inAddr_36 == 6'h14; // @[Switch.scala 30:53:@6558.4]
  assign valid_20_36 = io_inValid_36 & _T_25462; // @[Switch.scala 30:36:@6559.4]
  assign _T_25465 = io_inAddr_37 == 6'h14; // @[Switch.scala 30:53:@6561.4]
  assign valid_20_37 = io_inValid_37 & _T_25465; // @[Switch.scala 30:36:@6562.4]
  assign _T_25468 = io_inAddr_38 == 6'h14; // @[Switch.scala 30:53:@6564.4]
  assign valid_20_38 = io_inValid_38 & _T_25468; // @[Switch.scala 30:36:@6565.4]
  assign _T_25471 = io_inAddr_39 == 6'h14; // @[Switch.scala 30:53:@6567.4]
  assign valid_20_39 = io_inValid_39 & _T_25471; // @[Switch.scala 30:36:@6568.4]
  assign _T_25474 = io_inAddr_40 == 6'h14; // @[Switch.scala 30:53:@6570.4]
  assign valid_20_40 = io_inValid_40 & _T_25474; // @[Switch.scala 30:36:@6571.4]
  assign _T_25477 = io_inAddr_41 == 6'h14; // @[Switch.scala 30:53:@6573.4]
  assign valid_20_41 = io_inValid_41 & _T_25477; // @[Switch.scala 30:36:@6574.4]
  assign _T_25480 = io_inAddr_42 == 6'h14; // @[Switch.scala 30:53:@6576.4]
  assign valid_20_42 = io_inValid_42 & _T_25480; // @[Switch.scala 30:36:@6577.4]
  assign _T_25483 = io_inAddr_43 == 6'h14; // @[Switch.scala 30:53:@6579.4]
  assign valid_20_43 = io_inValid_43 & _T_25483; // @[Switch.scala 30:36:@6580.4]
  assign _T_25486 = io_inAddr_44 == 6'h14; // @[Switch.scala 30:53:@6582.4]
  assign valid_20_44 = io_inValid_44 & _T_25486; // @[Switch.scala 30:36:@6583.4]
  assign _T_25489 = io_inAddr_45 == 6'h14; // @[Switch.scala 30:53:@6585.4]
  assign valid_20_45 = io_inValid_45 & _T_25489; // @[Switch.scala 30:36:@6586.4]
  assign _T_25492 = io_inAddr_46 == 6'h14; // @[Switch.scala 30:53:@6588.4]
  assign valid_20_46 = io_inValid_46 & _T_25492; // @[Switch.scala 30:36:@6589.4]
  assign _T_25495 = io_inAddr_47 == 6'h14; // @[Switch.scala 30:53:@6591.4]
  assign valid_20_47 = io_inValid_47 & _T_25495; // @[Switch.scala 30:36:@6592.4]
  assign _T_25498 = io_inAddr_48 == 6'h14; // @[Switch.scala 30:53:@6594.4]
  assign valid_20_48 = io_inValid_48 & _T_25498; // @[Switch.scala 30:36:@6595.4]
  assign _T_25501 = io_inAddr_49 == 6'h14; // @[Switch.scala 30:53:@6597.4]
  assign valid_20_49 = io_inValid_49 & _T_25501; // @[Switch.scala 30:36:@6598.4]
  assign _T_25504 = io_inAddr_50 == 6'h14; // @[Switch.scala 30:53:@6600.4]
  assign valid_20_50 = io_inValid_50 & _T_25504; // @[Switch.scala 30:36:@6601.4]
  assign _T_25507 = io_inAddr_51 == 6'h14; // @[Switch.scala 30:53:@6603.4]
  assign valid_20_51 = io_inValid_51 & _T_25507; // @[Switch.scala 30:36:@6604.4]
  assign _T_25510 = io_inAddr_52 == 6'h14; // @[Switch.scala 30:53:@6606.4]
  assign valid_20_52 = io_inValid_52 & _T_25510; // @[Switch.scala 30:36:@6607.4]
  assign _T_25513 = io_inAddr_53 == 6'h14; // @[Switch.scala 30:53:@6609.4]
  assign valid_20_53 = io_inValid_53 & _T_25513; // @[Switch.scala 30:36:@6610.4]
  assign _T_25516 = io_inAddr_54 == 6'h14; // @[Switch.scala 30:53:@6612.4]
  assign valid_20_54 = io_inValid_54 & _T_25516; // @[Switch.scala 30:36:@6613.4]
  assign _T_25519 = io_inAddr_55 == 6'h14; // @[Switch.scala 30:53:@6615.4]
  assign valid_20_55 = io_inValid_55 & _T_25519; // @[Switch.scala 30:36:@6616.4]
  assign _T_25522 = io_inAddr_56 == 6'h14; // @[Switch.scala 30:53:@6618.4]
  assign valid_20_56 = io_inValid_56 & _T_25522; // @[Switch.scala 30:36:@6619.4]
  assign _T_25525 = io_inAddr_57 == 6'h14; // @[Switch.scala 30:53:@6621.4]
  assign valid_20_57 = io_inValid_57 & _T_25525; // @[Switch.scala 30:36:@6622.4]
  assign _T_25528 = io_inAddr_58 == 6'h14; // @[Switch.scala 30:53:@6624.4]
  assign valid_20_58 = io_inValid_58 & _T_25528; // @[Switch.scala 30:36:@6625.4]
  assign _T_25531 = io_inAddr_59 == 6'h14; // @[Switch.scala 30:53:@6627.4]
  assign valid_20_59 = io_inValid_59 & _T_25531; // @[Switch.scala 30:36:@6628.4]
  assign _T_25534 = io_inAddr_60 == 6'h14; // @[Switch.scala 30:53:@6630.4]
  assign valid_20_60 = io_inValid_60 & _T_25534; // @[Switch.scala 30:36:@6631.4]
  assign _T_25537 = io_inAddr_61 == 6'h14; // @[Switch.scala 30:53:@6633.4]
  assign valid_20_61 = io_inValid_61 & _T_25537; // @[Switch.scala 30:36:@6634.4]
  assign _T_25540 = io_inAddr_62 == 6'h14; // @[Switch.scala 30:53:@6636.4]
  assign valid_20_62 = io_inValid_62 & _T_25540; // @[Switch.scala 30:36:@6637.4]
  assign _T_25543 = io_inAddr_63 == 6'h14; // @[Switch.scala 30:53:@6639.4]
  assign valid_20_63 = io_inValid_63 & _T_25543; // @[Switch.scala 30:36:@6640.4]
  assign _T_25609 = valid_20_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@6642.4]
  assign _T_25610 = valid_20_61 ? 6'h3d : _T_25609; // @[Mux.scala 31:69:@6643.4]
  assign _T_25611 = valid_20_60 ? 6'h3c : _T_25610; // @[Mux.scala 31:69:@6644.4]
  assign _T_25612 = valid_20_59 ? 6'h3b : _T_25611; // @[Mux.scala 31:69:@6645.4]
  assign _T_25613 = valid_20_58 ? 6'h3a : _T_25612; // @[Mux.scala 31:69:@6646.4]
  assign _T_25614 = valid_20_57 ? 6'h39 : _T_25613; // @[Mux.scala 31:69:@6647.4]
  assign _T_25615 = valid_20_56 ? 6'h38 : _T_25614; // @[Mux.scala 31:69:@6648.4]
  assign _T_25616 = valid_20_55 ? 6'h37 : _T_25615; // @[Mux.scala 31:69:@6649.4]
  assign _T_25617 = valid_20_54 ? 6'h36 : _T_25616; // @[Mux.scala 31:69:@6650.4]
  assign _T_25618 = valid_20_53 ? 6'h35 : _T_25617; // @[Mux.scala 31:69:@6651.4]
  assign _T_25619 = valid_20_52 ? 6'h34 : _T_25618; // @[Mux.scala 31:69:@6652.4]
  assign _T_25620 = valid_20_51 ? 6'h33 : _T_25619; // @[Mux.scala 31:69:@6653.4]
  assign _T_25621 = valid_20_50 ? 6'h32 : _T_25620; // @[Mux.scala 31:69:@6654.4]
  assign _T_25622 = valid_20_49 ? 6'h31 : _T_25621; // @[Mux.scala 31:69:@6655.4]
  assign _T_25623 = valid_20_48 ? 6'h30 : _T_25622; // @[Mux.scala 31:69:@6656.4]
  assign _T_25624 = valid_20_47 ? 6'h2f : _T_25623; // @[Mux.scala 31:69:@6657.4]
  assign _T_25625 = valid_20_46 ? 6'h2e : _T_25624; // @[Mux.scala 31:69:@6658.4]
  assign _T_25626 = valid_20_45 ? 6'h2d : _T_25625; // @[Mux.scala 31:69:@6659.4]
  assign _T_25627 = valid_20_44 ? 6'h2c : _T_25626; // @[Mux.scala 31:69:@6660.4]
  assign _T_25628 = valid_20_43 ? 6'h2b : _T_25627; // @[Mux.scala 31:69:@6661.4]
  assign _T_25629 = valid_20_42 ? 6'h2a : _T_25628; // @[Mux.scala 31:69:@6662.4]
  assign _T_25630 = valid_20_41 ? 6'h29 : _T_25629; // @[Mux.scala 31:69:@6663.4]
  assign _T_25631 = valid_20_40 ? 6'h28 : _T_25630; // @[Mux.scala 31:69:@6664.4]
  assign _T_25632 = valid_20_39 ? 6'h27 : _T_25631; // @[Mux.scala 31:69:@6665.4]
  assign _T_25633 = valid_20_38 ? 6'h26 : _T_25632; // @[Mux.scala 31:69:@6666.4]
  assign _T_25634 = valid_20_37 ? 6'h25 : _T_25633; // @[Mux.scala 31:69:@6667.4]
  assign _T_25635 = valid_20_36 ? 6'h24 : _T_25634; // @[Mux.scala 31:69:@6668.4]
  assign _T_25636 = valid_20_35 ? 6'h23 : _T_25635; // @[Mux.scala 31:69:@6669.4]
  assign _T_25637 = valid_20_34 ? 6'h22 : _T_25636; // @[Mux.scala 31:69:@6670.4]
  assign _T_25638 = valid_20_33 ? 6'h21 : _T_25637; // @[Mux.scala 31:69:@6671.4]
  assign _T_25639 = valid_20_32 ? 6'h20 : _T_25638; // @[Mux.scala 31:69:@6672.4]
  assign _T_25640 = valid_20_31 ? 6'h1f : _T_25639; // @[Mux.scala 31:69:@6673.4]
  assign _T_25641 = valid_20_30 ? 6'h1e : _T_25640; // @[Mux.scala 31:69:@6674.4]
  assign _T_25642 = valid_20_29 ? 6'h1d : _T_25641; // @[Mux.scala 31:69:@6675.4]
  assign _T_25643 = valid_20_28 ? 6'h1c : _T_25642; // @[Mux.scala 31:69:@6676.4]
  assign _T_25644 = valid_20_27 ? 6'h1b : _T_25643; // @[Mux.scala 31:69:@6677.4]
  assign _T_25645 = valid_20_26 ? 6'h1a : _T_25644; // @[Mux.scala 31:69:@6678.4]
  assign _T_25646 = valid_20_25 ? 6'h19 : _T_25645; // @[Mux.scala 31:69:@6679.4]
  assign _T_25647 = valid_20_24 ? 6'h18 : _T_25646; // @[Mux.scala 31:69:@6680.4]
  assign _T_25648 = valid_20_23 ? 6'h17 : _T_25647; // @[Mux.scala 31:69:@6681.4]
  assign _T_25649 = valid_20_22 ? 6'h16 : _T_25648; // @[Mux.scala 31:69:@6682.4]
  assign _T_25650 = valid_20_21 ? 6'h15 : _T_25649; // @[Mux.scala 31:69:@6683.4]
  assign _T_25651 = valid_20_20 ? 6'h14 : _T_25650; // @[Mux.scala 31:69:@6684.4]
  assign _T_25652 = valid_20_19 ? 6'h13 : _T_25651; // @[Mux.scala 31:69:@6685.4]
  assign _T_25653 = valid_20_18 ? 6'h12 : _T_25652; // @[Mux.scala 31:69:@6686.4]
  assign _T_25654 = valid_20_17 ? 6'h11 : _T_25653; // @[Mux.scala 31:69:@6687.4]
  assign _T_25655 = valid_20_16 ? 6'h10 : _T_25654; // @[Mux.scala 31:69:@6688.4]
  assign _T_25656 = valid_20_15 ? 6'hf : _T_25655; // @[Mux.scala 31:69:@6689.4]
  assign _T_25657 = valid_20_14 ? 6'he : _T_25656; // @[Mux.scala 31:69:@6690.4]
  assign _T_25658 = valid_20_13 ? 6'hd : _T_25657; // @[Mux.scala 31:69:@6691.4]
  assign _T_25659 = valid_20_12 ? 6'hc : _T_25658; // @[Mux.scala 31:69:@6692.4]
  assign _T_25660 = valid_20_11 ? 6'hb : _T_25659; // @[Mux.scala 31:69:@6693.4]
  assign _T_25661 = valid_20_10 ? 6'ha : _T_25660; // @[Mux.scala 31:69:@6694.4]
  assign _T_25662 = valid_20_9 ? 6'h9 : _T_25661; // @[Mux.scala 31:69:@6695.4]
  assign _T_25663 = valid_20_8 ? 6'h8 : _T_25662; // @[Mux.scala 31:69:@6696.4]
  assign _T_25664 = valid_20_7 ? 6'h7 : _T_25663; // @[Mux.scala 31:69:@6697.4]
  assign _T_25665 = valid_20_6 ? 6'h6 : _T_25664; // @[Mux.scala 31:69:@6698.4]
  assign _T_25666 = valid_20_5 ? 6'h5 : _T_25665; // @[Mux.scala 31:69:@6699.4]
  assign _T_25667 = valid_20_4 ? 6'h4 : _T_25666; // @[Mux.scala 31:69:@6700.4]
  assign _T_25668 = valid_20_3 ? 6'h3 : _T_25667; // @[Mux.scala 31:69:@6701.4]
  assign _T_25669 = valid_20_2 ? 6'h2 : _T_25668; // @[Mux.scala 31:69:@6702.4]
  assign _T_25670 = valid_20_1 ? 6'h1 : _T_25669; // @[Mux.scala 31:69:@6703.4]
  assign select_20 = valid_20_0 ? 6'h0 : _T_25670; // @[Mux.scala 31:69:@6704.4]
  assign _GEN_1281 = 6'h1 == select_20 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1282 = 6'h2 == select_20 ? io_inData_2 : _GEN_1281; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1283 = 6'h3 == select_20 ? io_inData_3 : _GEN_1282; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1284 = 6'h4 == select_20 ? io_inData_4 : _GEN_1283; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1285 = 6'h5 == select_20 ? io_inData_5 : _GEN_1284; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1286 = 6'h6 == select_20 ? io_inData_6 : _GEN_1285; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1287 = 6'h7 == select_20 ? io_inData_7 : _GEN_1286; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1288 = 6'h8 == select_20 ? io_inData_8 : _GEN_1287; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1289 = 6'h9 == select_20 ? io_inData_9 : _GEN_1288; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1290 = 6'ha == select_20 ? io_inData_10 : _GEN_1289; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1291 = 6'hb == select_20 ? io_inData_11 : _GEN_1290; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1292 = 6'hc == select_20 ? io_inData_12 : _GEN_1291; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1293 = 6'hd == select_20 ? io_inData_13 : _GEN_1292; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1294 = 6'he == select_20 ? io_inData_14 : _GEN_1293; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1295 = 6'hf == select_20 ? io_inData_15 : _GEN_1294; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1296 = 6'h10 == select_20 ? io_inData_16 : _GEN_1295; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1297 = 6'h11 == select_20 ? io_inData_17 : _GEN_1296; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1298 = 6'h12 == select_20 ? io_inData_18 : _GEN_1297; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1299 = 6'h13 == select_20 ? io_inData_19 : _GEN_1298; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1300 = 6'h14 == select_20 ? io_inData_20 : _GEN_1299; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1301 = 6'h15 == select_20 ? io_inData_21 : _GEN_1300; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1302 = 6'h16 == select_20 ? io_inData_22 : _GEN_1301; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1303 = 6'h17 == select_20 ? io_inData_23 : _GEN_1302; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1304 = 6'h18 == select_20 ? io_inData_24 : _GEN_1303; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1305 = 6'h19 == select_20 ? io_inData_25 : _GEN_1304; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1306 = 6'h1a == select_20 ? io_inData_26 : _GEN_1305; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1307 = 6'h1b == select_20 ? io_inData_27 : _GEN_1306; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1308 = 6'h1c == select_20 ? io_inData_28 : _GEN_1307; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1309 = 6'h1d == select_20 ? io_inData_29 : _GEN_1308; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1310 = 6'h1e == select_20 ? io_inData_30 : _GEN_1309; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1311 = 6'h1f == select_20 ? io_inData_31 : _GEN_1310; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1312 = 6'h20 == select_20 ? io_inData_32 : _GEN_1311; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1313 = 6'h21 == select_20 ? io_inData_33 : _GEN_1312; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1314 = 6'h22 == select_20 ? io_inData_34 : _GEN_1313; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1315 = 6'h23 == select_20 ? io_inData_35 : _GEN_1314; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1316 = 6'h24 == select_20 ? io_inData_36 : _GEN_1315; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1317 = 6'h25 == select_20 ? io_inData_37 : _GEN_1316; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1318 = 6'h26 == select_20 ? io_inData_38 : _GEN_1317; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1319 = 6'h27 == select_20 ? io_inData_39 : _GEN_1318; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1320 = 6'h28 == select_20 ? io_inData_40 : _GEN_1319; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1321 = 6'h29 == select_20 ? io_inData_41 : _GEN_1320; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1322 = 6'h2a == select_20 ? io_inData_42 : _GEN_1321; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1323 = 6'h2b == select_20 ? io_inData_43 : _GEN_1322; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1324 = 6'h2c == select_20 ? io_inData_44 : _GEN_1323; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1325 = 6'h2d == select_20 ? io_inData_45 : _GEN_1324; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1326 = 6'h2e == select_20 ? io_inData_46 : _GEN_1325; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1327 = 6'h2f == select_20 ? io_inData_47 : _GEN_1326; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1328 = 6'h30 == select_20 ? io_inData_48 : _GEN_1327; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1329 = 6'h31 == select_20 ? io_inData_49 : _GEN_1328; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1330 = 6'h32 == select_20 ? io_inData_50 : _GEN_1329; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1331 = 6'h33 == select_20 ? io_inData_51 : _GEN_1330; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1332 = 6'h34 == select_20 ? io_inData_52 : _GEN_1331; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1333 = 6'h35 == select_20 ? io_inData_53 : _GEN_1332; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1334 = 6'h36 == select_20 ? io_inData_54 : _GEN_1333; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1335 = 6'h37 == select_20 ? io_inData_55 : _GEN_1334; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1336 = 6'h38 == select_20 ? io_inData_56 : _GEN_1335; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1337 = 6'h39 == select_20 ? io_inData_57 : _GEN_1336; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1338 = 6'h3a == select_20 ? io_inData_58 : _GEN_1337; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1339 = 6'h3b == select_20 ? io_inData_59 : _GEN_1338; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1340 = 6'h3c == select_20 ? io_inData_60 : _GEN_1339; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1341 = 6'h3d == select_20 ? io_inData_61 : _GEN_1340; // @[Switch.scala 33:19:@6706.4]
  assign _GEN_1342 = 6'h3e == select_20 ? io_inData_62 : _GEN_1341; // @[Switch.scala 33:19:@6706.4]
  assign _T_25679 = {valid_20_7,valid_20_6,valid_20_5,valid_20_4,valid_20_3,valid_20_2,valid_20_1,valid_20_0}; // @[Switch.scala 34:32:@6713.4]
  assign _T_25687 = {valid_20_15,valid_20_14,valid_20_13,valid_20_12,valid_20_11,valid_20_10,valid_20_9,valid_20_8,_T_25679}; // @[Switch.scala 34:32:@6721.4]
  assign _T_25694 = {valid_20_23,valid_20_22,valid_20_21,valid_20_20,valid_20_19,valid_20_18,valid_20_17,valid_20_16}; // @[Switch.scala 34:32:@6728.4]
  assign _T_25703 = {valid_20_31,valid_20_30,valid_20_29,valid_20_28,valid_20_27,valid_20_26,valid_20_25,valid_20_24,_T_25694,_T_25687}; // @[Switch.scala 34:32:@6737.4]
  assign _T_25710 = {valid_20_39,valid_20_38,valid_20_37,valid_20_36,valid_20_35,valid_20_34,valid_20_33,valid_20_32}; // @[Switch.scala 34:32:@6744.4]
  assign _T_25718 = {valid_20_47,valid_20_46,valid_20_45,valid_20_44,valid_20_43,valid_20_42,valid_20_41,valid_20_40,_T_25710}; // @[Switch.scala 34:32:@6752.4]
  assign _T_25725 = {valid_20_55,valid_20_54,valid_20_53,valid_20_52,valid_20_51,valid_20_50,valid_20_49,valid_20_48}; // @[Switch.scala 34:32:@6759.4]
  assign _T_25734 = {valid_20_63,valid_20_62,valid_20_61,valid_20_60,valid_20_59,valid_20_58,valid_20_57,valid_20_56,_T_25725,_T_25718}; // @[Switch.scala 34:32:@6768.4]
  assign _T_25735 = {_T_25734,_T_25703}; // @[Switch.scala 34:32:@6769.4]
  assign _T_25739 = io_inAddr_0 == 6'h15; // @[Switch.scala 30:53:@6772.4]
  assign valid_21_0 = io_inValid_0 & _T_25739; // @[Switch.scala 30:36:@6773.4]
  assign _T_25742 = io_inAddr_1 == 6'h15; // @[Switch.scala 30:53:@6775.4]
  assign valid_21_1 = io_inValid_1 & _T_25742; // @[Switch.scala 30:36:@6776.4]
  assign _T_25745 = io_inAddr_2 == 6'h15; // @[Switch.scala 30:53:@6778.4]
  assign valid_21_2 = io_inValid_2 & _T_25745; // @[Switch.scala 30:36:@6779.4]
  assign _T_25748 = io_inAddr_3 == 6'h15; // @[Switch.scala 30:53:@6781.4]
  assign valid_21_3 = io_inValid_3 & _T_25748; // @[Switch.scala 30:36:@6782.4]
  assign _T_25751 = io_inAddr_4 == 6'h15; // @[Switch.scala 30:53:@6784.4]
  assign valid_21_4 = io_inValid_4 & _T_25751; // @[Switch.scala 30:36:@6785.4]
  assign _T_25754 = io_inAddr_5 == 6'h15; // @[Switch.scala 30:53:@6787.4]
  assign valid_21_5 = io_inValid_5 & _T_25754; // @[Switch.scala 30:36:@6788.4]
  assign _T_25757 = io_inAddr_6 == 6'h15; // @[Switch.scala 30:53:@6790.4]
  assign valid_21_6 = io_inValid_6 & _T_25757; // @[Switch.scala 30:36:@6791.4]
  assign _T_25760 = io_inAddr_7 == 6'h15; // @[Switch.scala 30:53:@6793.4]
  assign valid_21_7 = io_inValid_7 & _T_25760; // @[Switch.scala 30:36:@6794.4]
  assign _T_25763 = io_inAddr_8 == 6'h15; // @[Switch.scala 30:53:@6796.4]
  assign valid_21_8 = io_inValid_8 & _T_25763; // @[Switch.scala 30:36:@6797.4]
  assign _T_25766 = io_inAddr_9 == 6'h15; // @[Switch.scala 30:53:@6799.4]
  assign valid_21_9 = io_inValid_9 & _T_25766; // @[Switch.scala 30:36:@6800.4]
  assign _T_25769 = io_inAddr_10 == 6'h15; // @[Switch.scala 30:53:@6802.4]
  assign valid_21_10 = io_inValid_10 & _T_25769; // @[Switch.scala 30:36:@6803.4]
  assign _T_25772 = io_inAddr_11 == 6'h15; // @[Switch.scala 30:53:@6805.4]
  assign valid_21_11 = io_inValid_11 & _T_25772; // @[Switch.scala 30:36:@6806.4]
  assign _T_25775 = io_inAddr_12 == 6'h15; // @[Switch.scala 30:53:@6808.4]
  assign valid_21_12 = io_inValid_12 & _T_25775; // @[Switch.scala 30:36:@6809.4]
  assign _T_25778 = io_inAddr_13 == 6'h15; // @[Switch.scala 30:53:@6811.4]
  assign valid_21_13 = io_inValid_13 & _T_25778; // @[Switch.scala 30:36:@6812.4]
  assign _T_25781 = io_inAddr_14 == 6'h15; // @[Switch.scala 30:53:@6814.4]
  assign valid_21_14 = io_inValid_14 & _T_25781; // @[Switch.scala 30:36:@6815.4]
  assign _T_25784 = io_inAddr_15 == 6'h15; // @[Switch.scala 30:53:@6817.4]
  assign valid_21_15 = io_inValid_15 & _T_25784; // @[Switch.scala 30:36:@6818.4]
  assign _T_25787 = io_inAddr_16 == 6'h15; // @[Switch.scala 30:53:@6820.4]
  assign valid_21_16 = io_inValid_16 & _T_25787; // @[Switch.scala 30:36:@6821.4]
  assign _T_25790 = io_inAddr_17 == 6'h15; // @[Switch.scala 30:53:@6823.4]
  assign valid_21_17 = io_inValid_17 & _T_25790; // @[Switch.scala 30:36:@6824.4]
  assign _T_25793 = io_inAddr_18 == 6'h15; // @[Switch.scala 30:53:@6826.4]
  assign valid_21_18 = io_inValid_18 & _T_25793; // @[Switch.scala 30:36:@6827.4]
  assign _T_25796 = io_inAddr_19 == 6'h15; // @[Switch.scala 30:53:@6829.4]
  assign valid_21_19 = io_inValid_19 & _T_25796; // @[Switch.scala 30:36:@6830.4]
  assign _T_25799 = io_inAddr_20 == 6'h15; // @[Switch.scala 30:53:@6832.4]
  assign valid_21_20 = io_inValid_20 & _T_25799; // @[Switch.scala 30:36:@6833.4]
  assign _T_25802 = io_inAddr_21 == 6'h15; // @[Switch.scala 30:53:@6835.4]
  assign valid_21_21 = io_inValid_21 & _T_25802; // @[Switch.scala 30:36:@6836.4]
  assign _T_25805 = io_inAddr_22 == 6'h15; // @[Switch.scala 30:53:@6838.4]
  assign valid_21_22 = io_inValid_22 & _T_25805; // @[Switch.scala 30:36:@6839.4]
  assign _T_25808 = io_inAddr_23 == 6'h15; // @[Switch.scala 30:53:@6841.4]
  assign valid_21_23 = io_inValid_23 & _T_25808; // @[Switch.scala 30:36:@6842.4]
  assign _T_25811 = io_inAddr_24 == 6'h15; // @[Switch.scala 30:53:@6844.4]
  assign valid_21_24 = io_inValid_24 & _T_25811; // @[Switch.scala 30:36:@6845.4]
  assign _T_25814 = io_inAddr_25 == 6'h15; // @[Switch.scala 30:53:@6847.4]
  assign valid_21_25 = io_inValid_25 & _T_25814; // @[Switch.scala 30:36:@6848.4]
  assign _T_25817 = io_inAddr_26 == 6'h15; // @[Switch.scala 30:53:@6850.4]
  assign valid_21_26 = io_inValid_26 & _T_25817; // @[Switch.scala 30:36:@6851.4]
  assign _T_25820 = io_inAddr_27 == 6'h15; // @[Switch.scala 30:53:@6853.4]
  assign valid_21_27 = io_inValid_27 & _T_25820; // @[Switch.scala 30:36:@6854.4]
  assign _T_25823 = io_inAddr_28 == 6'h15; // @[Switch.scala 30:53:@6856.4]
  assign valid_21_28 = io_inValid_28 & _T_25823; // @[Switch.scala 30:36:@6857.4]
  assign _T_25826 = io_inAddr_29 == 6'h15; // @[Switch.scala 30:53:@6859.4]
  assign valid_21_29 = io_inValid_29 & _T_25826; // @[Switch.scala 30:36:@6860.4]
  assign _T_25829 = io_inAddr_30 == 6'h15; // @[Switch.scala 30:53:@6862.4]
  assign valid_21_30 = io_inValid_30 & _T_25829; // @[Switch.scala 30:36:@6863.4]
  assign _T_25832 = io_inAddr_31 == 6'h15; // @[Switch.scala 30:53:@6865.4]
  assign valid_21_31 = io_inValid_31 & _T_25832; // @[Switch.scala 30:36:@6866.4]
  assign _T_25835 = io_inAddr_32 == 6'h15; // @[Switch.scala 30:53:@6868.4]
  assign valid_21_32 = io_inValid_32 & _T_25835; // @[Switch.scala 30:36:@6869.4]
  assign _T_25838 = io_inAddr_33 == 6'h15; // @[Switch.scala 30:53:@6871.4]
  assign valid_21_33 = io_inValid_33 & _T_25838; // @[Switch.scala 30:36:@6872.4]
  assign _T_25841 = io_inAddr_34 == 6'h15; // @[Switch.scala 30:53:@6874.4]
  assign valid_21_34 = io_inValid_34 & _T_25841; // @[Switch.scala 30:36:@6875.4]
  assign _T_25844 = io_inAddr_35 == 6'h15; // @[Switch.scala 30:53:@6877.4]
  assign valid_21_35 = io_inValid_35 & _T_25844; // @[Switch.scala 30:36:@6878.4]
  assign _T_25847 = io_inAddr_36 == 6'h15; // @[Switch.scala 30:53:@6880.4]
  assign valid_21_36 = io_inValid_36 & _T_25847; // @[Switch.scala 30:36:@6881.4]
  assign _T_25850 = io_inAddr_37 == 6'h15; // @[Switch.scala 30:53:@6883.4]
  assign valid_21_37 = io_inValid_37 & _T_25850; // @[Switch.scala 30:36:@6884.4]
  assign _T_25853 = io_inAddr_38 == 6'h15; // @[Switch.scala 30:53:@6886.4]
  assign valid_21_38 = io_inValid_38 & _T_25853; // @[Switch.scala 30:36:@6887.4]
  assign _T_25856 = io_inAddr_39 == 6'h15; // @[Switch.scala 30:53:@6889.4]
  assign valid_21_39 = io_inValid_39 & _T_25856; // @[Switch.scala 30:36:@6890.4]
  assign _T_25859 = io_inAddr_40 == 6'h15; // @[Switch.scala 30:53:@6892.4]
  assign valid_21_40 = io_inValid_40 & _T_25859; // @[Switch.scala 30:36:@6893.4]
  assign _T_25862 = io_inAddr_41 == 6'h15; // @[Switch.scala 30:53:@6895.4]
  assign valid_21_41 = io_inValid_41 & _T_25862; // @[Switch.scala 30:36:@6896.4]
  assign _T_25865 = io_inAddr_42 == 6'h15; // @[Switch.scala 30:53:@6898.4]
  assign valid_21_42 = io_inValid_42 & _T_25865; // @[Switch.scala 30:36:@6899.4]
  assign _T_25868 = io_inAddr_43 == 6'h15; // @[Switch.scala 30:53:@6901.4]
  assign valid_21_43 = io_inValid_43 & _T_25868; // @[Switch.scala 30:36:@6902.4]
  assign _T_25871 = io_inAddr_44 == 6'h15; // @[Switch.scala 30:53:@6904.4]
  assign valid_21_44 = io_inValid_44 & _T_25871; // @[Switch.scala 30:36:@6905.4]
  assign _T_25874 = io_inAddr_45 == 6'h15; // @[Switch.scala 30:53:@6907.4]
  assign valid_21_45 = io_inValid_45 & _T_25874; // @[Switch.scala 30:36:@6908.4]
  assign _T_25877 = io_inAddr_46 == 6'h15; // @[Switch.scala 30:53:@6910.4]
  assign valid_21_46 = io_inValid_46 & _T_25877; // @[Switch.scala 30:36:@6911.4]
  assign _T_25880 = io_inAddr_47 == 6'h15; // @[Switch.scala 30:53:@6913.4]
  assign valid_21_47 = io_inValid_47 & _T_25880; // @[Switch.scala 30:36:@6914.4]
  assign _T_25883 = io_inAddr_48 == 6'h15; // @[Switch.scala 30:53:@6916.4]
  assign valid_21_48 = io_inValid_48 & _T_25883; // @[Switch.scala 30:36:@6917.4]
  assign _T_25886 = io_inAddr_49 == 6'h15; // @[Switch.scala 30:53:@6919.4]
  assign valid_21_49 = io_inValid_49 & _T_25886; // @[Switch.scala 30:36:@6920.4]
  assign _T_25889 = io_inAddr_50 == 6'h15; // @[Switch.scala 30:53:@6922.4]
  assign valid_21_50 = io_inValid_50 & _T_25889; // @[Switch.scala 30:36:@6923.4]
  assign _T_25892 = io_inAddr_51 == 6'h15; // @[Switch.scala 30:53:@6925.4]
  assign valid_21_51 = io_inValid_51 & _T_25892; // @[Switch.scala 30:36:@6926.4]
  assign _T_25895 = io_inAddr_52 == 6'h15; // @[Switch.scala 30:53:@6928.4]
  assign valid_21_52 = io_inValid_52 & _T_25895; // @[Switch.scala 30:36:@6929.4]
  assign _T_25898 = io_inAddr_53 == 6'h15; // @[Switch.scala 30:53:@6931.4]
  assign valid_21_53 = io_inValid_53 & _T_25898; // @[Switch.scala 30:36:@6932.4]
  assign _T_25901 = io_inAddr_54 == 6'h15; // @[Switch.scala 30:53:@6934.4]
  assign valid_21_54 = io_inValid_54 & _T_25901; // @[Switch.scala 30:36:@6935.4]
  assign _T_25904 = io_inAddr_55 == 6'h15; // @[Switch.scala 30:53:@6937.4]
  assign valid_21_55 = io_inValid_55 & _T_25904; // @[Switch.scala 30:36:@6938.4]
  assign _T_25907 = io_inAddr_56 == 6'h15; // @[Switch.scala 30:53:@6940.4]
  assign valid_21_56 = io_inValid_56 & _T_25907; // @[Switch.scala 30:36:@6941.4]
  assign _T_25910 = io_inAddr_57 == 6'h15; // @[Switch.scala 30:53:@6943.4]
  assign valid_21_57 = io_inValid_57 & _T_25910; // @[Switch.scala 30:36:@6944.4]
  assign _T_25913 = io_inAddr_58 == 6'h15; // @[Switch.scala 30:53:@6946.4]
  assign valid_21_58 = io_inValid_58 & _T_25913; // @[Switch.scala 30:36:@6947.4]
  assign _T_25916 = io_inAddr_59 == 6'h15; // @[Switch.scala 30:53:@6949.4]
  assign valid_21_59 = io_inValid_59 & _T_25916; // @[Switch.scala 30:36:@6950.4]
  assign _T_25919 = io_inAddr_60 == 6'h15; // @[Switch.scala 30:53:@6952.4]
  assign valid_21_60 = io_inValid_60 & _T_25919; // @[Switch.scala 30:36:@6953.4]
  assign _T_25922 = io_inAddr_61 == 6'h15; // @[Switch.scala 30:53:@6955.4]
  assign valid_21_61 = io_inValid_61 & _T_25922; // @[Switch.scala 30:36:@6956.4]
  assign _T_25925 = io_inAddr_62 == 6'h15; // @[Switch.scala 30:53:@6958.4]
  assign valid_21_62 = io_inValid_62 & _T_25925; // @[Switch.scala 30:36:@6959.4]
  assign _T_25928 = io_inAddr_63 == 6'h15; // @[Switch.scala 30:53:@6961.4]
  assign valid_21_63 = io_inValid_63 & _T_25928; // @[Switch.scala 30:36:@6962.4]
  assign _T_25994 = valid_21_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@6964.4]
  assign _T_25995 = valid_21_61 ? 6'h3d : _T_25994; // @[Mux.scala 31:69:@6965.4]
  assign _T_25996 = valid_21_60 ? 6'h3c : _T_25995; // @[Mux.scala 31:69:@6966.4]
  assign _T_25997 = valid_21_59 ? 6'h3b : _T_25996; // @[Mux.scala 31:69:@6967.4]
  assign _T_25998 = valid_21_58 ? 6'h3a : _T_25997; // @[Mux.scala 31:69:@6968.4]
  assign _T_25999 = valid_21_57 ? 6'h39 : _T_25998; // @[Mux.scala 31:69:@6969.4]
  assign _T_26000 = valid_21_56 ? 6'h38 : _T_25999; // @[Mux.scala 31:69:@6970.4]
  assign _T_26001 = valid_21_55 ? 6'h37 : _T_26000; // @[Mux.scala 31:69:@6971.4]
  assign _T_26002 = valid_21_54 ? 6'h36 : _T_26001; // @[Mux.scala 31:69:@6972.4]
  assign _T_26003 = valid_21_53 ? 6'h35 : _T_26002; // @[Mux.scala 31:69:@6973.4]
  assign _T_26004 = valid_21_52 ? 6'h34 : _T_26003; // @[Mux.scala 31:69:@6974.4]
  assign _T_26005 = valid_21_51 ? 6'h33 : _T_26004; // @[Mux.scala 31:69:@6975.4]
  assign _T_26006 = valid_21_50 ? 6'h32 : _T_26005; // @[Mux.scala 31:69:@6976.4]
  assign _T_26007 = valid_21_49 ? 6'h31 : _T_26006; // @[Mux.scala 31:69:@6977.4]
  assign _T_26008 = valid_21_48 ? 6'h30 : _T_26007; // @[Mux.scala 31:69:@6978.4]
  assign _T_26009 = valid_21_47 ? 6'h2f : _T_26008; // @[Mux.scala 31:69:@6979.4]
  assign _T_26010 = valid_21_46 ? 6'h2e : _T_26009; // @[Mux.scala 31:69:@6980.4]
  assign _T_26011 = valid_21_45 ? 6'h2d : _T_26010; // @[Mux.scala 31:69:@6981.4]
  assign _T_26012 = valid_21_44 ? 6'h2c : _T_26011; // @[Mux.scala 31:69:@6982.4]
  assign _T_26013 = valid_21_43 ? 6'h2b : _T_26012; // @[Mux.scala 31:69:@6983.4]
  assign _T_26014 = valid_21_42 ? 6'h2a : _T_26013; // @[Mux.scala 31:69:@6984.4]
  assign _T_26015 = valid_21_41 ? 6'h29 : _T_26014; // @[Mux.scala 31:69:@6985.4]
  assign _T_26016 = valid_21_40 ? 6'h28 : _T_26015; // @[Mux.scala 31:69:@6986.4]
  assign _T_26017 = valid_21_39 ? 6'h27 : _T_26016; // @[Mux.scala 31:69:@6987.4]
  assign _T_26018 = valid_21_38 ? 6'h26 : _T_26017; // @[Mux.scala 31:69:@6988.4]
  assign _T_26019 = valid_21_37 ? 6'h25 : _T_26018; // @[Mux.scala 31:69:@6989.4]
  assign _T_26020 = valid_21_36 ? 6'h24 : _T_26019; // @[Mux.scala 31:69:@6990.4]
  assign _T_26021 = valid_21_35 ? 6'h23 : _T_26020; // @[Mux.scala 31:69:@6991.4]
  assign _T_26022 = valid_21_34 ? 6'h22 : _T_26021; // @[Mux.scala 31:69:@6992.4]
  assign _T_26023 = valid_21_33 ? 6'h21 : _T_26022; // @[Mux.scala 31:69:@6993.4]
  assign _T_26024 = valid_21_32 ? 6'h20 : _T_26023; // @[Mux.scala 31:69:@6994.4]
  assign _T_26025 = valid_21_31 ? 6'h1f : _T_26024; // @[Mux.scala 31:69:@6995.4]
  assign _T_26026 = valid_21_30 ? 6'h1e : _T_26025; // @[Mux.scala 31:69:@6996.4]
  assign _T_26027 = valid_21_29 ? 6'h1d : _T_26026; // @[Mux.scala 31:69:@6997.4]
  assign _T_26028 = valid_21_28 ? 6'h1c : _T_26027; // @[Mux.scala 31:69:@6998.4]
  assign _T_26029 = valid_21_27 ? 6'h1b : _T_26028; // @[Mux.scala 31:69:@6999.4]
  assign _T_26030 = valid_21_26 ? 6'h1a : _T_26029; // @[Mux.scala 31:69:@7000.4]
  assign _T_26031 = valid_21_25 ? 6'h19 : _T_26030; // @[Mux.scala 31:69:@7001.4]
  assign _T_26032 = valid_21_24 ? 6'h18 : _T_26031; // @[Mux.scala 31:69:@7002.4]
  assign _T_26033 = valid_21_23 ? 6'h17 : _T_26032; // @[Mux.scala 31:69:@7003.4]
  assign _T_26034 = valid_21_22 ? 6'h16 : _T_26033; // @[Mux.scala 31:69:@7004.4]
  assign _T_26035 = valid_21_21 ? 6'h15 : _T_26034; // @[Mux.scala 31:69:@7005.4]
  assign _T_26036 = valid_21_20 ? 6'h14 : _T_26035; // @[Mux.scala 31:69:@7006.4]
  assign _T_26037 = valid_21_19 ? 6'h13 : _T_26036; // @[Mux.scala 31:69:@7007.4]
  assign _T_26038 = valid_21_18 ? 6'h12 : _T_26037; // @[Mux.scala 31:69:@7008.4]
  assign _T_26039 = valid_21_17 ? 6'h11 : _T_26038; // @[Mux.scala 31:69:@7009.4]
  assign _T_26040 = valid_21_16 ? 6'h10 : _T_26039; // @[Mux.scala 31:69:@7010.4]
  assign _T_26041 = valid_21_15 ? 6'hf : _T_26040; // @[Mux.scala 31:69:@7011.4]
  assign _T_26042 = valid_21_14 ? 6'he : _T_26041; // @[Mux.scala 31:69:@7012.4]
  assign _T_26043 = valid_21_13 ? 6'hd : _T_26042; // @[Mux.scala 31:69:@7013.4]
  assign _T_26044 = valid_21_12 ? 6'hc : _T_26043; // @[Mux.scala 31:69:@7014.4]
  assign _T_26045 = valid_21_11 ? 6'hb : _T_26044; // @[Mux.scala 31:69:@7015.4]
  assign _T_26046 = valid_21_10 ? 6'ha : _T_26045; // @[Mux.scala 31:69:@7016.4]
  assign _T_26047 = valid_21_9 ? 6'h9 : _T_26046; // @[Mux.scala 31:69:@7017.4]
  assign _T_26048 = valid_21_8 ? 6'h8 : _T_26047; // @[Mux.scala 31:69:@7018.4]
  assign _T_26049 = valid_21_7 ? 6'h7 : _T_26048; // @[Mux.scala 31:69:@7019.4]
  assign _T_26050 = valid_21_6 ? 6'h6 : _T_26049; // @[Mux.scala 31:69:@7020.4]
  assign _T_26051 = valid_21_5 ? 6'h5 : _T_26050; // @[Mux.scala 31:69:@7021.4]
  assign _T_26052 = valid_21_4 ? 6'h4 : _T_26051; // @[Mux.scala 31:69:@7022.4]
  assign _T_26053 = valid_21_3 ? 6'h3 : _T_26052; // @[Mux.scala 31:69:@7023.4]
  assign _T_26054 = valid_21_2 ? 6'h2 : _T_26053; // @[Mux.scala 31:69:@7024.4]
  assign _T_26055 = valid_21_1 ? 6'h1 : _T_26054; // @[Mux.scala 31:69:@7025.4]
  assign select_21 = valid_21_0 ? 6'h0 : _T_26055; // @[Mux.scala 31:69:@7026.4]
  assign _GEN_1345 = 6'h1 == select_21 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1346 = 6'h2 == select_21 ? io_inData_2 : _GEN_1345; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1347 = 6'h3 == select_21 ? io_inData_3 : _GEN_1346; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1348 = 6'h4 == select_21 ? io_inData_4 : _GEN_1347; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1349 = 6'h5 == select_21 ? io_inData_5 : _GEN_1348; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1350 = 6'h6 == select_21 ? io_inData_6 : _GEN_1349; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1351 = 6'h7 == select_21 ? io_inData_7 : _GEN_1350; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1352 = 6'h8 == select_21 ? io_inData_8 : _GEN_1351; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1353 = 6'h9 == select_21 ? io_inData_9 : _GEN_1352; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1354 = 6'ha == select_21 ? io_inData_10 : _GEN_1353; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1355 = 6'hb == select_21 ? io_inData_11 : _GEN_1354; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1356 = 6'hc == select_21 ? io_inData_12 : _GEN_1355; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1357 = 6'hd == select_21 ? io_inData_13 : _GEN_1356; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1358 = 6'he == select_21 ? io_inData_14 : _GEN_1357; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1359 = 6'hf == select_21 ? io_inData_15 : _GEN_1358; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1360 = 6'h10 == select_21 ? io_inData_16 : _GEN_1359; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1361 = 6'h11 == select_21 ? io_inData_17 : _GEN_1360; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1362 = 6'h12 == select_21 ? io_inData_18 : _GEN_1361; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1363 = 6'h13 == select_21 ? io_inData_19 : _GEN_1362; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1364 = 6'h14 == select_21 ? io_inData_20 : _GEN_1363; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1365 = 6'h15 == select_21 ? io_inData_21 : _GEN_1364; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1366 = 6'h16 == select_21 ? io_inData_22 : _GEN_1365; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1367 = 6'h17 == select_21 ? io_inData_23 : _GEN_1366; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1368 = 6'h18 == select_21 ? io_inData_24 : _GEN_1367; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1369 = 6'h19 == select_21 ? io_inData_25 : _GEN_1368; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1370 = 6'h1a == select_21 ? io_inData_26 : _GEN_1369; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1371 = 6'h1b == select_21 ? io_inData_27 : _GEN_1370; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1372 = 6'h1c == select_21 ? io_inData_28 : _GEN_1371; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1373 = 6'h1d == select_21 ? io_inData_29 : _GEN_1372; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1374 = 6'h1e == select_21 ? io_inData_30 : _GEN_1373; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1375 = 6'h1f == select_21 ? io_inData_31 : _GEN_1374; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1376 = 6'h20 == select_21 ? io_inData_32 : _GEN_1375; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1377 = 6'h21 == select_21 ? io_inData_33 : _GEN_1376; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1378 = 6'h22 == select_21 ? io_inData_34 : _GEN_1377; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1379 = 6'h23 == select_21 ? io_inData_35 : _GEN_1378; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1380 = 6'h24 == select_21 ? io_inData_36 : _GEN_1379; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1381 = 6'h25 == select_21 ? io_inData_37 : _GEN_1380; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1382 = 6'h26 == select_21 ? io_inData_38 : _GEN_1381; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1383 = 6'h27 == select_21 ? io_inData_39 : _GEN_1382; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1384 = 6'h28 == select_21 ? io_inData_40 : _GEN_1383; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1385 = 6'h29 == select_21 ? io_inData_41 : _GEN_1384; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1386 = 6'h2a == select_21 ? io_inData_42 : _GEN_1385; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1387 = 6'h2b == select_21 ? io_inData_43 : _GEN_1386; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1388 = 6'h2c == select_21 ? io_inData_44 : _GEN_1387; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1389 = 6'h2d == select_21 ? io_inData_45 : _GEN_1388; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1390 = 6'h2e == select_21 ? io_inData_46 : _GEN_1389; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1391 = 6'h2f == select_21 ? io_inData_47 : _GEN_1390; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1392 = 6'h30 == select_21 ? io_inData_48 : _GEN_1391; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1393 = 6'h31 == select_21 ? io_inData_49 : _GEN_1392; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1394 = 6'h32 == select_21 ? io_inData_50 : _GEN_1393; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1395 = 6'h33 == select_21 ? io_inData_51 : _GEN_1394; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1396 = 6'h34 == select_21 ? io_inData_52 : _GEN_1395; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1397 = 6'h35 == select_21 ? io_inData_53 : _GEN_1396; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1398 = 6'h36 == select_21 ? io_inData_54 : _GEN_1397; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1399 = 6'h37 == select_21 ? io_inData_55 : _GEN_1398; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1400 = 6'h38 == select_21 ? io_inData_56 : _GEN_1399; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1401 = 6'h39 == select_21 ? io_inData_57 : _GEN_1400; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1402 = 6'h3a == select_21 ? io_inData_58 : _GEN_1401; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1403 = 6'h3b == select_21 ? io_inData_59 : _GEN_1402; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1404 = 6'h3c == select_21 ? io_inData_60 : _GEN_1403; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1405 = 6'h3d == select_21 ? io_inData_61 : _GEN_1404; // @[Switch.scala 33:19:@7028.4]
  assign _GEN_1406 = 6'h3e == select_21 ? io_inData_62 : _GEN_1405; // @[Switch.scala 33:19:@7028.4]
  assign _T_26064 = {valid_21_7,valid_21_6,valid_21_5,valid_21_4,valid_21_3,valid_21_2,valid_21_1,valid_21_0}; // @[Switch.scala 34:32:@7035.4]
  assign _T_26072 = {valid_21_15,valid_21_14,valid_21_13,valid_21_12,valid_21_11,valid_21_10,valid_21_9,valid_21_8,_T_26064}; // @[Switch.scala 34:32:@7043.4]
  assign _T_26079 = {valid_21_23,valid_21_22,valid_21_21,valid_21_20,valid_21_19,valid_21_18,valid_21_17,valid_21_16}; // @[Switch.scala 34:32:@7050.4]
  assign _T_26088 = {valid_21_31,valid_21_30,valid_21_29,valid_21_28,valid_21_27,valid_21_26,valid_21_25,valid_21_24,_T_26079,_T_26072}; // @[Switch.scala 34:32:@7059.4]
  assign _T_26095 = {valid_21_39,valid_21_38,valid_21_37,valid_21_36,valid_21_35,valid_21_34,valid_21_33,valid_21_32}; // @[Switch.scala 34:32:@7066.4]
  assign _T_26103 = {valid_21_47,valid_21_46,valid_21_45,valid_21_44,valid_21_43,valid_21_42,valid_21_41,valid_21_40,_T_26095}; // @[Switch.scala 34:32:@7074.4]
  assign _T_26110 = {valid_21_55,valid_21_54,valid_21_53,valid_21_52,valid_21_51,valid_21_50,valid_21_49,valid_21_48}; // @[Switch.scala 34:32:@7081.4]
  assign _T_26119 = {valid_21_63,valid_21_62,valid_21_61,valid_21_60,valid_21_59,valid_21_58,valid_21_57,valid_21_56,_T_26110,_T_26103}; // @[Switch.scala 34:32:@7090.4]
  assign _T_26120 = {_T_26119,_T_26088}; // @[Switch.scala 34:32:@7091.4]
  assign _T_26124 = io_inAddr_0 == 6'h16; // @[Switch.scala 30:53:@7094.4]
  assign valid_22_0 = io_inValid_0 & _T_26124; // @[Switch.scala 30:36:@7095.4]
  assign _T_26127 = io_inAddr_1 == 6'h16; // @[Switch.scala 30:53:@7097.4]
  assign valid_22_1 = io_inValid_1 & _T_26127; // @[Switch.scala 30:36:@7098.4]
  assign _T_26130 = io_inAddr_2 == 6'h16; // @[Switch.scala 30:53:@7100.4]
  assign valid_22_2 = io_inValid_2 & _T_26130; // @[Switch.scala 30:36:@7101.4]
  assign _T_26133 = io_inAddr_3 == 6'h16; // @[Switch.scala 30:53:@7103.4]
  assign valid_22_3 = io_inValid_3 & _T_26133; // @[Switch.scala 30:36:@7104.4]
  assign _T_26136 = io_inAddr_4 == 6'h16; // @[Switch.scala 30:53:@7106.4]
  assign valid_22_4 = io_inValid_4 & _T_26136; // @[Switch.scala 30:36:@7107.4]
  assign _T_26139 = io_inAddr_5 == 6'h16; // @[Switch.scala 30:53:@7109.4]
  assign valid_22_5 = io_inValid_5 & _T_26139; // @[Switch.scala 30:36:@7110.4]
  assign _T_26142 = io_inAddr_6 == 6'h16; // @[Switch.scala 30:53:@7112.4]
  assign valid_22_6 = io_inValid_6 & _T_26142; // @[Switch.scala 30:36:@7113.4]
  assign _T_26145 = io_inAddr_7 == 6'h16; // @[Switch.scala 30:53:@7115.4]
  assign valid_22_7 = io_inValid_7 & _T_26145; // @[Switch.scala 30:36:@7116.4]
  assign _T_26148 = io_inAddr_8 == 6'h16; // @[Switch.scala 30:53:@7118.4]
  assign valid_22_8 = io_inValid_8 & _T_26148; // @[Switch.scala 30:36:@7119.4]
  assign _T_26151 = io_inAddr_9 == 6'h16; // @[Switch.scala 30:53:@7121.4]
  assign valid_22_9 = io_inValid_9 & _T_26151; // @[Switch.scala 30:36:@7122.4]
  assign _T_26154 = io_inAddr_10 == 6'h16; // @[Switch.scala 30:53:@7124.4]
  assign valid_22_10 = io_inValid_10 & _T_26154; // @[Switch.scala 30:36:@7125.4]
  assign _T_26157 = io_inAddr_11 == 6'h16; // @[Switch.scala 30:53:@7127.4]
  assign valid_22_11 = io_inValid_11 & _T_26157; // @[Switch.scala 30:36:@7128.4]
  assign _T_26160 = io_inAddr_12 == 6'h16; // @[Switch.scala 30:53:@7130.4]
  assign valid_22_12 = io_inValid_12 & _T_26160; // @[Switch.scala 30:36:@7131.4]
  assign _T_26163 = io_inAddr_13 == 6'h16; // @[Switch.scala 30:53:@7133.4]
  assign valid_22_13 = io_inValid_13 & _T_26163; // @[Switch.scala 30:36:@7134.4]
  assign _T_26166 = io_inAddr_14 == 6'h16; // @[Switch.scala 30:53:@7136.4]
  assign valid_22_14 = io_inValid_14 & _T_26166; // @[Switch.scala 30:36:@7137.4]
  assign _T_26169 = io_inAddr_15 == 6'h16; // @[Switch.scala 30:53:@7139.4]
  assign valid_22_15 = io_inValid_15 & _T_26169; // @[Switch.scala 30:36:@7140.4]
  assign _T_26172 = io_inAddr_16 == 6'h16; // @[Switch.scala 30:53:@7142.4]
  assign valid_22_16 = io_inValid_16 & _T_26172; // @[Switch.scala 30:36:@7143.4]
  assign _T_26175 = io_inAddr_17 == 6'h16; // @[Switch.scala 30:53:@7145.4]
  assign valid_22_17 = io_inValid_17 & _T_26175; // @[Switch.scala 30:36:@7146.4]
  assign _T_26178 = io_inAddr_18 == 6'h16; // @[Switch.scala 30:53:@7148.4]
  assign valid_22_18 = io_inValid_18 & _T_26178; // @[Switch.scala 30:36:@7149.4]
  assign _T_26181 = io_inAddr_19 == 6'h16; // @[Switch.scala 30:53:@7151.4]
  assign valid_22_19 = io_inValid_19 & _T_26181; // @[Switch.scala 30:36:@7152.4]
  assign _T_26184 = io_inAddr_20 == 6'h16; // @[Switch.scala 30:53:@7154.4]
  assign valid_22_20 = io_inValid_20 & _T_26184; // @[Switch.scala 30:36:@7155.4]
  assign _T_26187 = io_inAddr_21 == 6'h16; // @[Switch.scala 30:53:@7157.4]
  assign valid_22_21 = io_inValid_21 & _T_26187; // @[Switch.scala 30:36:@7158.4]
  assign _T_26190 = io_inAddr_22 == 6'h16; // @[Switch.scala 30:53:@7160.4]
  assign valid_22_22 = io_inValid_22 & _T_26190; // @[Switch.scala 30:36:@7161.4]
  assign _T_26193 = io_inAddr_23 == 6'h16; // @[Switch.scala 30:53:@7163.4]
  assign valid_22_23 = io_inValid_23 & _T_26193; // @[Switch.scala 30:36:@7164.4]
  assign _T_26196 = io_inAddr_24 == 6'h16; // @[Switch.scala 30:53:@7166.4]
  assign valid_22_24 = io_inValid_24 & _T_26196; // @[Switch.scala 30:36:@7167.4]
  assign _T_26199 = io_inAddr_25 == 6'h16; // @[Switch.scala 30:53:@7169.4]
  assign valid_22_25 = io_inValid_25 & _T_26199; // @[Switch.scala 30:36:@7170.4]
  assign _T_26202 = io_inAddr_26 == 6'h16; // @[Switch.scala 30:53:@7172.4]
  assign valid_22_26 = io_inValid_26 & _T_26202; // @[Switch.scala 30:36:@7173.4]
  assign _T_26205 = io_inAddr_27 == 6'h16; // @[Switch.scala 30:53:@7175.4]
  assign valid_22_27 = io_inValid_27 & _T_26205; // @[Switch.scala 30:36:@7176.4]
  assign _T_26208 = io_inAddr_28 == 6'h16; // @[Switch.scala 30:53:@7178.4]
  assign valid_22_28 = io_inValid_28 & _T_26208; // @[Switch.scala 30:36:@7179.4]
  assign _T_26211 = io_inAddr_29 == 6'h16; // @[Switch.scala 30:53:@7181.4]
  assign valid_22_29 = io_inValid_29 & _T_26211; // @[Switch.scala 30:36:@7182.4]
  assign _T_26214 = io_inAddr_30 == 6'h16; // @[Switch.scala 30:53:@7184.4]
  assign valid_22_30 = io_inValid_30 & _T_26214; // @[Switch.scala 30:36:@7185.4]
  assign _T_26217 = io_inAddr_31 == 6'h16; // @[Switch.scala 30:53:@7187.4]
  assign valid_22_31 = io_inValid_31 & _T_26217; // @[Switch.scala 30:36:@7188.4]
  assign _T_26220 = io_inAddr_32 == 6'h16; // @[Switch.scala 30:53:@7190.4]
  assign valid_22_32 = io_inValid_32 & _T_26220; // @[Switch.scala 30:36:@7191.4]
  assign _T_26223 = io_inAddr_33 == 6'h16; // @[Switch.scala 30:53:@7193.4]
  assign valid_22_33 = io_inValid_33 & _T_26223; // @[Switch.scala 30:36:@7194.4]
  assign _T_26226 = io_inAddr_34 == 6'h16; // @[Switch.scala 30:53:@7196.4]
  assign valid_22_34 = io_inValid_34 & _T_26226; // @[Switch.scala 30:36:@7197.4]
  assign _T_26229 = io_inAddr_35 == 6'h16; // @[Switch.scala 30:53:@7199.4]
  assign valid_22_35 = io_inValid_35 & _T_26229; // @[Switch.scala 30:36:@7200.4]
  assign _T_26232 = io_inAddr_36 == 6'h16; // @[Switch.scala 30:53:@7202.4]
  assign valid_22_36 = io_inValid_36 & _T_26232; // @[Switch.scala 30:36:@7203.4]
  assign _T_26235 = io_inAddr_37 == 6'h16; // @[Switch.scala 30:53:@7205.4]
  assign valid_22_37 = io_inValid_37 & _T_26235; // @[Switch.scala 30:36:@7206.4]
  assign _T_26238 = io_inAddr_38 == 6'h16; // @[Switch.scala 30:53:@7208.4]
  assign valid_22_38 = io_inValid_38 & _T_26238; // @[Switch.scala 30:36:@7209.4]
  assign _T_26241 = io_inAddr_39 == 6'h16; // @[Switch.scala 30:53:@7211.4]
  assign valid_22_39 = io_inValid_39 & _T_26241; // @[Switch.scala 30:36:@7212.4]
  assign _T_26244 = io_inAddr_40 == 6'h16; // @[Switch.scala 30:53:@7214.4]
  assign valid_22_40 = io_inValid_40 & _T_26244; // @[Switch.scala 30:36:@7215.4]
  assign _T_26247 = io_inAddr_41 == 6'h16; // @[Switch.scala 30:53:@7217.4]
  assign valid_22_41 = io_inValid_41 & _T_26247; // @[Switch.scala 30:36:@7218.4]
  assign _T_26250 = io_inAddr_42 == 6'h16; // @[Switch.scala 30:53:@7220.4]
  assign valid_22_42 = io_inValid_42 & _T_26250; // @[Switch.scala 30:36:@7221.4]
  assign _T_26253 = io_inAddr_43 == 6'h16; // @[Switch.scala 30:53:@7223.4]
  assign valid_22_43 = io_inValid_43 & _T_26253; // @[Switch.scala 30:36:@7224.4]
  assign _T_26256 = io_inAddr_44 == 6'h16; // @[Switch.scala 30:53:@7226.4]
  assign valid_22_44 = io_inValid_44 & _T_26256; // @[Switch.scala 30:36:@7227.4]
  assign _T_26259 = io_inAddr_45 == 6'h16; // @[Switch.scala 30:53:@7229.4]
  assign valid_22_45 = io_inValid_45 & _T_26259; // @[Switch.scala 30:36:@7230.4]
  assign _T_26262 = io_inAddr_46 == 6'h16; // @[Switch.scala 30:53:@7232.4]
  assign valid_22_46 = io_inValid_46 & _T_26262; // @[Switch.scala 30:36:@7233.4]
  assign _T_26265 = io_inAddr_47 == 6'h16; // @[Switch.scala 30:53:@7235.4]
  assign valid_22_47 = io_inValid_47 & _T_26265; // @[Switch.scala 30:36:@7236.4]
  assign _T_26268 = io_inAddr_48 == 6'h16; // @[Switch.scala 30:53:@7238.4]
  assign valid_22_48 = io_inValid_48 & _T_26268; // @[Switch.scala 30:36:@7239.4]
  assign _T_26271 = io_inAddr_49 == 6'h16; // @[Switch.scala 30:53:@7241.4]
  assign valid_22_49 = io_inValid_49 & _T_26271; // @[Switch.scala 30:36:@7242.4]
  assign _T_26274 = io_inAddr_50 == 6'h16; // @[Switch.scala 30:53:@7244.4]
  assign valid_22_50 = io_inValid_50 & _T_26274; // @[Switch.scala 30:36:@7245.4]
  assign _T_26277 = io_inAddr_51 == 6'h16; // @[Switch.scala 30:53:@7247.4]
  assign valid_22_51 = io_inValid_51 & _T_26277; // @[Switch.scala 30:36:@7248.4]
  assign _T_26280 = io_inAddr_52 == 6'h16; // @[Switch.scala 30:53:@7250.4]
  assign valid_22_52 = io_inValid_52 & _T_26280; // @[Switch.scala 30:36:@7251.4]
  assign _T_26283 = io_inAddr_53 == 6'h16; // @[Switch.scala 30:53:@7253.4]
  assign valid_22_53 = io_inValid_53 & _T_26283; // @[Switch.scala 30:36:@7254.4]
  assign _T_26286 = io_inAddr_54 == 6'h16; // @[Switch.scala 30:53:@7256.4]
  assign valid_22_54 = io_inValid_54 & _T_26286; // @[Switch.scala 30:36:@7257.4]
  assign _T_26289 = io_inAddr_55 == 6'h16; // @[Switch.scala 30:53:@7259.4]
  assign valid_22_55 = io_inValid_55 & _T_26289; // @[Switch.scala 30:36:@7260.4]
  assign _T_26292 = io_inAddr_56 == 6'h16; // @[Switch.scala 30:53:@7262.4]
  assign valid_22_56 = io_inValid_56 & _T_26292; // @[Switch.scala 30:36:@7263.4]
  assign _T_26295 = io_inAddr_57 == 6'h16; // @[Switch.scala 30:53:@7265.4]
  assign valid_22_57 = io_inValid_57 & _T_26295; // @[Switch.scala 30:36:@7266.4]
  assign _T_26298 = io_inAddr_58 == 6'h16; // @[Switch.scala 30:53:@7268.4]
  assign valid_22_58 = io_inValid_58 & _T_26298; // @[Switch.scala 30:36:@7269.4]
  assign _T_26301 = io_inAddr_59 == 6'h16; // @[Switch.scala 30:53:@7271.4]
  assign valid_22_59 = io_inValid_59 & _T_26301; // @[Switch.scala 30:36:@7272.4]
  assign _T_26304 = io_inAddr_60 == 6'h16; // @[Switch.scala 30:53:@7274.4]
  assign valid_22_60 = io_inValid_60 & _T_26304; // @[Switch.scala 30:36:@7275.4]
  assign _T_26307 = io_inAddr_61 == 6'h16; // @[Switch.scala 30:53:@7277.4]
  assign valid_22_61 = io_inValid_61 & _T_26307; // @[Switch.scala 30:36:@7278.4]
  assign _T_26310 = io_inAddr_62 == 6'h16; // @[Switch.scala 30:53:@7280.4]
  assign valid_22_62 = io_inValid_62 & _T_26310; // @[Switch.scala 30:36:@7281.4]
  assign _T_26313 = io_inAddr_63 == 6'h16; // @[Switch.scala 30:53:@7283.4]
  assign valid_22_63 = io_inValid_63 & _T_26313; // @[Switch.scala 30:36:@7284.4]
  assign _T_26379 = valid_22_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@7286.4]
  assign _T_26380 = valid_22_61 ? 6'h3d : _T_26379; // @[Mux.scala 31:69:@7287.4]
  assign _T_26381 = valid_22_60 ? 6'h3c : _T_26380; // @[Mux.scala 31:69:@7288.4]
  assign _T_26382 = valid_22_59 ? 6'h3b : _T_26381; // @[Mux.scala 31:69:@7289.4]
  assign _T_26383 = valid_22_58 ? 6'h3a : _T_26382; // @[Mux.scala 31:69:@7290.4]
  assign _T_26384 = valid_22_57 ? 6'h39 : _T_26383; // @[Mux.scala 31:69:@7291.4]
  assign _T_26385 = valid_22_56 ? 6'h38 : _T_26384; // @[Mux.scala 31:69:@7292.4]
  assign _T_26386 = valid_22_55 ? 6'h37 : _T_26385; // @[Mux.scala 31:69:@7293.4]
  assign _T_26387 = valid_22_54 ? 6'h36 : _T_26386; // @[Mux.scala 31:69:@7294.4]
  assign _T_26388 = valid_22_53 ? 6'h35 : _T_26387; // @[Mux.scala 31:69:@7295.4]
  assign _T_26389 = valid_22_52 ? 6'h34 : _T_26388; // @[Mux.scala 31:69:@7296.4]
  assign _T_26390 = valid_22_51 ? 6'h33 : _T_26389; // @[Mux.scala 31:69:@7297.4]
  assign _T_26391 = valid_22_50 ? 6'h32 : _T_26390; // @[Mux.scala 31:69:@7298.4]
  assign _T_26392 = valid_22_49 ? 6'h31 : _T_26391; // @[Mux.scala 31:69:@7299.4]
  assign _T_26393 = valid_22_48 ? 6'h30 : _T_26392; // @[Mux.scala 31:69:@7300.4]
  assign _T_26394 = valid_22_47 ? 6'h2f : _T_26393; // @[Mux.scala 31:69:@7301.4]
  assign _T_26395 = valid_22_46 ? 6'h2e : _T_26394; // @[Mux.scala 31:69:@7302.4]
  assign _T_26396 = valid_22_45 ? 6'h2d : _T_26395; // @[Mux.scala 31:69:@7303.4]
  assign _T_26397 = valid_22_44 ? 6'h2c : _T_26396; // @[Mux.scala 31:69:@7304.4]
  assign _T_26398 = valid_22_43 ? 6'h2b : _T_26397; // @[Mux.scala 31:69:@7305.4]
  assign _T_26399 = valid_22_42 ? 6'h2a : _T_26398; // @[Mux.scala 31:69:@7306.4]
  assign _T_26400 = valid_22_41 ? 6'h29 : _T_26399; // @[Mux.scala 31:69:@7307.4]
  assign _T_26401 = valid_22_40 ? 6'h28 : _T_26400; // @[Mux.scala 31:69:@7308.4]
  assign _T_26402 = valid_22_39 ? 6'h27 : _T_26401; // @[Mux.scala 31:69:@7309.4]
  assign _T_26403 = valid_22_38 ? 6'h26 : _T_26402; // @[Mux.scala 31:69:@7310.4]
  assign _T_26404 = valid_22_37 ? 6'h25 : _T_26403; // @[Mux.scala 31:69:@7311.4]
  assign _T_26405 = valid_22_36 ? 6'h24 : _T_26404; // @[Mux.scala 31:69:@7312.4]
  assign _T_26406 = valid_22_35 ? 6'h23 : _T_26405; // @[Mux.scala 31:69:@7313.4]
  assign _T_26407 = valid_22_34 ? 6'h22 : _T_26406; // @[Mux.scala 31:69:@7314.4]
  assign _T_26408 = valid_22_33 ? 6'h21 : _T_26407; // @[Mux.scala 31:69:@7315.4]
  assign _T_26409 = valid_22_32 ? 6'h20 : _T_26408; // @[Mux.scala 31:69:@7316.4]
  assign _T_26410 = valid_22_31 ? 6'h1f : _T_26409; // @[Mux.scala 31:69:@7317.4]
  assign _T_26411 = valid_22_30 ? 6'h1e : _T_26410; // @[Mux.scala 31:69:@7318.4]
  assign _T_26412 = valid_22_29 ? 6'h1d : _T_26411; // @[Mux.scala 31:69:@7319.4]
  assign _T_26413 = valid_22_28 ? 6'h1c : _T_26412; // @[Mux.scala 31:69:@7320.4]
  assign _T_26414 = valid_22_27 ? 6'h1b : _T_26413; // @[Mux.scala 31:69:@7321.4]
  assign _T_26415 = valid_22_26 ? 6'h1a : _T_26414; // @[Mux.scala 31:69:@7322.4]
  assign _T_26416 = valid_22_25 ? 6'h19 : _T_26415; // @[Mux.scala 31:69:@7323.4]
  assign _T_26417 = valid_22_24 ? 6'h18 : _T_26416; // @[Mux.scala 31:69:@7324.4]
  assign _T_26418 = valid_22_23 ? 6'h17 : _T_26417; // @[Mux.scala 31:69:@7325.4]
  assign _T_26419 = valid_22_22 ? 6'h16 : _T_26418; // @[Mux.scala 31:69:@7326.4]
  assign _T_26420 = valid_22_21 ? 6'h15 : _T_26419; // @[Mux.scala 31:69:@7327.4]
  assign _T_26421 = valid_22_20 ? 6'h14 : _T_26420; // @[Mux.scala 31:69:@7328.4]
  assign _T_26422 = valid_22_19 ? 6'h13 : _T_26421; // @[Mux.scala 31:69:@7329.4]
  assign _T_26423 = valid_22_18 ? 6'h12 : _T_26422; // @[Mux.scala 31:69:@7330.4]
  assign _T_26424 = valid_22_17 ? 6'h11 : _T_26423; // @[Mux.scala 31:69:@7331.4]
  assign _T_26425 = valid_22_16 ? 6'h10 : _T_26424; // @[Mux.scala 31:69:@7332.4]
  assign _T_26426 = valid_22_15 ? 6'hf : _T_26425; // @[Mux.scala 31:69:@7333.4]
  assign _T_26427 = valid_22_14 ? 6'he : _T_26426; // @[Mux.scala 31:69:@7334.4]
  assign _T_26428 = valid_22_13 ? 6'hd : _T_26427; // @[Mux.scala 31:69:@7335.4]
  assign _T_26429 = valid_22_12 ? 6'hc : _T_26428; // @[Mux.scala 31:69:@7336.4]
  assign _T_26430 = valid_22_11 ? 6'hb : _T_26429; // @[Mux.scala 31:69:@7337.4]
  assign _T_26431 = valid_22_10 ? 6'ha : _T_26430; // @[Mux.scala 31:69:@7338.4]
  assign _T_26432 = valid_22_9 ? 6'h9 : _T_26431; // @[Mux.scala 31:69:@7339.4]
  assign _T_26433 = valid_22_8 ? 6'h8 : _T_26432; // @[Mux.scala 31:69:@7340.4]
  assign _T_26434 = valid_22_7 ? 6'h7 : _T_26433; // @[Mux.scala 31:69:@7341.4]
  assign _T_26435 = valid_22_6 ? 6'h6 : _T_26434; // @[Mux.scala 31:69:@7342.4]
  assign _T_26436 = valid_22_5 ? 6'h5 : _T_26435; // @[Mux.scala 31:69:@7343.4]
  assign _T_26437 = valid_22_4 ? 6'h4 : _T_26436; // @[Mux.scala 31:69:@7344.4]
  assign _T_26438 = valid_22_3 ? 6'h3 : _T_26437; // @[Mux.scala 31:69:@7345.4]
  assign _T_26439 = valid_22_2 ? 6'h2 : _T_26438; // @[Mux.scala 31:69:@7346.4]
  assign _T_26440 = valid_22_1 ? 6'h1 : _T_26439; // @[Mux.scala 31:69:@7347.4]
  assign select_22 = valid_22_0 ? 6'h0 : _T_26440; // @[Mux.scala 31:69:@7348.4]
  assign _GEN_1409 = 6'h1 == select_22 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1410 = 6'h2 == select_22 ? io_inData_2 : _GEN_1409; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1411 = 6'h3 == select_22 ? io_inData_3 : _GEN_1410; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1412 = 6'h4 == select_22 ? io_inData_4 : _GEN_1411; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1413 = 6'h5 == select_22 ? io_inData_5 : _GEN_1412; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1414 = 6'h6 == select_22 ? io_inData_6 : _GEN_1413; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1415 = 6'h7 == select_22 ? io_inData_7 : _GEN_1414; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1416 = 6'h8 == select_22 ? io_inData_8 : _GEN_1415; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1417 = 6'h9 == select_22 ? io_inData_9 : _GEN_1416; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1418 = 6'ha == select_22 ? io_inData_10 : _GEN_1417; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1419 = 6'hb == select_22 ? io_inData_11 : _GEN_1418; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1420 = 6'hc == select_22 ? io_inData_12 : _GEN_1419; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1421 = 6'hd == select_22 ? io_inData_13 : _GEN_1420; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1422 = 6'he == select_22 ? io_inData_14 : _GEN_1421; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1423 = 6'hf == select_22 ? io_inData_15 : _GEN_1422; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1424 = 6'h10 == select_22 ? io_inData_16 : _GEN_1423; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1425 = 6'h11 == select_22 ? io_inData_17 : _GEN_1424; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1426 = 6'h12 == select_22 ? io_inData_18 : _GEN_1425; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1427 = 6'h13 == select_22 ? io_inData_19 : _GEN_1426; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1428 = 6'h14 == select_22 ? io_inData_20 : _GEN_1427; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1429 = 6'h15 == select_22 ? io_inData_21 : _GEN_1428; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1430 = 6'h16 == select_22 ? io_inData_22 : _GEN_1429; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1431 = 6'h17 == select_22 ? io_inData_23 : _GEN_1430; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1432 = 6'h18 == select_22 ? io_inData_24 : _GEN_1431; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1433 = 6'h19 == select_22 ? io_inData_25 : _GEN_1432; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1434 = 6'h1a == select_22 ? io_inData_26 : _GEN_1433; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1435 = 6'h1b == select_22 ? io_inData_27 : _GEN_1434; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1436 = 6'h1c == select_22 ? io_inData_28 : _GEN_1435; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1437 = 6'h1d == select_22 ? io_inData_29 : _GEN_1436; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1438 = 6'h1e == select_22 ? io_inData_30 : _GEN_1437; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1439 = 6'h1f == select_22 ? io_inData_31 : _GEN_1438; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1440 = 6'h20 == select_22 ? io_inData_32 : _GEN_1439; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1441 = 6'h21 == select_22 ? io_inData_33 : _GEN_1440; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1442 = 6'h22 == select_22 ? io_inData_34 : _GEN_1441; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1443 = 6'h23 == select_22 ? io_inData_35 : _GEN_1442; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1444 = 6'h24 == select_22 ? io_inData_36 : _GEN_1443; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1445 = 6'h25 == select_22 ? io_inData_37 : _GEN_1444; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1446 = 6'h26 == select_22 ? io_inData_38 : _GEN_1445; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1447 = 6'h27 == select_22 ? io_inData_39 : _GEN_1446; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1448 = 6'h28 == select_22 ? io_inData_40 : _GEN_1447; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1449 = 6'h29 == select_22 ? io_inData_41 : _GEN_1448; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1450 = 6'h2a == select_22 ? io_inData_42 : _GEN_1449; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1451 = 6'h2b == select_22 ? io_inData_43 : _GEN_1450; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1452 = 6'h2c == select_22 ? io_inData_44 : _GEN_1451; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1453 = 6'h2d == select_22 ? io_inData_45 : _GEN_1452; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1454 = 6'h2e == select_22 ? io_inData_46 : _GEN_1453; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1455 = 6'h2f == select_22 ? io_inData_47 : _GEN_1454; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1456 = 6'h30 == select_22 ? io_inData_48 : _GEN_1455; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1457 = 6'h31 == select_22 ? io_inData_49 : _GEN_1456; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1458 = 6'h32 == select_22 ? io_inData_50 : _GEN_1457; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1459 = 6'h33 == select_22 ? io_inData_51 : _GEN_1458; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1460 = 6'h34 == select_22 ? io_inData_52 : _GEN_1459; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1461 = 6'h35 == select_22 ? io_inData_53 : _GEN_1460; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1462 = 6'h36 == select_22 ? io_inData_54 : _GEN_1461; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1463 = 6'h37 == select_22 ? io_inData_55 : _GEN_1462; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1464 = 6'h38 == select_22 ? io_inData_56 : _GEN_1463; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1465 = 6'h39 == select_22 ? io_inData_57 : _GEN_1464; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1466 = 6'h3a == select_22 ? io_inData_58 : _GEN_1465; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1467 = 6'h3b == select_22 ? io_inData_59 : _GEN_1466; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1468 = 6'h3c == select_22 ? io_inData_60 : _GEN_1467; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1469 = 6'h3d == select_22 ? io_inData_61 : _GEN_1468; // @[Switch.scala 33:19:@7350.4]
  assign _GEN_1470 = 6'h3e == select_22 ? io_inData_62 : _GEN_1469; // @[Switch.scala 33:19:@7350.4]
  assign _T_26449 = {valid_22_7,valid_22_6,valid_22_5,valid_22_4,valid_22_3,valid_22_2,valid_22_1,valid_22_0}; // @[Switch.scala 34:32:@7357.4]
  assign _T_26457 = {valid_22_15,valid_22_14,valid_22_13,valid_22_12,valid_22_11,valid_22_10,valid_22_9,valid_22_8,_T_26449}; // @[Switch.scala 34:32:@7365.4]
  assign _T_26464 = {valid_22_23,valid_22_22,valid_22_21,valid_22_20,valid_22_19,valid_22_18,valid_22_17,valid_22_16}; // @[Switch.scala 34:32:@7372.4]
  assign _T_26473 = {valid_22_31,valid_22_30,valid_22_29,valid_22_28,valid_22_27,valid_22_26,valid_22_25,valid_22_24,_T_26464,_T_26457}; // @[Switch.scala 34:32:@7381.4]
  assign _T_26480 = {valid_22_39,valid_22_38,valid_22_37,valid_22_36,valid_22_35,valid_22_34,valid_22_33,valid_22_32}; // @[Switch.scala 34:32:@7388.4]
  assign _T_26488 = {valid_22_47,valid_22_46,valid_22_45,valid_22_44,valid_22_43,valid_22_42,valid_22_41,valid_22_40,_T_26480}; // @[Switch.scala 34:32:@7396.4]
  assign _T_26495 = {valid_22_55,valid_22_54,valid_22_53,valid_22_52,valid_22_51,valid_22_50,valid_22_49,valid_22_48}; // @[Switch.scala 34:32:@7403.4]
  assign _T_26504 = {valid_22_63,valid_22_62,valid_22_61,valid_22_60,valid_22_59,valid_22_58,valid_22_57,valid_22_56,_T_26495,_T_26488}; // @[Switch.scala 34:32:@7412.4]
  assign _T_26505 = {_T_26504,_T_26473}; // @[Switch.scala 34:32:@7413.4]
  assign _T_26509 = io_inAddr_0 == 6'h17; // @[Switch.scala 30:53:@7416.4]
  assign valid_23_0 = io_inValid_0 & _T_26509; // @[Switch.scala 30:36:@7417.4]
  assign _T_26512 = io_inAddr_1 == 6'h17; // @[Switch.scala 30:53:@7419.4]
  assign valid_23_1 = io_inValid_1 & _T_26512; // @[Switch.scala 30:36:@7420.4]
  assign _T_26515 = io_inAddr_2 == 6'h17; // @[Switch.scala 30:53:@7422.4]
  assign valid_23_2 = io_inValid_2 & _T_26515; // @[Switch.scala 30:36:@7423.4]
  assign _T_26518 = io_inAddr_3 == 6'h17; // @[Switch.scala 30:53:@7425.4]
  assign valid_23_3 = io_inValid_3 & _T_26518; // @[Switch.scala 30:36:@7426.4]
  assign _T_26521 = io_inAddr_4 == 6'h17; // @[Switch.scala 30:53:@7428.4]
  assign valid_23_4 = io_inValid_4 & _T_26521; // @[Switch.scala 30:36:@7429.4]
  assign _T_26524 = io_inAddr_5 == 6'h17; // @[Switch.scala 30:53:@7431.4]
  assign valid_23_5 = io_inValid_5 & _T_26524; // @[Switch.scala 30:36:@7432.4]
  assign _T_26527 = io_inAddr_6 == 6'h17; // @[Switch.scala 30:53:@7434.4]
  assign valid_23_6 = io_inValid_6 & _T_26527; // @[Switch.scala 30:36:@7435.4]
  assign _T_26530 = io_inAddr_7 == 6'h17; // @[Switch.scala 30:53:@7437.4]
  assign valid_23_7 = io_inValid_7 & _T_26530; // @[Switch.scala 30:36:@7438.4]
  assign _T_26533 = io_inAddr_8 == 6'h17; // @[Switch.scala 30:53:@7440.4]
  assign valid_23_8 = io_inValid_8 & _T_26533; // @[Switch.scala 30:36:@7441.4]
  assign _T_26536 = io_inAddr_9 == 6'h17; // @[Switch.scala 30:53:@7443.4]
  assign valid_23_9 = io_inValid_9 & _T_26536; // @[Switch.scala 30:36:@7444.4]
  assign _T_26539 = io_inAddr_10 == 6'h17; // @[Switch.scala 30:53:@7446.4]
  assign valid_23_10 = io_inValid_10 & _T_26539; // @[Switch.scala 30:36:@7447.4]
  assign _T_26542 = io_inAddr_11 == 6'h17; // @[Switch.scala 30:53:@7449.4]
  assign valid_23_11 = io_inValid_11 & _T_26542; // @[Switch.scala 30:36:@7450.4]
  assign _T_26545 = io_inAddr_12 == 6'h17; // @[Switch.scala 30:53:@7452.4]
  assign valid_23_12 = io_inValid_12 & _T_26545; // @[Switch.scala 30:36:@7453.4]
  assign _T_26548 = io_inAddr_13 == 6'h17; // @[Switch.scala 30:53:@7455.4]
  assign valid_23_13 = io_inValid_13 & _T_26548; // @[Switch.scala 30:36:@7456.4]
  assign _T_26551 = io_inAddr_14 == 6'h17; // @[Switch.scala 30:53:@7458.4]
  assign valid_23_14 = io_inValid_14 & _T_26551; // @[Switch.scala 30:36:@7459.4]
  assign _T_26554 = io_inAddr_15 == 6'h17; // @[Switch.scala 30:53:@7461.4]
  assign valid_23_15 = io_inValid_15 & _T_26554; // @[Switch.scala 30:36:@7462.4]
  assign _T_26557 = io_inAddr_16 == 6'h17; // @[Switch.scala 30:53:@7464.4]
  assign valid_23_16 = io_inValid_16 & _T_26557; // @[Switch.scala 30:36:@7465.4]
  assign _T_26560 = io_inAddr_17 == 6'h17; // @[Switch.scala 30:53:@7467.4]
  assign valid_23_17 = io_inValid_17 & _T_26560; // @[Switch.scala 30:36:@7468.4]
  assign _T_26563 = io_inAddr_18 == 6'h17; // @[Switch.scala 30:53:@7470.4]
  assign valid_23_18 = io_inValid_18 & _T_26563; // @[Switch.scala 30:36:@7471.4]
  assign _T_26566 = io_inAddr_19 == 6'h17; // @[Switch.scala 30:53:@7473.4]
  assign valid_23_19 = io_inValid_19 & _T_26566; // @[Switch.scala 30:36:@7474.4]
  assign _T_26569 = io_inAddr_20 == 6'h17; // @[Switch.scala 30:53:@7476.4]
  assign valid_23_20 = io_inValid_20 & _T_26569; // @[Switch.scala 30:36:@7477.4]
  assign _T_26572 = io_inAddr_21 == 6'h17; // @[Switch.scala 30:53:@7479.4]
  assign valid_23_21 = io_inValid_21 & _T_26572; // @[Switch.scala 30:36:@7480.4]
  assign _T_26575 = io_inAddr_22 == 6'h17; // @[Switch.scala 30:53:@7482.4]
  assign valid_23_22 = io_inValid_22 & _T_26575; // @[Switch.scala 30:36:@7483.4]
  assign _T_26578 = io_inAddr_23 == 6'h17; // @[Switch.scala 30:53:@7485.4]
  assign valid_23_23 = io_inValid_23 & _T_26578; // @[Switch.scala 30:36:@7486.4]
  assign _T_26581 = io_inAddr_24 == 6'h17; // @[Switch.scala 30:53:@7488.4]
  assign valid_23_24 = io_inValid_24 & _T_26581; // @[Switch.scala 30:36:@7489.4]
  assign _T_26584 = io_inAddr_25 == 6'h17; // @[Switch.scala 30:53:@7491.4]
  assign valid_23_25 = io_inValid_25 & _T_26584; // @[Switch.scala 30:36:@7492.4]
  assign _T_26587 = io_inAddr_26 == 6'h17; // @[Switch.scala 30:53:@7494.4]
  assign valid_23_26 = io_inValid_26 & _T_26587; // @[Switch.scala 30:36:@7495.4]
  assign _T_26590 = io_inAddr_27 == 6'h17; // @[Switch.scala 30:53:@7497.4]
  assign valid_23_27 = io_inValid_27 & _T_26590; // @[Switch.scala 30:36:@7498.4]
  assign _T_26593 = io_inAddr_28 == 6'h17; // @[Switch.scala 30:53:@7500.4]
  assign valid_23_28 = io_inValid_28 & _T_26593; // @[Switch.scala 30:36:@7501.4]
  assign _T_26596 = io_inAddr_29 == 6'h17; // @[Switch.scala 30:53:@7503.4]
  assign valid_23_29 = io_inValid_29 & _T_26596; // @[Switch.scala 30:36:@7504.4]
  assign _T_26599 = io_inAddr_30 == 6'h17; // @[Switch.scala 30:53:@7506.4]
  assign valid_23_30 = io_inValid_30 & _T_26599; // @[Switch.scala 30:36:@7507.4]
  assign _T_26602 = io_inAddr_31 == 6'h17; // @[Switch.scala 30:53:@7509.4]
  assign valid_23_31 = io_inValid_31 & _T_26602; // @[Switch.scala 30:36:@7510.4]
  assign _T_26605 = io_inAddr_32 == 6'h17; // @[Switch.scala 30:53:@7512.4]
  assign valid_23_32 = io_inValid_32 & _T_26605; // @[Switch.scala 30:36:@7513.4]
  assign _T_26608 = io_inAddr_33 == 6'h17; // @[Switch.scala 30:53:@7515.4]
  assign valid_23_33 = io_inValid_33 & _T_26608; // @[Switch.scala 30:36:@7516.4]
  assign _T_26611 = io_inAddr_34 == 6'h17; // @[Switch.scala 30:53:@7518.4]
  assign valid_23_34 = io_inValid_34 & _T_26611; // @[Switch.scala 30:36:@7519.4]
  assign _T_26614 = io_inAddr_35 == 6'h17; // @[Switch.scala 30:53:@7521.4]
  assign valid_23_35 = io_inValid_35 & _T_26614; // @[Switch.scala 30:36:@7522.4]
  assign _T_26617 = io_inAddr_36 == 6'h17; // @[Switch.scala 30:53:@7524.4]
  assign valid_23_36 = io_inValid_36 & _T_26617; // @[Switch.scala 30:36:@7525.4]
  assign _T_26620 = io_inAddr_37 == 6'h17; // @[Switch.scala 30:53:@7527.4]
  assign valid_23_37 = io_inValid_37 & _T_26620; // @[Switch.scala 30:36:@7528.4]
  assign _T_26623 = io_inAddr_38 == 6'h17; // @[Switch.scala 30:53:@7530.4]
  assign valid_23_38 = io_inValid_38 & _T_26623; // @[Switch.scala 30:36:@7531.4]
  assign _T_26626 = io_inAddr_39 == 6'h17; // @[Switch.scala 30:53:@7533.4]
  assign valid_23_39 = io_inValid_39 & _T_26626; // @[Switch.scala 30:36:@7534.4]
  assign _T_26629 = io_inAddr_40 == 6'h17; // @[Switch.scala 30:53:@7536.4]
  assign valid_23_40 = io_inValid_40 & _T_26629; // @[Switch.scala 30:36:@7537.4]
  assign _T_26632 = io_inAddr_41 == 6'h17; // @[Switch.scala 30:53:@7539.4]
  assign valid_23_41 = io_inValid_41 & _T_26632; // @[Switch.scala 30:36:@7540.4]
  assign _T_26635 = io_inAddr_42 == 6'h17; // @[Switch.scala 30:53:@7542.4]
  assign valid_23_42 = io_inValid_42 & _T_26635; // @[Switch.scala 30:36:@7543.4]
  assign _T_26638 = io_inAddr_43 == 6'h17; // @[Switch.scala 30:53:@7545.4]
  assign valid_23_43 = io_inValid_43 & _T_26638; // @[Switch.scala 30:36:@7546.4]
  assign _T_26641 = io_inAddr_44 == 6'h17; // @[Switch.scala 30:53:@7548.4]
  assign valid_23_44 = io_inValid_44 & _T_26641; // @[Switch.scala 30:36:@7549.4]
  assign _T_26644 = io_inAddr_45 == 6'h17; // @[Switch.scala 30:53:@7551.4]
  assign valid_23_45 = io_inValid_45 & _T_26644; // @[Switch.scala 30:36:@7552.4]
  assign _T_26647 = io_inAddr_46 == 6'h17; // @[Switch.scala 30:53:@7554.4]
  assign valid_23_46 = io_inValid_46 & _T_26647; // @[Switch.scala 30:36:@7555.4]
  assign _T_26650 = io_inAddr_47 == 6'h17; // @[Switch.scala 30:53:@7557.4]
  assign valid_23_47 = io_inValid_47 & _T_26650; // @[Switch.scala 30:36:@7558.4]
  assign _T_26653 = io_inAddr_48 == 6'h17; // @[Switch.scala 30:53:@7560.4]
  assign valid_23_48 = io_inValid_48 & _T_26653; // @[Switch.scala 30:36:@7561.4]
  assign _T_26656 = io_inAddr_49 == 6'h17; // @[Switch.scala 30:53:@7563.4]
  assign valid_23_49 = io_inValid_49 & _T_26656; // @[Switch.scala 30:36:@7564.4]
  assign _T_26659 = io_inAddr_50 == 6'h17; // @[Switch.scala 30:53:@7566.4]
  assign valid_23_50 = io_inValid_50 & _T_26659; // @[Switch.scala 30:36:@7567.4]
  assign _T_26662 = io_inAddr_51 == 6'h17; // @[Switch.scala 30:53:@7569.4]
  assign valid_23_51 = io_inValid_51 & _T_26662; // @[Switch.scala 30:36:@7570.4]
  assign _T_26665 = io_inAddr_52 == 6'h17; // @[Switch.scala 30:53:@7572.4]
  assign valid_23_52 = io_inValid_52 & _T_26665; // @[Switch.scala 30:36:@7573.4]
  assign _T_26668 = io_inAddr_53 == 6'h17; // @[Switch.scala 30:53:@7575.4]
  assign valid_23_53 = io_inValid_53 & _T_26668; // @[Switch.scala 30:36:@7576.4]
  assign _T_26671 = io_inAddr_54 == 6'h17; // @[Switch.scala 30:53:@7578.4]
  assign valid_23_54 = io_inValid_54 & _T_26671; // @[Switch.scala 30:36:@7579.4]
  assign _T_26674 = io_inAddr_55 == 6'h17; // @[Switch.scala 30:53:@7581.4]
  assign valid_23_55 = io_inValid_55 & _T_26674; // @[Switch.scala 30:36:@7582.4]
  assign _T_26677 = io_inAddr_56 == 6'h17; // @[Switch.scala 30:53:@7584.4]
  assign valid_23_56 = io_inValid_56 & _T_26677; // @[Switch.scala 30:36:@7585.4]
  assign _T_26680 = io_inAddr_57 == 6'h17; // @[Switch.scala 30:53:@7587.4]
  assign valid_23_57 = io_inValid_57 & _T_26680; // @[Switch.scala 30:36:@7588.4]
  assign _T_26683 = io_inAddr_58 == 6'h17; // @[Switch.scala 30:53:@7590.4]
  assign valid_23_58 = io_inValid_58 & _T_26683; // @[Switch.scala 30:36:@7591.4]
  assign _T_26686 = io_inAddr_59 == 6'h17; // @[Switch.scala 30:53:@7593.4]
  assign valid_23_59 = io_inValid_59 & _T_26686; // @[Switch.scala 30:36:@7594.4]
  assign _T_26689 = io_inAddr_60 == 6'h17; // @[Switch.scala 30:53:@7596.4]
  assign valid_23_60 = io_inValid_60 & _T_26689; // @[Switch.scala 30:36:@7597.4]
  assign _T_26692 = io_inAddr_61 == 6'h17; // @[Switch.scala 30:53:@7599.4]
  assign valid_23_61 = io_inValid_61 & _T_26692; // @[Switch.scala 30:36:@7600.4]
  assign _T_26695 = io_inAddr_62 == 6'h17; // @[Switch.scala 30:53:@7602.4]
  assign valid_23_62 = io_inValid_62 & _T_26695; // @[Switch.scala 30:36:@7603.4]
  assign _T_26698 = io_inAddr_63 == 6'h17; // @[Switch.scala 30:53:@7605.4]
  assign valid_23_63 = io_inValid_63 & _T_26698; // @[Switch.scala 30:36:@7606.4]
  assign _T_26764 = valid_23_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@7608.4]
  assign _T_26765 = valid_23_61 ? 6'h3d : _T_26764; // @[Mux.scala 31:69:@7609.4]
  assign _T_26766 = valid_23_60 ? 6'h3c : _T_26765; // @[Mux.scala 31:69:@7610.4]
  assign _T_26767 = valid_23_59 ? 6'h3b : _T_26766; // @[Mux.scala 31:69:@7611.4]
  assign _T_26768 = valid_23_58 ? 6'h3a : _T_26767; // @[Mux.scala 31:69:@7612.4]
  assign _T_26769 = valid_23_57 ? 6'h39 : _T_26768; // @[Mux.scala 31:69:@7613.4]
  assign _T_26770 = valid_23_56 ? 6'h38 : _T_26769; // @[Mux.scala 31:69:@7614.4]
  assign _T_26771 = valid_23_55 ? 6'h37 : _T_26770; // @[Mux.scala 31:69:@7615.4]
  assign _T_26772 = valid_23_54 ? 6'h36 : _T_26771; // @[Mux.scala 31:69:@7616.4]
  assign _T_26773 = valid_23_53 ? 6'h35 : _T_26772; // @[Mux.scala 31:69:@7617.4]
  assign _T_26774 = valid_23_52 ? 6'h34 : _T_26773; // @[Mux.scala 31:69:@7618.4]
  assign _T_26775 = valid_23_51 ? 6'h33 : _T_26774; // @[Mux.scala 31:69:@7619.4]
  assign _T_26776 = valid_23_50 ? 6'h32 : _T_26775; // @[Mux.scala 31:69:@7620.4]
  assign _T_26777 = valid_23_49 ? 6'h31 : _T_26776; // @[Mux.scala 31:69:@7621.4]
  assign _T_26778 = valid_23_48 ? 6'h30 : _T_26777; // @[Mux.scala 31:69:@7622.4]
  assign _T_26779 = valid_23_47 ? 6'h2f : _T_26778; // @[Mux.scala 31:69:@7623.4]
  assign _T_26780 = valid_23_46 ? 6'h2e : _T_26779; // @[Mux.scala 31:69:@7624.4]
  assign _T_26781 = valid_23_45 ? 6'h2d : _T_26780; // @[Mux.scala 31:69:@7625.4]
  assign _T_26782 = valid_23_44 ? 6'h2c : _T_26781; // @[Mux.scala 31:69:@7626.4]
  assign _T_26783 = valid_23_43 ? 6'h2b : _T_26782; // @[Mux.scala 31:69:@7627.4]
  assign _T_26784 = valid_23_42 ? 6'h2a : _T_26783; // @[Mux.scala 31:69:@7628.4]
  assign _T_26785 = valid_23_41 ? 6'h29 : _T_26784; // @[Mux.scala 31:69:@7629.4]
  assign _T_26786 = valid_23_40 ? 6'h28 : _T_26785; // @[Mux.scala 31:69:@7630.4]
  assign _T_26787 = valid_23_39 ? 6'h27 : _T_26786; // @[Mux.scala 31:69:@7631.4]
  assign _T_26788 = valid_23_38 ? 6'h26 : _T_26787; // @[Mux.scala 31:69:@7632.4]
  assign _T_26789 = valid_23_37 ? 6'h25 : _T_26788; // @[Mux.scala 31:69:@7633.4]
  assign _T_26790 = valid_23_36 ? 6'h24 : _T_26789; // @[Mux.scala 31:69:@7634.4]
  assign _T_26791 = valid_23_35 ? 6'h23 : _T_26790; // @[Mux.scala 31:69:@7635.4]
  assign _T_26792 = valid_23_34 ? 6'h22 : _T_26791; // @[Mux.scala 31:69:@7636.4]
  assign _T_26793 = valid_23_33 ? 6'h21 : _T_26792; // @[Mux.scala 31:69:@7637.4]
  assign _T_26794 = valid_23_32 ? 6'h20 : _T_26793; // @[Mux.scala 31:69:@7638.4]
  assign _T_26795 = valid_23_31 ? 6'h1f : _T_26794; // @[Mux.scala 31:69:@7639.4]
  assign _T_26796 = valid_23_30 ? 6'h1e : _T_26795; // @[Mux.scala 31:69:@7640.4]
  assign _T_26797 = valid_23_29 ? 6'h1d : _T_26796; // @[Mux.scala 31:69:@7641.4]
  assign _T_26798 = valid_23_28 ? 6'h1c : _T_26797; // @[Mux.scala 31:69:@7642.4]
  assign _T_26799 = valid_23_27 ? 6'h1b : _T_26798; // @[Mux.scala 31:69:@7643.4]
  assign _T_26800 = valid_23_26 ? 6'h1a : _T_26799; // @[Mux.scala 31:69:@7644.4]
  assign _T_26801 = valid_23_25 ? 6'h19 : _T_26800; // @[Mux.scala 31:69:@7645.4]
  assign _T_26802 = valid_23_24 ? 6'h18 : _T_26801; // @[Mux.scala 31:69:@7646.4]
  assign _T_26803 = valid_23_23 ? 6'h17 : _T_26802; // @[Mux.scala 31:69:@7647.4]
  assign _T_26804 = valid_23_22 ? 6'h16 : _T_26803; // @[Mux.scala 31:69:@7648.4]
  assign _T_26805 = valid_23_21 ? 6'h15 : _T_26804; // @[Mux.scala 31:69:@7649.4]
  assign _T_26806 = valid_23_20 ? 6'h14 : _T_26805; // @[Mux.scala 31:69:@7650.4]
  assign _T_26807 = valid_23_19 ? 6'h13 : _T_26806; // @[Mux.scala 31:69:@7651.4]
  assign _T_26808 = valid_23_18 ? 6'h12 : _T_26807; // @[Mux.scala 31:69:@7652.4]
  assign _T_26809 = valid_23_17 ? 6'h11 : _T_26808; // @[Mux.scala 31:69:@7653.4]
  assign _T_26810 = valid_23_16 ? 6'h10 : _T_26809; // @[Mux.scala 31:69:@7654.4]
  assign _T_26811 = valid_23_15 ? 6'hf : _T_26810; // @[Mux.scala 31:69:@7655.4]
  assign _T_26812 = valid_23_14 ? 6'he : _T_26811; // @[Mux.scala 31:69:@7656.4]
  assign _T_26813 = valid_23_13 ? 6'hd : _T_26812; // @[Mux.scala 31:69:@7657.4]
  assign _T_26814 = valid_23_12 ? 6'hc : _T_26813; // @[Mux.scala 31:69:@7658.4]
  assign _T_26815 = valid_23_11 ? 6'hb : _T_26814; // @[Mux.scala 31:69:@7659.4]
  assign _T_26816 = valid_23_10 ? 6'ha : _T_26815; // @[Mux.scala 31:69:@7660.4]
  assign _T_26817 = valid_23_9 ? 6'h9 : _T_26816; // @[Mux.scala 31:69:@7661.4]
  assign _T_26818 = valid_23_8 ? 6'h8 : _T_26817; // @[Mux.scala 31:69:@7662.4]
  assign _T_26819 = valid_23_7 ? 6'h7 : _T_26818; // @[Mux.scala 31:69:@7663.4]
  assign _T_26820 = valid_23_6 ? 6'h6 : _T_26819; // @[Mux.scala 31:69:@7664.4]
  assign _T_26821 = valid_23_5 ? 6'h5 : _T_26820; // @[Mux.scala 31:69:@7665.4]
  assign _T_26822 = valid_23_4 ? 6'h4 : _T_26821; // @[Mux.scala 31:69:@7666.4]
  assign _T_26823 = valid_23_3 ? 6'h3 : _T_26822; // @[Mux.scala 31:69:@7667.4]
  assign _T_26824 = valid_23_2 ? 6'h2 : _T_26823; // @[Mux.scala 31:69:@7668.4]
  assign _T_26825 = valid_23_1 ? 6'h1 : _T_26824; // @[Mux.scala 31:69:@7669.4]
  assign select_23 = valid_23_0 ? 6'h0 : _T_26825; // @[Mux.scala 31:69:@7670.4]
  assign _GEN_1473 = 6'h1 == select_23 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1474 = 6'h2 == select_23 ? io_inData_2 : _GEN_1473; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1475 = 6'h3 == select_23 ? io_inData_3 : _GEN_1474; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1476 = 6'h4 == select_23 ? io_inData_4 : _GEN_1475; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1477 = 6'h5 == select_23 ? io_inData_5 : _GEN_1476; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1478 = 6'h6 == select_23 ? io_inData_6 : _GEN_1477; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1479 = 6'h7 == select_23 ? io_inData_7 : _GEN_1478; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1480 = 6'h8 == select_23 ? io_inData_8 : _GEN_1479; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1481 = 6'h9 == select_23 ? io_inData_9 : _GEN_1480; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1482 = 6'ha == select_23 ? io_inData_10 : _GEN_1481; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1483 = 6'hb == select_23 ? io_inData_11 : _GEN_1482; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1484 = 6'hc == select_23 ? io_inData_12 : _GEN_1483; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1485 = 6'hd == select_23 ? io_inData_13 : _GEN_1484; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1486 = 6'he == select_23 ? io_inData_14 : _GEN_1485; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1487 = 6'hf == select_23 ? io_inData_15 : _GEN_1486; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1488 = 6'h10 == select_23 ? io_inData_16 : _GEN_1487; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1489 = 6'h11 == select_23 ? io_inData_17 : _GEN_1488; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1490 = 6'h12 == select_23 ? io_inData_18 : _GEN_1489; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1491 = 6'h13 == select_23 ? io_inData_19 : _GEN_1490; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1492 = 6'h14 == select_23 ? io_inData_20 : _GEN_1491; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1493 = 6'h15 == select_23 ? io_inData_21 : _GEN_1492; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1494 = 6'h16 == select_23 ? io_inData_22 : _GEN_1493; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1495 = 6'h17 == select_23 ? io_inData_23 : _GEN_1494; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1496 = 6'h18 == select_23 ? io_inData_24 : _GEN_1495; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1497 = 6'h19 == select_23 ? io_inData_25 : _GEN_1496; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1498 = 6'h1a == select_23 ? io_inData_26 : _GEN_1497; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1499 = 6'h1b == select_23 ? io_inData_27 : _GEN_1498; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1500 = 6'h1c == select_23 ? io_inData_28 : _GEN_1499; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1501 = 6'h1d == select_23 ? io_inData_29 : _GEN_1500; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1502 = 6'h1e == select_23 ? io_inData_30 : _GEN_1501; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1503 = 6'h1f == select_23 ? io_inData_31 : _GEN_1502; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1504 = 6'h20 == select_23 ? io_inData_32 : _GEN_1503; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1505 = 6'h21 == select_23 ? io_inData_33 : _GEN_1504; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1506 = 6'h22 == select_23 ? io_inData_34 : _GEN_1505; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1507 = 6'h23 == select_23 ? io_inData_35 : _GEN_1506; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1508 = 6'h24 == select_23 ? io_inData_36 : _GEN_1507; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1509 = 6'h25 == select_23 ? io_inData_37 : _GEN_1508; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1510 = 6'h26 == select_23 ? io_inData_38 : _GEN_1509; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1511 = 6'h27 == select_23 ? io_inData_39 : _GEN_1510; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1512 = 6'h28 == select_23 ? io_inData_40 : _GEN_1511; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1513 = 6'h29 == select_23 ? io_inData_41 : _GEN_1512; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1514 = 6'h2a == select_23 ? io_inData_42 : _GEN_1513; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1515 = 6'h2b == select_23 ? io_inData_43 : _GEN_1514; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1516 = 6'h2c == select_23 ? io_inData_44 : _GEN_1515; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1517 = 6'h2d == select_23 ? io_inData_45 : _GEN_1516; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1518 = 6'h2e == select_23 ? io_inData_46 : _GEN_1517; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1519 = 6'h2f == select_23 ? io_inData_47 : _GEN_1518; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1520 = 6'h30 == select_23 ? io_inData_48 : _GEN_1519; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1521 = 6'h31 == select_23 ? io_inData_49 : _GEN_1520; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1522 = 6'h32 == select_23 ? io_inData_50 : _GEN_1521; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1523 = 6'h33 == select_23 ? io_inData_51 : _GEN_1522; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1524 = 6'h34 == select_23 ? io_inData_52 : _GEN_1523; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1525 = 6'h35 == select_23 ? io_inData_53 : _GEN_1524; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1526 = 6'h36 == select_23 ? io_inData_54 : _GEN_1525; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1527 = 6'h37 == select_23 ? io_inData_55 : _GEN_1526; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1528 = 6'h38 == select_23 ? io_inData_56 : _GEN_1527; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1529 = 6'h39 == select_23 ? io_inData_57 : _GEN_1528; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1530 = 6'h3a == select_23 ? io_inData_58 : _GEN_1529; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1531 = 6'h3b == select_23 ? io_inData_59 : _GEN_1530; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1532 = 6'h3c == select_23 ? io_inData_60 : _GEN_1531; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1533 = 6'h3d == select_23 ? io_inData_61 : _GEN_1532; // @[Switch.scala 33:19:@7672.4]
  assign _GEN_1534 = 6'h3e == select_23 ? io_inData_62 : _GEN_1533; // @[Switch.scala 33:19:@7672.4]
  assign _T_26834 = {valid_23_7,valid_23_6,valid_23_5,valid_23_4,valid_23_3,valid_23_2,valid_23_1,valid_23_0}; // @[Switch.scala 34:32:@7679.4]
  assign _T_26842 = {valid_23_15,valid_23_14,valid_23_13,valid_23_12,valid_23_11,valid_23_10,valid_23_9,valid_23_8,_T_26834}; // @[Switch.scala 34:32:@7687.4]
  assign _T_26849 = {valid_23_23,valid_23_22,valid_23_21,valid_23_20,valid_23_19,valid_23_18,valid_23_17,valid_23_16}; // @[Switch.scala 34:32:@7694.4]
  assign _T_26858 = {valid_23_31,valid_23_30,valid_23_29,valid_23_28,valid_23_27,valid_23_26,valid_23_25,valid_23_24,_T_26849,_T_26842}; // @[Switch.scala 34:32:@7703.4]
  assign _T_26865 = {valid_23_39,valid_23_38,valid_23_37,valid_23_36,valid_23_35,valid_23_34,valid_23_33,valid_23_32}; // @[Switch.scala 34:32:@7710.4]
  assign _T_26873 = {valid_23_47,valid_23_46,valid_23_45,valid_23_44,valid_23_43,valid_23_42,valid_23_41,valid_23_40,_T_26865}; // @[Switch.scala 34:32:@7718.4]
  assign _T_26880 = {valid_23_55,valid_23_54,valid_23_53,valid_23_52,valid_23_51,valid_23_50,valid_23_49,valid_23_48}; // @[Switch.scala 34:32:@7725.4]
  assign _T_26889 = {valid_23_63,valid_23_62,valid_23_61,valid_23_60,valid_23_59,valid_23_58,valid_23_57,valid_23_56,_T_26880,_T_26873}; // @[Switch.scala 34:32:@7734.4]
  assign _T_26890 = {_T_26889,_T_26858}; // @[Switch.scala 34:32:@7735.4]
  assign _T_26894 = io_inAddr_0 == 6'h18; // @[Switch.scala 30:53:@7738.4]
  assign valid_24_0 = io_inValid_0 & _T_26894; // @[Switch.scala 30:36:@7739.4]
  assign _T_26897 = io_inAddr_1 == 6'h18; // @[Switch.scala 30:53:@7741.4]
  assign valid_24_1 = io_inValid_1 & _T_26897; // @[Switch.scala 30:36:@7742.4]
  assign _T_26900 = io_inAddr_2 == 6'h18; // @[Switch.scala 30:53:@7744.4]
  assign valid_24_2 = io_inValid_2 & _T_26900; // @[Switch.scala 30:36:@7745.4]
  assign _T_26903 = io_inAddr_3 == 6'h18; // @[Switch.scala 30:53:@7747.4]
  assign valid_24_3 = io_inValid_3 & _T_26903; // @[Switch.scala 30:36:@7748.4]
  assign _T_26906 = io_inAddr_4 == 6'h18; // @[Switch.scala 30:53:@7750.4]
  assign valid_24_4 = io_inValid_4 & _T_26906; // @[Switch.scala 30:36:@7751.4]
  assign _T_26909 = io_inAddr_5 == 6'h18; // @[Switch.scala 30:53:@7753.4]
  assign valid_24_5 = io_inValid_5 & _T_26909; // @[Switch.scala 30:36:@7754.4]
  assign _T_26912 = io_inAddr_6 == 6'h18; // @[Switch.scala 30:53:@7756.4]
  assign valid_24_6 = io_inValid_6 & _T_26912; // @[Switch.scala 30:36:@7757.4]
  assign _T_26915 = io_inAddr_7 == 6'h18; // @[Switch.scala 30:53:@7759.4]
  assign valid_24_7 = io_inValid_7 & _T_26915; // @[Switch.scala 30:36:@7760.4]
  assign _T_26918 = io_inAddr_8 == 6'h18; // @[Switch.scala 30:53:@7762.4]
  assign valid_24_8 = io_inValid_8 & _T_26918; // @[Switch.scala 30:36:@7763.4]
  assign _T_26921 = io_inAddr_9 == 6'h18; // @[Switch.scala 30:53:@7765.4]
  assign valid_24_9 = io_inValid_9 & _T_26921; // @[Switch.scala 30:36:@7766.4]
  assign _T_26924 = io_inAddr_10 == 6'h18; // @[Switch.scala 30:53:@7768.4]
  assign valid_24_10 = io_inValid_10 & _T_26924; // @[Switch.scala 30:36:@7769.4]
  assign _T_26927 = io_inAddr_11 == 6'h18; // @[Switch.scala 30:53:@7771.4]
  assign valid_24_11 = io_inValid_11 & _T_26927; // @[Switch.scala 30:36:@7772.4]
  assign _T_26930 = io_inAddr_12 == 6'h18; // @[Switch.scala 30:53:@7774.4]
  assign valid_24_12 = io_inValid_12 & _T_26930; // @[Switch.scala 30:36:@7775.4]
  assign _T_26933 = io_inAddr_13 == 6'h18; // @[Switch.scala 30:53:@7777.4]
  assign valid_24_13 = io_inValid_13 & _T_26933; // @[Switch.scala 30:36:@7778.4]
  assign _T_26936 = io_inAddr_14 == 6'h18; // @[Switch.scala 30:53:@7780.4]
  assign valid_24_14 = io_inValid_14 & _T_26936; // @[Switch.scala 30:36:@7781.4]
  assign _T_26939 = io_inAddr_15 == 6'h18; // @[Switch.scala 30:53:@7783.4]
  assign valid_24_15 = io_inValid_15 & _T_26939; // @[Switch.scala 30:36:@7784.4]
  assign _T_26942 = io_inAddr_16 == 6'h18; // @[Switch.scala 30:53:@7786.4]
  assign valid_24_16 = io_inValid_16 & _T_26942; // @[Switch.scala 30:36:@7787.4]
  assign _T_26945 = io_inAddr_17 == 6'h18; // @[Switch.scala 30:53:@7789.4]
  assign valid_24_17 = io_inValid_17 & _T_26945; // @[Switch.scala 30:36:@7790.4]
  assign _T_26948 = io_inAddr_18 == 6'h18; // @[Switch.scala 30:53:@7792.4]
  assign valid_24_18 = io_inValid_18 & _T_26948; // @[Switch.scala 30:36:@7793.4]
  assign _T_26951 = io_inAddr_19 == 6'h18; // @[Switch.scala 30:53:@7795.4]
  assign valid_24_19 = io_inValid_19 & _T_26951; // @[Switch.scala 30:36:@7796.4]
  assign _T_26954 = io_inAddr_20 == 6'h18; // @[Switch.scala 30:53:@7798.4]
  assign valid_24_20 = io_inValid_20 & _T_26954; // @[Switch.scala 30:36:@7799.4]
  assign _T_26957 = io_inAddr_21 == 6'h18; // @[Switch.scala 30:53:@7801.4]
  assign valid_24_21 = io_inValid_21 & _T_26957; // @[Switch.scala 30:36:@7802.4]
  assign _T_26960 = io_inAddr_22 == 6'h18; // @[Switch.scala 30:53:@7804.4]
  assign valid_24_22 = io_inValid_22 & _T_26960; // @[Switch.scala 30:36:@7805.4]
  assign _T_26963 = io_inAddr_23 == 6'h18; // @[Switch.scala 30:53:@7807.4]
  assign valid_24_23 = io_inValid_23 & _T_26963; // @[Switch.scala 30:36:@7808.4]
  assign _T_26966 = io_inAddr_24 == 6'h18; // @[Switch.scala 30:53:@7810.4]
  assign valid_24_24 = io_inValid_24 & _T_26966; // @[Switch.scala 30:36:@7811.4]
  assign _T_26969 = io_inAddr_25 == 6'h18; // @[Switch.scala 30:53:@7813.4]
  assign valid_24_25 = io_inValid_25 & _T_26969; // @[Switch.scala 30:36:@7814.4]
  assign _T_26972 = io_inAddr_26 == 6'h18; // @[Switch.scala 30:53:@7816.4]
  assign valid_24_26 = io_inValid_26 & _T_26972; // @[Switch.scala 30:36:@7817.4]
  assign _T_26975 = io_inAddr_27 == 6'h18; // @[Switch.scala 30:53:@7819.4]
  assign valid_24_27 = io_inValid_27 & _T_26975; // @[Switch.scala 30:36:@7820.4]
  assign _T_26978 = io_inAddr_28 == 6'h18; // @[Switch.scala 30:53:@7822.4]
  assign valid_24_28 = io_inValid_28 & _T_26978; // @[Switch.scala 30:36:@7823.4]
  assign _T_26981 = io_inAddr_29 == 6'h18; // @[Switch.scala 30:53:@7825.4]
  assign valid_24_29 = io_inValid_29 & _T_26981; // @[Switch.scala 30:36:@7826.4]
  assign _T_26984 = io_inAddr_30 == 6'h18; // @[Switch.scala 30:53:@7828.4]
  assign valid_24_30 = io_inValid_30 & _T_26984; // @[Switch.scala 30:36:@7829.4]
  assign _T_26987 = io_inAddr_31 == 6'h18; // @[Switch.scala 30:53:@7831.4]
  assign valid_24_31 = io_inValid_31 & _T_26987; // @[Switch.scala 30:36:@7832.4]
  assign _T_26990 = io_inAddr_32 == 6'h18; // @[Switch.scala 30:53:@7834.4]
  assign valid_24_32 = io_inValid_32 & _T_26990; // @[Switch.scala 30:36:@7835.4]
  assign _T_26993 = io_inAddr_33 == 6'h18; // @[Switch.scala 30:53:@7837.4]
  assign valid_24_33 = io_inValid_33 & _T_26993; // @[Switch.scala 30:36:@7838.4]
  assign _T_26996 = io_inAddr_34 == 6'h18; // @[Switch.scala 30:53:@7840.4]
  assign valid_24_34 = io_inValid_34 & _T_26996; // @[Switch.scala 30:36:@7841.4]
  assign _T_26999 = io_inAddr_35 == 6'h18; // @[Switch.scala 30:53:@7843.4]
  assign valid_24_35 = io_inValid_35 & _T_26999; // @[Switch.scala 30:36:@7844.4]
  assign _T_27002 = io_inAddr_36 == 6'h18; // @[Switch.scala 30:53:@7846.4]
  assign valid_24_36 = io_inValid_36 & _T_27002; // @[Switch.scala 30:36:@7847.4]
  assign _T_27005 = io_inAddr_37 == 6'h18; // @[Switch.scala 30:53:@7849.4]
  assign valid_24_37 = io_inValid_37 & _T_27005; // @[Switch.scala 30:36:@7850.4]
  assign _T_27008 = io_inAddr_38 == 6'h18; // @[Switch.scala 30:53:@7852.4]
  assign valid_24_38 = io_inValid_38 & _T_27008; // @[Switch.scala 30:36:@7853.4]
  assign _T_27011 = io_inAddr_39 == 6'h18; // @[Switch.scala 30:53:@7855.4]
  assign valid_24_39 = io_inValid_39 & _T_27011; // @[Switch.scala 30:36:@7856.4]
  assign _T_27014 = io_inAddr_40 == 6'h18; // @[Switch.scala 30:53:@7858.4]
  assign valid_24_40 = io_inValid_40 & _T_27014; // @[Switch.scala 30:36:@7859.4]
  assign _T_27017 = io_inAddr_41 == 6'h18; // @[Switch.scala 30:53:@7861.4]
  assign valid_24_41 = io_inValid_41 & _T_27017; // @[Switch.scala 30:36:@7862.4]
  assign _T_27020 = io_inAddr_42 == 6'h18; // @[Switch.scala 30:53:@7864.4]
  assign valid_24_42 = io_inValid_42 & _T_27020; // @[Switch.scala 30:36:@7865.4]
  assign _T_27023 = io_inAddr_43 == 6'h18; // @[Switch.scala 30:53:@7867.4]
  assign valid_24_43 = io_inValid_43 & _T_27023; // @[Switch.scala 30:36:@7868.4]
  assign _T_27026 = io_inAddr_44 == 6'h18; // @[Switch.scala 30:53:@7870.4]
  assign valid_24_44 = io_inValid_44 & _T_27026; // @[Switch.scala 30:36:@7871.4]
  assign _T_27029 = io_inAddr_45 == 6'h18; // @[Switch.scala 30:53:@7873.4]
  assign valid_24_45 = io_inValid_45 & _T_27029; // @[Switch.scala 30:36:@7874.4]
  assign _T_27032 = io_inAddr_46 == 6'h18; // @[Switch.scala 30:53:@7876.4]
  assign valid_24_46 = io_inValid_46 & _T_27032; // @[Switch.scala 30:36:@7877.4]
  assign _T_27035 = io_inAddr_47 == 6'h18; // @[Switch.scala 30:53:@7879.4]
  assign valid_24_47 = io_inValid_47 & _T_27035; // @[Switch.scala 30:36:@7880.4]
  assign _T_27038 = io_inAddr_48 == 6'h18; // @[Switch.scala 30:53:@7882.4]
  assign valid_24_48 = io_inValid_48 & _T_27038; // @[Switch.scala 30:36:@7883.4]
  assign _T_27041 = io_inAddr_49 == 6'h18; // @[Switch.scala 30:53:@7885.4]
  assign valid_24_49 = io_inValid_49 & _T_27041; // @[Switch.scala 30:36:@7886.4]
  assign _T_27044 = io_inAddr_50 == 6'h18; // @[Switch.scala 30:53:@7888.4]
  assign valid_24_50 = io_inValid_50 & _T_27044; // @[Switch.scala 30:36:@7889.4]
  assign _T_27047 = io_inAddr_51 == 6'h18; // @[Switch.scala 30:53:@7891.4]
  assign valid_24_51 = io_inValid_51 & _T_27047; // @[Switch.scala 30:36:@7892.4]
  assign _T_27050 = io_inAddr_52 == 6'h18; // @[Switch.scala 30:53:@7894.4]
  assign valid_24_52 = io_inValid_52 & _T_27050; // @[Switch.scala 30:36:@7895.4]
  assign _T_27053 = io_inAddr_53 == 6'h18; // @[Switch.scala 30:53:@7897.4]
  assign valid_24_53 = io_inValid_53 & _T_27053; // @[Switch.scala 30:36:@7898.4]
  assign _T_27056 = io_inAddr_54 == 6'h18; // @[Switch.scala 30:53:@7900.4]
  assign valid_24_54 = io_inValid_54 & _T_27056; // @[Switch.scala 30:36:@7901.4]
  assign _T_27059 = io_inAddr_55 == 6'h18; // @[Switch.scala 30:53:@7903.4]
  assign valid_24_55 = io_inValid_55 & _T_27059; // @[Switch.scala 30:36:@7904.4]
  assign _T_27062 = io_inAddr_56 == 6'h18; // @[Switch.scala 30:53:@7906.4]
  assign valid_24_56 = io_inValid_56 & _T_27062; // @[Switch.scala 30:36:@7907.4]
  assign _T_27065 = io_inAddr_57 == 6'h18; // @[Switch.scala 30:53:@7909.4]
  assign valid_24_57 = io_inValid_57 & _T_27065; // @[Switch.scala 30:36:@7910.4]
  assign _T_27068 = io_inAddr_58 == 6'h18; // @[Switch.scala 30:53:@7912.4]
  assign valid_24_58 = io_inValid_58 & _T_27068; // @[Switch.scala 30:36:@7913.4]
  assign _T_27071 = io_inAddr_59 == 6'h18; // @[Switch.scala 30:53:@7915.4]
  assign valid_24_59 = io_inValid_59 & _T_27071; // @[Switch.scala 30:36:@7916.4]
  assign _T_27074 = io_inAddr_60 == 6'h18; // @[Switch.scala 30:53:@7918.4]
  assign valid_24_60 = io_inValid_60 & _T_27074; // @[Switch.scala 30:36:@7919.4]
  assign _T_27077 = io_inAddr_61 == 6'h18; // @[Switch.scala 30:53:@7921.4]
  assign valid_24_61 = io_inValid_61 & _T_27077; // @[Switch.scala 30:36:@7922.4]
  assign _T_27080 = io_inAddr_62 == 6'h18; // @[Switch.scala 30:53:@7924.4]
  assign valid_24_62 = io_inValid_62 & _T_27080; // @[Switch.scala 30:36:@7925.4]
  assign _T_27083 = io_inAddr_63 == 6'h18; // @[Switch.scala 30:53:@7927.4]
  assign valid_24_63 = io_inValid_63 & _T_27083; // @[Switch.scala 30:36:@7928.4]
  assign _T_27149 = valid_24_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@7930.4]
  assign _T_27150 = valid_24_61 ? 6'h3d : _T_27149; // @[Mux.scala 31:69:@7931.4]
  assign _T_27151 = valid_24_60 ? 6'h3c : _T_27150; // @[Mux.scala 31:69:@7932.4]
  assign _T_27152 = valid_24_59 ? 6'h3b : _T_27151; // @[Mux.scala 31:69:@7933.4]
  assign _T_27153 = valid_24_58 ? 6'h3a : _T_27152; // @[Mux.scala 31:69:@7934.4]
  assign _T_27154 = valid_24_57 ? 6'h39 : _T_27153; // @[Mux.scala 31:69:@7935.4]
  assign _T_27155 = valid_24_56 ? 6'h38 : _T_27154; // @[Mux.scala 31:69:@7936.4]
  assign _T_27156 = valid_24_55 ? 6'h37 : _T_27155; // @[Mux.scala 31:69:@7937.4]
  assign _T_27157 = valid_24_54 ? 6'h36 : _T_27156; // @[Mux.scala 31:69:@7938.4]
  assign _T_27158 = valid_24_53 ? 6'h35 : _T_27157; // @[Mux.scala 31:69:@7939.4]
  assign _T_27159 = valid_24_52 ? 6'h34 : _T_27158; // @[Mux.scala 31:69:@7940.4]
  assign _T_27160 = valid_24_51 ? 6'h33 : _T_27159; // @[Mux.scala 31:69:@7941.4]
  assign _T_27161 = valid_24_50 ? 6'h32 : _T_27160; // @[Mux.scala 31:69:@7942.4]
  assign _T_27162 = valid_24_49 ? 6'h31 : _T_27161; // @[Mux.scala 31:69:@7943.4]
  assign _T_27163 = valid_24_48 ? 6'h30 : _T_27162; // @[Mux.scala 31:69:@7944.4]
  assign _T_27164 = valid_24_47 ? 6'h2f : _T_27163; // @[Mux.scala 31:69:@7945.4]
  assign _T_27165 = valid_24_46 ? 6'h2e : _T_27164; // @[Mux.scala 31:69:@7946.4]
  assign _T_27166 = valid_24_45 ? 6'h2d : _T_27165; // @[Mux.scala 31:69:@7947.4]
  assign _T_27167 = valid_24_44 ? 6'h2c : _T_27166; // @[Mux.scala 31:69:@7948.4]
  assign _T_27168 = valid_24_43 ? 6'h2b : _T_27167; // @[Mux.scala 31:69:@7949.4]
  assign _T_27169 = valid_24_42 ? 6'h2a : _T_27168; // @[Mux.scala 31:69:@7950.4]
  assign _T_27170 = valid_24_41 ? 6'h29 : _T_27169; // @[Mux.scala 31:69:@7951.4]
  assign _T_27171 = valid_24_40 ? 6'h28 : _T_27170; // @[Mux.scala 31:69:@7952.4]
  assign _T_27172 = valid_24_39 ? 6'h27 : _T_27171; // @[Mux.scala 31:69:@7953.4]
  assign _T_27173 = valid_24_38 ? 6'h26 : _T_27172; // @[Mux.scala 31:69:@7954.4]
  assign _T_27174 = valid_24_37 ? 6'h25 : _T_27173; // @[Mux.scala 31:69:@7955.4]
  assign _T_27175 = valid_24_36 ? 6'h24 : _T_27174; // @[Mux.scala 31:69:@7956.4]
  assign _T_27176 = valid_24_35 ? 6'h23 : _T_27175; // @[Mux.scala 31:69:@7957.4]
  assign _T_27177 = valid_24_34 ? 6'h22 : _T_27176; // @[Mux.scala 31:69:@7958.4]
  assign _T_27178 = valid_24_33 ? 6'h21 : _T_27177; // @[Mux.scala 31:69:@7959.4]
  assign _T_27179 = valid_24_32 ? 6'h20 : _T_27178; // @[Mux.scala 31:69:@7960.4]
  assign _T_27180 = valid_24_31 ? 6'h1f : _T_27179; // @[Mux.scala 31:69:@7961.4]
  assign _T_27181 = valid_24_30 ? 6'h1e : _T_27180; // @[Mux.scala 31:69:@7962.4]
  assign _T_27182 = valid_24_29 ? 6'h1d : _T_27181; // @[Mux.scala 31:69:@7963.4]
  assign _T_27183 = valid_24_28 ? 6'h1c : _T_27182; // @[Mux.scala 31:69:@7964.4]
  assign _T_27184 = valid_24_27 ? 6'h1b : _T_27183; // @[Mux.scala 31:69:@7965.4]
  assign _T_27185 = valid_24_26 ? 6'h1a : _T_27184; // @[Mux.scala 31:69:@7966.4]
  assign _T_27186 = valid_24_25 ? 6'h19 : _T_27185; // @[Mux.scala 31:69:@7967.4]
  assign _T_27187 = valid_24_24 ? 6'h18 : _T_27186; // @[Mux.scala 31:69:@7968.4]
  assign _T_27188 = valid_24_23 ? 6'h17 : _T_27187; // @[Mux.scala 31:69:@7969.4]
  assign _T_27189 = valid_24_22 ? 6'h16 : _T_27188; // @[Mux.scala 31:69:@7970.4]
  assign _T_27190 = valid_24_21 ? 6'h15 : _T_27189; // @[Mux.scala 31:69:@7971.4]
  assign _T_27191 = valid_24_20 ? 6'h14 : _T_27190; // @[Mux.scala 31:69:@7972.4]
  assign _T_27192 = valid_24_19 ? 6'h13 : _T_27191; // @[Mux.scala 31:69:@7973.4]
  assign _T_27193 = valid_24_18 ? 6'h12 : _T_27192; // @[Mux.scala 31:69:@7974.4]
  assign _T_27194 = valid_24_17 ? 6'h11 : _T_27193; // @[Mux.scala 31:69:@7975.4]
  assign _T_27195 = valid_24_16 ? 6'h10 : _T_27194; // @[Mux.scala 31:69:@7976.4]
  assign _T_27196 = valid_24_15 ? 6'hf : _T_27195; // @[Mux.scala 31:69:@7977.4]
  assign _T_27197 = valid_24_14 ? 6'he : _T_27196; // @[Mux.scala 31:69:@7978.4]
  assign _T_27198 = valid_24_13 ? 6'hd : _T_27197; // @[Mux.scala 31:69:@7979.4]
  assign _T_27199 = valid_24_12 ? 6'hc : _T_27198; // @[Mux.scala 31:69:@7980.4]
  assign _T_27200 = valid_24_11 ? 6'hb : _T_27199; // @[Mux.scala 31:69:@7981.4]
  assign _T_27201 = valid_24_10 ? 6'ha : _T_27200; // @[Mux.scala 31:69:@7982.4]
  assign _T_27202 = valid_24_9 ? 6'h9 : _T_27201; // @[Mux.scala 31:69:@7983.4]
  assign _T_27203 = valid_24_8 ? 6'h8 : _T_27202; // @[Mux.scala 31:69:@7984.4]
  assign _T_27204 = valid_24_7 ? 6'h7 : _T_27203; // @[Mux.scala 31:69:@7985.4]
  assign _T_27205 = valid_24_6 ? 6'h6 : _T_27204; // @[Mux.scala 31:69:@7986.4]
  assign _T_27206 = valid_24_5 ? 6'h5 : _T_27205; // @[Mux.scala 31:69:@7987.4]
  assign _T_27207 = valid_24_4 ? 6'h4 : _T_27206; // @[Mux.scala 31:69:@7988.4]
  assign _T_27208 = valid_24_3 ? 6'h3 : _T_27207; // @[Mux.scala 31:69:@7989.4]
  assign _T_27209 = valid_24_2 ? 6'h2 : _T_27208; // @[Mux.scala 31:69:@7990.4]
  assign _T_27210 = valid_24_1 ? 6'h1 : _T_27209; // @[Mux.scala 31:69:@7991.4]
  assign select_24 = valid_24_0 ? 6'h0 : _T_27210; // @[Mux.scala 31:69:@7992.4]
  assign _GEN_1537 = 6'h1 == select_24 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1538 = 6'h2 == select_24 ? io_inData_2 : _GEN_1537; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1539 = 6'h3 == select_24 ? io_inData_3 : _GEN_1538; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1540 = 6'h4 == select_24 ? io_inData_4 : _GEN_1539; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1541 = 6'h5 == select_24 ? io_inData_5 : _GEN_1540; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1542 = 6'h6 == select_24 ? io_inData_6 : _GEN_1541; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1543 = 6'h7 == select_24 ? io_inData_7 : _GEN_1542; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1544 = 6'h8 == select_24 ? io_inData_8 : _GEN_1543; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1545 = 6'h9 == select_24 ? io_inData_9 : _GEN_1544; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1546 = 6'ha == select_24 ? io_inData_10 : _GEN_1545; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1547 = 6'hb == select_24 ? io_inData_11 : _GEN_1546; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1548 = 6'hc == select_24 ? io_inData_12 : _GEN_1547; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1549 = 6'hd == select_24 ? io_inData_13 : _GEN_1548; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1550 = 6'he == select_24 ? io_inData_14 : _GEN_1549; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1551 = 6'hf == select_24 ? io_inData_15 : _GEN_1550; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1552 = 6'h10 == select_24 ? io_inData_16 : _GEN_1551; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1553 = 6'h11 == select_24 ? io_inData_17 : _GEN_1552; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1554 = 6'h12 == select_24 ? io_inData_18 : _GEN_1553; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1555 = 6'h13 == select_24 ? io_inData_19 : _GEN_1554; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1556 = 6'h14 == select_24 ? io_inData_20 : _GEN_1555; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1557 = 6'h15 == select_24 ? io_inData_21 : _GEN_1556; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1558 = 6'h16 == select_24 ? io_inData_22 : _GEN_1557; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1559 = 6'h17 == select_24 ? io_inData_23 : _GEN_1558; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1560 = 6'h18 == select_24 ? io_inData_24 : _GEN_1559; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1561 = 6'h19 == select_24 ? io_inData_25 : _GEN_1560; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1562 = 6'h1a == select_24 ? io_inData_26 : _GEN_1561; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1563 = 6'h1b == select_24 ? io_inData_27 : _GEN_1562; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1564 = 6'h1c == select_24 ? io_inData_28 : _GEN_1563; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1565 = 6'h1d == select_24 ? io_inData_29 : _GEN_1564; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1566 = 6'h1e == select_24 ? io_inData_30 : _GEN_1565; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1567 = 6'h1f == select_24 ? io_inData_31 : _GEN_1566; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1568 = 6'h20 == select_24 ? io_inData_32 : _GEN_1567; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1569 = 6'h21 == select_24 ? io_inData_33 : _GEN_1568; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1570 = 6'h22 == select_24 ? io_inData_34 : _GEN_1569; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1571 = 6'h23 == select_24 ? io_inData_35 : _GEN_1570; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1572 = 6'h24 == select_24 ? io_inData_36 : _GEN_1571; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1573 = 6'h25 == select_24 ? io_inData_37 : _GEN_1572; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1574 = 6'h26 == select_24 ? io_inData_38 : _GEN_1573; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1575 = 6'h27 == select_24 ? io_inData_39 : _GEN_1574; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1576 = 6'h28 == select_24 ? io_inData_40 : _GEN_1575; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1577 = 6'h29 == select_24 ? io_inData_41 : _GEN_1576; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1578 = 6'h2a == select_24 ? io_inData_42 : _GEN_1577; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1579 = 6'h2b == select_24 ? io_inData_43 : _GEN_1578; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1580 = 6'h2c == select_24 ? io_inData_44 : _GEN_1579; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1581 = 6'h2d == select_24 ? io_inData_45 : _GEN_1580; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1582 = 6'h2e == select_24 ? io_inData_46 : _GEN_1581; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1583 = 6'h2f == select_24 ? io_inData_47 : _GEN_1582; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1584 = 6'h30 == select_24 ? io_inData_48 : _GEN_1583; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1585 = 6'h31 == select_24 ? io_inData_49 : _GEN_1584; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1586 = 6'h32 == select_24 ? io_inData_50 : _GEN_1585; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1587 = 6'h33 == select_24 ? io_inData_51 : _GEN_1586; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1588 = 6'h34 == select_24 ? io_inData_52 : _GEN_1587; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1589 = 6'h35 == select_24 ? io_inData_53 : _GEN_1588; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1590 = 6'h36 == select_24 ? io_inData_54 : _GEN_1589; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1591 = 6'h37 == select_24 ? io_inData_55 : _GEN_1590; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1592 = 6'h38 == select_24 ? io_inData_56 : _GEN_1591; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1593 = 6'h39 == select_24 ? io_inData_57 : _GEN_1592; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1594 = 6'h3a == select_24 ? io_inData_58 : _GEN_1593; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1595 = 6'h3b == select_24 ? io_inData_59 : _GEN_1594; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1596 = 6'h3c == select_24 ? io_inData_60 : _GEN_1595; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1597 = 6'h3d == select_24 ? io_inData_61 : _GEN_1596; // @[Switch.scala 33:19:@7994.4]
  assign _GEN_1598 = 6'h3e == select_24 ? io_inData_62 : _GEN_1597; // @[Switch.scala 33:19:@7994.4]
  assign _T_27219 = {valid_24_7,valid_24_6,valid_24_5,valid_24_4,valid_24_3,valid_24_2,valid_24_1,valid_24_0}; // @[Switch.scala 34:32:@8001.4]
  assign _T_27227 = {valid_24_15,valid_24_14,valid_24_13,valid_24_12,valid_24_11,valid_24_10,valid_24_9,valid_24_8,_T_27219}; // @[Switch.scala 34:32:@8009.4]
  assign _T_27234 = {valid_24_23,valid_24_22,valid_24_21,valid_24_20,valid_24_19,valid_24_18,valid_24_17,valid_24_16}; // @[Switch.scala 34:32:@8016.4]
  assign _T_27243 = {valid_24_31,valid_24_30,valid_24_29,valid_24_28,valid_24_27,valid_24_26,valid_24_25,valid_24_24,_T_27234,_T_27227}; // @[Switch.scala 34:32:@8025.4]
  assign _T_27250 = {valid_24_39,valid_24_38,valid_24_37,valid_24_36,valid_24_35,valid_24_34,valid_24_33,valid_24_32}; // @[Switch.scala 34:32:@8032.4]
  assign _T_27258 = {valid_24_47,valid_24_46,valid_24_45,valid_24_44,valid_24_43,valid_24_42,valid_24_41,valid_24_40,_T_27250}; // @[Switch.scala 34:32:@8040.4]
  assign _T_27265 = {valid_24_55,valid_24_54,valid_24_53,valid_24_52,valid_24_51,valid_24_50,valid_24_49,valid_24_48}; // @[Switch.scala 34:32:@8047.4]
  assign _T_27274 = {valid_24_63,valid_24_62,valid_24_61,valid_24_60,valid_24_59,valid_24_58,valid_24_57,valid_24_56,_T_27265,_T_27258}; // @[Switch.scala 34:32:@8056.4]
  assign _T_27275 = {_T_27274,_T_27243}; // @[Switch.scala 34:32:@8057.4]
  assign _T_27279 = io_inAddr_0 == 6'h19; // @[Switch.scala 30:53:@8060.4]
  assign valid_25_0 = io_inValid_0 & _T_27279; // @[Switch.scala 30:36:@8061.4]
  assign _T_27282 = io_inAddr_1 == 6'h19; // @[Switch.scala 30:53:@8063.4]
  assign valid_25_1 = io_inValid_1 & _T_27282; // @[Switch.scala 30:36:@8064.4]
  assign _T_27285 = io_inAddr_2 == 6'h19; // @[Switch.scala 30:53:@8066.4]
  assign valid_25_2 = io_inValid_2 & _T_27285; // @[Switch.scala 30:36:@8067.4]
  assign _T_27288 = io_inAddr_3 == 6'h19; // @[Switch.scala 30:53:@8069.4]
  assign valid_25_3 = io_inValid_3 & _T_27288; // @[Switch.scala 30:36:@8070.4]
  assign _T_27291 = io_inAddr_4 == 6'h19; // @[Switch.scala 30:53:@8072.4]
  assign valid_25_4 = io_inValid_4 & _T_27291; // @[Switch.scala 30:36:@8073.4]
  assign _T_27294 = io_inAddr_5 == 6'h19; // @[Switch.scala 30:53:@8075.4]
  assign valid_25_5 = io_inValid_5 & _T_27294; // @[Switch.scala 30:36:@8076.4]
  assign _T_27297 = io_inAddr_6 == 6'h19; // @[Switch.scala 30:53:@8078.4]
  assign valid_25_6 = io_inValid_6 & _T_27297; // @[Switch.scala 30:36:@8079.4]
  assign _T_27300 = io_inAddr_7 == 6'h19; // @[Switch.scala 30:53:@8081.4]
  assign valid_25_7 = io_inValid_7 & _T_27300; // @[Switch.scala 30:36:@8082.4]
  assign _T_27303 = io_inAddr_8 == 6'h19; // @[Switch.scala 30:53:@8084.4]
  assign valid_25_8 = io_inValid_8 & _T_27303; // @[Switch.scala 30:36:@8085.4]
  assign _T_27306 = io_inAddr_9 == 6'h19; // @[Switch.scala 30:53:@8087.4]
  assign valid_25_9 = io_inValid_9 & _T_27306; // @[Switch.scala 30:36:@8088.4]
  assign _T_27309 = io_inAddr_10 == 6'h19; // @[Switch.scala 30:53:@8090.4]
  assign valid_25_10 = io_inValid_10 & _T_27309; // @[Switch.scala 30:36:@8091.4]
  assign _T_27312 = io_inAddr_11 == 6'h19; // @[Switch.scala 30:53:@8093.4]
  assign valid_25_11 = io_inValid_11 & _T_27312; // @[Switch.scala 30:36:@8094.4]
  assign _T_27315 = io_inAddr_12 == 6'h19; // @[Switch.scala 30:53:@8096.4]
  assign valid_25_12 = io_inValid_12 & _T_27315; // @[Switch.scala 30:36:@8097.4]
  assign _T_27318 = io_inAddr_13 == 6'h19; // @[Switch.scala 30:53:@8099.4]
  assign valid_25_13 = io_inValid_13 & _T_27318; // @[Switch.scala 30:36:@8100.4]
  assign _T_27321 = io_inAddr_14 == 6'h19; // @[Switch.scala 30:53:@8102.4]
  assign valid_25_14 = io_inValid_14 & _T_27321; // @[Switch.scala 30:36:@8103.4]
  assign _T_27324 = io_inAddr_15 == 6'h19; // @[Switch.scala 30:53:@8105.4]
  assign valid_25_15 = io_inValid_15 & _T_27324; // @[Switch.scala 30:36:@8106.4]
  assign _T_27327 = io_inAddr_16 == 6'h19; // @[Switch.scala 30:53:@8108.4]
  assign valid_25_16 = io_inValid_16 & _T_27327; // @[Switch.scala 30:36:@8109.4]
  assign _T_27330 = io_inAddr_17 == 6'h19; // @[Switch.scala 30:53:@8111.4]
  assign valid_25_17 = io_inValid_17 & _T_27330; // @[Switch.scala 30:36:@8112.4]
  assign _T_27333 = io_inAddr_18 == 6'h19; // @[Switch.scala 30:53:@8114.4]
  assign valid_25_18 = io_inValid_18 & _T_27333; // @[Switch.scala 30:36:@8115.4]
  assign _T_27336 = io_inAddr_19 == 6'h19; // @[Switch.scala 30:53:@8117.4]
  assign valid_25_19 = io_inValid_19 & _T_27336; // @[Switch.scala 30:36:@8118.4]
  assign _T_27339 = io_inAddr_20 == 6'h19; // @[Switch.scala 30:53:@8120.4]
  assign valid_25_20 = io_inValid_20 & _T_27339; // @[Switch.scala 30:36:@8121.4]
  assign _T_27342 = io_inAddr_21 == 6'h19; // @[Switch.scala 30:53:@8123.4]
  assign valid_25_21 = io_inValid_21 & _T_27342; // @[Switch.scala 30:36:@8124.4]
  assign _T_27345 = io_inAddr_22 == 6'h19; // @[Switch.scala 30:53:@8126.4]
  assign valid_25_22 = io_inValid_22 & _T_27345; // @[Switch.scala 30:36:@8127.4]
  assign _T_27348 = io_inAddr_23 == 6'h19; // @[Switch.scala 30:53:@8129.4]
  assign valid_25_23 = io_inValid_23 & _T_27348; // @[Switch.scala 30:36:@8130.4]
  assign _T_27351 = io_inAddr_24 == 6'h19; // @[Switch.scala 30:53:@8132.4]
  assign valid_25_24 = io_inValid_24 & _T_27351; // @[Switch.scala 30:36:@8133.4]
  assign _T_27354 = io_inAddr_25 == 6'h19; // @[Switch.scala 30:53:@8135.4]
  assign valid_25_25 = io_inValid_25 & _T_27354; // @[Switch.scala 30:36:@8136.4]
  assign _T_27357 = io_inAddr_26 == 6'h19; // @[Switch.scala 30:53:@8138.4]
  assign valid_25_26 = io_inValid_26 & _T_27357; // @[Switch.scala 30:36:@8139.4]
  assign _T_27360 = io_inAddr_27 == 6'h19; // @[Switch.scala 30:53:@8141.4]
  assign valid_25_27 = io_inValid_27 & _T_27360; // @[Switch.scala 30:36:@8142.4]
  assign _T_27363 = io_inAddr_28 == 6'h19; // @[Switch.scala 30:53:@8144.4]
  assign valid_25_28 = io_inValid_28 & _T_27363; // @[Switch.scala 30:36:@8145.4]
  assign _T_27366 = io_inAddr_29 == 6'h19; // @[Switch.scala 30:53:@8147.4]
  assign valid_25_29 = io_inValid_29 & _T_27366; // @[Switch.scala 30:36:@8148.4]
  assign _T_27369 = io_inAddr_30 == 6'h19; // @[Switch.scala 30:53:@8150.4]
  assign valid_25_30 = io_inValid_30 & _T_27369; // @[Switch.scala 30:36:@8151.4]
  assign _T_27372 = io_inAddr_31 == 6'h19; // @[Switch.scala 30:53:@8153.4]
  assign valid_25_31 = io_inValid_31 & _T_27372; // @[Switch.scala 30:36:@8154.4]
  assign _T_27375 = io_inAddr_32 == 6'h19; // @[Switch.scala 30:53:@8156.4]
  assign valid_25_32 = io_inValid_32 & _T_27375; // @[Switch.scala 30:36:@8157.4]
  assign _T_27378 = io_inAddr_33 == 6'h19; // @[Switch.scala 30:53:@8159.4]
  assign valid_25_33 = io_inValid_33 & _T_27378; // @[Switch.scala 30:36:@8160.4]
  assign _T_27381 = io_inAddr_34 == 6'h19; // @[Switch.scala 30:53:@8162.4]
  assign valid_25_34 = io_inValid_34 & _T_27381; // @[Switch.scala 30:36:@8163.4]
  assign _T_27384 = io_inAddr_35 == 6'h19; // @[Switch.scala 30:53:@8165.4]
  assign valid_25_35 = io_inValid_35 & _T_27384; // @[Switch.scala 30:36:@8166.4]
  assign _T_27387 = io_inAddr_36 == 6'h19; // @[Switch.scala 30:53:@8168.4]
  assign valid_25_36 = io_inValid_36 & _T_27387; // @[Switch.scala 30:36:@8169.4]
  assign _T_27390 = io_inAddr_37 == 6'h19; // @[Switch.scala 30:53:@8171.4]
  assign valid_25_37 = io_inValid_37 & _T_27390; // @[Switch.scala 30:36:@8172.4]
  assign _T_27393 = io_inAddr_38 == 6'h19; // @[Switch.scala 30:53:@8174.4]
  assign valid_25_38 = io_inValid_38 & _T_27393; // @[Switch.scala 30:36:@8175.4]
  assign _T_27396 = io_inAddr_39 == 6'h19; // @[Switch.scala 30:53:@8177.4]
  assign valid_25_39 = io_inValid_39 & _T_27396; // @[Switch.scala 30:36:@8178.4]
  assign _T_27399 = io_inAddr_40 == 6'h19; // @[Switch.scala 30:53:@8180.4]
  assign valid_25_40 = io_inValid_40 & _T_27399; // @[Switch.scala 30:36:@8181.4]
  assign _T_27402 = io_inAddr_41 == 6'h19; // @[Switch.scala 30:53:@8183.4]
  assign valid_25_41 = io_inValid_41 & _T_27402; // @[Switch.scala 30:36:@8184.4]
  assign _T_27405 = io_inAddr_42 == 6'h19; // @[Switch.scala 30:53:@8186.4]
  assign valid_25_42 = io_inValid_42 & _T_27405; // @[Switch.scala 30:36:@8187.4]
  assign _T_27408 = io_inAddr_43 == 6'h19; // @[Switch.scala 30:53:@8189.4]
  assign valid_25_43 = io_inValid_43 & _T_27408; // @[Switch.scala 30:36:@8190.4]
  assign _T_27411 = io_inAddr_44 == 6'h19; // @[Switch.scala 30:53:@8192.4]
  assign valid_25_44 = io_inValid_44 & _T_27411; // @[Switch.scala 30:36:@8193.4]
  assign _T_27414 = io_inAddr_45 == 6'h19; // @[Switch.scala 30:53:@8195.4]
  assign valid_25_45 = io_inValid_45 & _T_27414; // @[Switch.scala 30:36:@8196.4]
  assign _T_27417 = io_inAddr_46 == 6'h19; // @[Switch.scala 30:53:@8198.4]
  assign valid_25_46 = io_inValid_46 & _T_27417; // @[Switch.scala 30:36:@8199.4]
  assign _T_27420 = io_inAddr_47 == 6'h19; // @[Switch.scala 30:53:@8201.4]
  assign valid_25_47 = io_inValid_47 & _T_27420; // @[Switch.scala 30:36:@8202.4]
  assign _T_27423 = io_inAddr_48 == 6'h19; // @[Switch.scala 30:53:@8204.4]
  assign valid_25_48 = io_inValid_48 & _T_27423; // @[Switch.scala 30:36:@8205.4]
  assign _T_27426 = io_inAddr_49 == 6'h19; // @[Switch.scala 30:53:@8207.4]
  assign valid_25_49 = io_inValid_49 & _T_27426; // @[Switch.scala 30:36:@8208.4]
  assign _T_27429 = io_inAddr_50 == 6'h19; // @[Switch.scala 30:53:@8210.4]
  assign valid_25_50 = io_inValid_50 & _T_27429; // @[Switch.scala 30:36:@8211.4]
  assign _T_27432 = io_inAddr_51 == 6'h19; // @[Switch.scala 30:53:@8213.4]
  assign valid_25_51 = io_inValid_51 & _T_27432; // @[Switch.scala 30:36:@8214.4]
  assign _T_27435 = io_inAddr_52 == 6'h19; // @[Switch.scala 30:53:@8216.4]
  assign valid_25_52 = io_inValid_52 & _T_27435; // @[Switch.scala 30:36:@8217.4]
  assign _T_27438 = io_inAddr_53 == 6'h19; // @[Switch.scala 30:53:@8219.4]
  assign valid_25_53 = io_inValid_53 & _T_27438; // @[Switch.scala 30:36:@8220.4]
  assign _T_27441 = io_inAddr_54 == 6'h19; // @[Switch.scala 30:53:@8222.4]
  assign valid_25_54 = io_inValid_54 & _T_27441; // @[Switch.scala 30:36:@8223.4]
  assign _T_27444 = io_inAddr_55 == 6'h19; // @[Switch.scala 30:53:@8225.4]
  assign valid_25_55 = io_inValid_55 & _T_27444; // @[Switch.scala 30:36:@8226.4]
  assign _T_27447 = io_inAddr_56 == 6'h19; // @[Switch.scala 30:53:@8228.4]
  assign valid_25_56 = io_inValid_56 & _T_27447; // @[Switch.scala 30:36:@8229.4]
  assign _T_27450 = io_inAddr_57 == 6'h19; // @[Switch.scala 30:53:@8231.4]
  assign valid_25_57 = io_inValid_57 & _T_27450; // @[Switch.scala 30:36:@8232.4]
  assign _T_27453 = io_inAddr_58 == 6'h19; // @[Switch.scala 30:53:@8234.4]
  assign valid_25_58 = io_inValid_58 & _T_27453; // @[Switch.scala 30:36:@8235.4]
  assign _T_27456 = io_inAddr_59 == 6'h19; // @[Switch.scala 30:53:@8237.4]
  assign valid_25_59 = io_inValid_59 & _T_27456; // @[Switch.scala 30:36:@8238.4]
  assign _T_27459 = io_inAddr_60 == 6'h19; // @[Switch.scala 30:53:@8240.4]
  assign valid_25_60 = io_inValid_60 & _T_27459; // @[Switch.scala 30:36:@8241.4]
  assign _T_27462 = io_inAddr_61 == 6'h19; // @[Switch.scala 30:53:@8243.4]
  assign valid_25_61 = io_inValid_61 & _T_27462; // @[Switch.scala 30:36:@8244.4]
  assign _T_27465 = io_inAddr_62 == 6'h19; // @[Switch.scala 30:53:@8246.4]
  assign valid_25_62 = io_inValid_62 & _T_27465; // @[Switch.scala 30:36:@8247.4]
  assign _T_27468 = io_inAddr_63 == 6'h19; // @[Switch.scala 30:53:@8249.4]
  assign valid_25_63 = io_inValid_63 & _T_27468; // @[Switch.scala 30:36:@8250.4]
  assign _T_27534 = valid_25_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@8252.4]
  assign _T_27535 = valid_25_61 ? 6'h3d : _T_27534; // @[Mux.scala 31:69:@8253.4]
  assign _T_27536 = valid_25_60 ? 6'h3c : _T_27535; // @[Mux.scala 31:69:@8254.4]
  assign _T_27537 = valid_25_59 ? 6'h3b : _T_27536; // @[Mux.scala 31:69:@8255.4]
  assign _T_27538 = valid_25_58 ? 6'h3a : _T_27537; // @[Mux.scala 31:69:@8256.4]
  assign _T_27539 = valid_25_57 ? 6'h39 : _T_27538; // @[Mux.scala 31:69:@8257.4]
  assign _T_27540 = valid_25_56 ? 6'h38 : _T_27539; // @[Mux.scala 31:69:@8258.4]
  assign _T_27541 = valid_25_55 ? 6'h37 : _T_27540; // @[Mux.scala 31:69:@8259.4]
  assign _T_27542 = valid_25_54 ? 6'h36 : _T_27541; // @[Mux.scala 31:69:@8260.4]
  assign _T_27543 = valid_25_53 ? 6'h35 : _T_27542; // @[Mux.scala 31:69:@8261.4]
  assign _T_27544 = valid_25_52 ? 6'h34 : _T_27543; // @[Mux.scala 31:69:@8262.4]
  assign _T_27545 = valid_25_51 ? 6'h33 : _T_27544; // @[Mux.scala 31:69:@8263.4]
  assign _T_27546 = valid_25_50 ? 6'h32 : _T_27545; // @[Mux.scala 31:69:@8264.4]
  assign _T_27547 = valid_25_49 ? 6'h31 : _T_27546; // @[Mux.scala 31:69:@8265.4]
  assign _T_27548 = valid_25_48 ? 6'h30 : _T_27547; // @[Mux.scala 31:69:@8266.4]
  assign _T_27549 = valid_25_47 ? 6'h2f : _T_27548; // @[Mux.scala 31:69:@8267.4]
  assign _T_27550 = valid_25_46 ? 6'h2e : _T_27549; // @[Mux.scala 31:69:@8268.4]
  assign _T_27551 = valid_25_45 ? 6'h2d : _T_27550; // @[Mux.scala 31:69:@8269.4]
  assign _T_27552 = valid_25_44 ? 6'h2c : _T_27551; // @[Mux.scala 31:69:@8270.4]
  assign _T_27553 = valid_25_43 ? 6'h2b : _T_27552; // @[Mux.scala 31:69:@8271.4]
  assign _T_27554 = valid_25_42 ? 6'h2a : _T_27553; // @[Mux.scala 31:69:@8272.4]
  assign _T_27555 = valid_25_41 ? 6'h29 : _T_27554; // @[Mux.scala 31:69:@8273.4]
  assign _T_27556 = valid_25_40 ? 6'h28 : _T_27555; // @[Mux.scala 31:69:@8274.4]
  assign _T_27557 = valid_25_39 ? 6'h27 : _T_27556; // @[Mux.scala 31:69:@8275.4]
  assign _T_27558 = valid_25_38 ? 6'h26 : _T_27557; // @[Mux.scala 31:69:@8276.4]
  assign _T_27559 = valid_25_37 ? 6'h25 : _T_27558; // @[Mux.scala 31:69:@8277.4]
  assign _T_27560 = valid_25_36 ? 6'h24 : _T_27559; // @[Mux.scala 31:69:@8278.4]
  assign _T_27561 = valid_25_35 ? 6'h23 : _T_27560; // @[Mux.scala 31:69:@8279.4]
  assign _T_27562 = valid_25_34 ? 6'h22 : _T_27561; // @[Mux.scala 31:69:@8280.4]
  assign _T_27563 = valid_25_33 ? 6'h21 : _T_27562; // @[Mux.scala 31:69:@8281.4]
  assign _T_27564 = valid_25_32 ? 6'h20 : _T_27563; // @[Mux.scala 31:69:@8282.4]
  assign _T_27565 = valid_25_31 ? 6'h1f : _T_27564; // @[Mux.scala 31:69:@8283.4]
  assign _T_27566 = valid_25_30 ? 6'h1e : _T_27565; // @[Mux.scala 31:69:@8284.4]
  assign _T_27567 = valid_25_29 ? 6'h1d : _T_27566; // @[Mux.scala 31:69:@8285.4]
  assign _T_27568 = valid_25_28 ? 6'h1c : _T_27567; // @[Mux.scala 31:69:@8286.4]
  assign _T_27569 = valid_25_27 ? 6'h1b : _T_27568; // @[Mux.scala 31:69:@8287.4]
  assign _T_27570 = valid_25_26 ? 6'h1a : _T_27569; // @[Mux.scala 31:69:@8288.4]
  assign _T_27571 = valid_25_25 ? 6'h19 : _T_27570; // @[Mux.scala 31:69:@8289.4]
  assign _T_27572 = valid_25_24 ? 6'h18 : _T_27571; // @[Mux.scala 31:69:@8290.4]
  assign _T_27573 = valid_25_23 ? 6'h17 : _T_27572; // @[Mux.scala 31:69:@8291.4]
  assign _T_27574 = valid_25_22 ? 6'h16 : _T_27573; // @[Mux.scala 31:69:@8292.4]
  assign _T_27575 = valid_25_21 ? 6'h15 : _T_27574; // @[Mux.scala 31:69:@8293.4]
  assign _T_27576 = valid_25_20 ? 6'h14 : _T_27575; // @[Mux.scala 31:69:@8294.4]
  assign _T_27577 = valid_25_19 ? 6'h13 : _T_27576; // @[Mux.scala 31:69:@8295.4]
  assign _T_27578 = valid_25_18 ? 6'h12 : _T_27577; // @[Mux.scala 31:69:@8296.4]
  assign _T_27579 = valid_25_17 ? 6'h11 : _T_27578; // @[Mux.scala 31:69:@8297.4]
  assign _T_27580 = valid_25_16 ? 6'h10 : _T_27579; // @[Mux.scala 31:69:@8298.4]
  assign _T_27581 = valid_25_15 ? 6'hf : _T_27580; // @[Mux.scala 31:69:@8299.4]
  assign _T_27582 = valid_25_14 ? 6'he : _T_27581; // @[Mux.scala 31:69:@8300.4]
  assign _T_27583 = valid_25_13 ? 6'hd : _T_27582; // @[Mux.scala 31:69:@8301.4]
  assign _T_27584 = valid_25_12 ? 6'hc : _T_27583; // @[Mux.scala 31:69:@8302.4]
  assign _T_27585 = valid_25_11 ? 6'hb : _T_27584; // @[Mux.scala 31:69:@8303.4]
  assign _T_27586 = valid_25_10 ? 6'ha : _T_27585; // @[Mux.scala 31:69:@8304.4]
  assign _T_27587 = valid_25_9 ? 6'h9 : _T_27586; // @[Mux.scala 31:69:@8305.4]
  assign _T_27588 = valid_25_8 ? 6'h8 : _T_27587; // @[Mux.scala 31:69:@8306.4]
  assign _T_27589 = valid_25_7 ? 6'h7 : _T_27588; // @[Mux.scala 31:69:@8307.4]
  assign _T_27590 = valid_25_6 ? 6'h6 : _T_27589; // @[Mux.scala 31:69:@8308.4]
  assign _T_27591 = valid_25_5 ? 6'h5 : _T_27590; // @[Mux.scala 31:69:@8309.4]
  assign _T_27592 = valid_25_4 ? 6'h4 : _T_27591; // @[Mux.scala 31:69:@8310.4]
  assign _T_27593 = valid_25_3 ? 6'h3 : _T_27592; // @[Mux.scala 31:69:@8311.4]
  assign _T_27594 = valid_25_2 ? 6'h2 : _T_27593; // @[Mux.scala 31:69:@8312.4]
  assign _T_27595 = valid_25_1 ? 6'h1 : _T_27594; // @[Mux.scala 31:69:@8313.4]
  assign select_25 = valid_25_0 ? 6'h0 : _T_27595; // @[Mux.scala 31:69:@8314.4]
  assign _GEN_1601 = 6'h1 == select_25 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1602 = 6'h2 == select_25 ? io_inData_2 : _GEN_1601; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1603 = 6'h3 == select_25 ? io_inData_3 : _GEN_1602; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1604 = 6'h4 == select_25 ? io_inData_4 : _GEN_1603; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1605 = 6'h5 == select_25 ? io_inData_5 : _GEN_1604; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1606 = 6'h6 == select_25 ? io_inData_6 : _GEN_1605; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1607 = 6'h7 == select_25 ? io_inData_7 : _GEN_1606; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1608 = 6'h8 == select_25 ? io_inData_8 : _GEN_1607; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1609 = 6'h9 == select_25 ? io_inData_9 : _GEN_1608; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1610 = 6'ha == select_25 ? io_inData_10 : _GEN_1609; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1611 = 6'hb == select_25 ? io_inData_11 : _GEN_1610; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1612 = 6'hc == select_25 ? io_inData_12 : _GEN_1611; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1613 = 6'hd == select_25 ? io_inData_13 : _GEN_1612; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1614 = 6'he == select_25 ? io_inData_14 : _GEN_1613; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1615 = 6'hf == select_25 ? io_inData_15 : _GEN_1614; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1616 = 6'h10 == select_25 ? io_inData_16 : _GEN_1615; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1617 = 6'h11 == select_25 ? io_inData_17 : _GEN_1616; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1618 = 6'h12 == select_25 ? io_inData_18 : _GEN_1617; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1619 = 6'h13 == select_25 ? io_inData_19 : _GEN_1618; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1620 = 6'h14 == select_25 ? io_inData_20 : _GEN_1619; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1621 = 6'h15 == select_25 ? io_inData_21 : _GEN_1620; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1622 = 6'h16 == select_25 ? io_inData_22 : _GEN_1621; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1623 = 6'h17 == select_25 ? io_inData_23 : _GEN_1622; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1624 = 6'h18 == select_25 ? io_inData_24 : _GEN_1623; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1625 = 6'h19 == select_25 ? io_inData_25 : _GEN_1624; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1626 = 6'h1a == select_25 ? io_inData_26 : _GEN_1625; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1627 = 6'h1b == select_25 ? io_inData_27 : _GEN_1626; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1628 = 6'h1c == select_25 ? io_inData_28 : _GEN_1627; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1629 = 6'h1d == select_25 ? io_inData_29 : _GEN_1628; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1630 = 6'h1e == select_25 ? io_inData_30 : _GEN_1629; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1631 = 6'h1f == select_25 ? io_inData_31 : _GEN_1630; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1632 = 6'h20 == select_25 ? io_inData_32 : _GEN_1631; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1633 = 6'h21 == select_25 ? io_inData_33 : _GEN_1632; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1634 = 6'h22 == select_25 ? io_inData_34 : _GEN_1633; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1635 = 6'h23 == select_25 ? io_inData_35 : _GEN_1634; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1636 = 6'h24 == select_25 ? io_inData_36 : _GEN_1635; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1637 = 6'h25 == select_25 ? io_inData_37 : _GEN_1636; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1638 = 6'h26 == select_25 ? io_inData_38 : _GEN_1637; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1639 = 6'h27 == select_25 ? io_inData_39 : _GEN_1638; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1640 = 6'h28 == select_25 ? io_inData_40 : _GEN_1639; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1641 = 6'h29 == select_25 ? io_inData_41 : _GEN_1640; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1642 = 6'h2a == select_25 ? io_inData_42 : _GEN_1641; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1643 = 6'h2b == select_25 ? io_inData_43 : _GEN_1642; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1644 = 6'h2c == select_25 ? io_inData_44 : _GEN_1643; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1645 = 6'h2d == select_25 ? io_inData_45 : _GEN_1644; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1646 = 6'h2e == select_25 ? io_inData_46 : _GEN_1645; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1647 = 6'h2f == select_25 ? io_inData_47 : _GEN_1646; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1648 = 6'h30 == select_25 ? io_inData_48 : _GEN_1647; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1649 = 6'h31 == select_25 ? io_inData_49 : _GEN_1648; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1650 = 6'h32 == select_25 ? io_inData_50 : _GEN_1649; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1651 = 6'h33 == select_25 ? io_inData_51 : _GEN_1650; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1652 = 6'h34 == select_25 ? io_inData_52 : _GEN_1651; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1653 = 6'h35 == select_25 ? io_inData_53 : _GEN_1652; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1654 = 6'h36 == select_25 ? io_inData_54 : _GEN_1653; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1655 = 6'h37 == select_25 ? io_inData_55 : _GEN_1654; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1656 = 6'h38 == select_25 ? io_inData_56 : _GEN_1655; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1657 = 6'h39 == select_25 ? io_inData_57 : _GEN_1656; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1658 = 6'h3a == select_25 ? io_inData_58 : _GEN_1657; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1659 = 6'h3b == select_25 ? io_inData_59 : _GEN_1658; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1660 = 6'h3c == select_25 ? io_inData_60 : _GEN_1659; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1661 = 6'h3d == select_25 ? io_inData_61 : _GEN_1660; // @[Switch.scala 33:19:@8316.4]
  assign _GEN_1662 = 6'h3e == select_25 ? io_inData_62 : _GEN_1661; // @[Switch.scala 33:19:@8316.4]
  assign _T_27604 = {valid_25_7,valid_25_6,valid_25_5,valid_25_4,valid_25_3,valid_25_2,valid_25_1,valid_25_0}; // @[Switch.scala 34:32:@8323.4]
  assign _T_27612 = {valid_25_15,valid_25_14,valid_25_13,valid_25_12,valid_25_11,valid_25_10,valid_25_9,valid_25_8,_T_27604}; // @[Switch.scala 34:32:@8331.4]
  assign _T_27619 = {valid_25_23,valid_25_22,valid_25_21,valid_25_20,valid_25_19,valid_25_18,valid_25_17,valid_25_16}; // @[Switch.scala 34:32:@8338.4]
  assign _T_27628 = {valid_25_31,valid_25_30,valid_25_29,valid_25_28,valid_25_27,valid_25_26,valid_25_25,valid_25_24,_T_27619,_T_27612}; // @[Switch.scala 34:32:@8347.4]
  assign _T_27635 = {valid_25_39,valid_25_38,valid_25_37,valid_25_36,valid_25_35,valid_25_34,valid_25_33,valid_25_32}; // @[Switch.scala 34:32:@8354.4]
  assign _T_27643 = {valid_25_47,valid_25_46,valid_25_45,valid_25_44,valid_25_43,valid_25_42,valid_25_41,valid_25_40,_T_27635}; // @[Switch.scala 34:32:@8362.4]
  assign _T_27650 = {valid_25_55,valid_25_54,valid_25_53,valid_25_52,valid_25_51,valid_25_50,valid_25_49,valid_25_48}; // @[Switch.scala 34:32:@8369.4]
  assign _T_27659 = {valid_25_63,valid_25_62,valid_25_61,valid_25_60,valid_25_59,valid_25_58,valid_25_57,valid_25_56,_T_27650,_T_27643}; // @[Switch.scala 34:32:@8378.4]
  assign _T_27660 = {_T_27659,_T_27628}; // @[Switch.scala 34:32:@8379.4]
  assign _T_27664 = io_inAddr_0 == 6'h1a; // @[Switch.scala 30:53:@8382.4]
  assign valid_26_0 = io_inValid_0 & _T_27664; // @[Switch.scala 30:36:@8383.4]
  assign _T_27667 = io_inAddr_1 == 6'h1a; // @[Switch.scala 30:53:@8385.4]
  assign valid_26_1 = io_inValid_1 & _T_27667; // @[Switch.scala 30:36:@8386.4]
  assign _T_27670 = io_inAddr_2 == 6'h1a; // @[Switch.scala 30:53:@8388.4]
  assign valid_26_2 = io_inValid_2 & _T_27670; // @[Switch.scala 30:36:@8389.4]
  assign _T_27673 = io_inAddr_3 == 6'h1a; // @[Switch.scala 30:53:@8391.4]
  assign valid_26_3 = io_inValid_3 & _T_27673; // @[Switch.scala 30:36:@8392.4]
  assign _T_27676 = io_inAddr_4 == 6'h1a; // @[Switch.scala 30:53:@8394.4]
  assign valid_26_4 = io_inValid_4 & _T_27676; // @[Switch.scala 30:36:@8395.4]
  assign _T_27679 = io_inAddr_5 == 6'h1a; // @[Switch.scala 30:53:@8397.4]
  assign valid_26_5 = io_inValid_5 & _T_27679; // @[Switch.scala 30:36:@8398.4]
  assign _T_27682 = io_inAddr_6 == 6'h1a; // @[Switch.scala 30:53:@8400.4]
  assign valid_26_6 = io_inValid_6 & _T_27682; // @[Switch.scala 30:36:@8401.4]
  assign _T_27685 = io_inAddr_7 == 6'h1a; // @[Switch.scala 30:53:@8403.4]
  assign valid_26_7 = io_inValid_7 & _T_27685; // @[Switch.scala 30:36:@8404.4]
  assign _T_27688 = io_inAddr_8 == 6'h1a; // @[Switch.scala 30:53:@8406.4]
  assign valid_26_8 = io_inValid_8 & _T_27688; // @[Switch.scala 30:36:@8407.4]
  assign _T_27691 = io_inAddr_9 == 6'h1a; // @[Switch.scala 30:53:@8409.4]
  assign valid_26_9 = io_inValid_9 & _T_27691; // @[Switch.scala 30:36:@8410.4]
  assign _T_27694 = io_inAddr_10 == 6'h1a; // @[Switch.scala 30:53:@8412.4]
  assign valid_26_10 = io_inValid_10 & _T_27694; // @[Switch.scala 30:36:@8413.4]
  assign _T_27697 = io_inAddr_11 == 6'h1a; // @[Switch.scala 30:53:@8415.4]
  assign valid_26_11 = io_inValid_11 & _T_27697; // @[Switch.scala 30:36:@8416.4]
  assign _T_27700 = io_inAddr_12 == 6'h1a; // @[Switch.scala 30:53:@8418.4]
  assign valid_26_12 = io_inValid_12 & _T_27700; // @[Switch.scala 30:36:@8419.4]
  assign _T_27703 = io_inAddr_13 == 6'h1a; // @[Switch.scala 30:53:@8421.4]
  assign valid_26_13 = io_inValid_13 & _T_27703; // @[Switch.scala 30:36:@8422.4]
  assign _T_27706 = io_inAddr_14 == 6'h1a; // @[Switch.scala 30:53:@8424.4]
  assign valid_26_14 = io_inValid_14 & _T_27706; // @[Switch.scala 30:36:@8425.4]
  assign _T_27709 = io_inAddr_15 == 6'h1a; // @[Switch.scala 30:53:@8427.4]
  assign valid_26_15 = io_inValid_15 & _T_27709; // @[Switch.scala 30:36:@8428.4]
  assign _T_27712 = io_inAddr_16 == 6'h1a; // @[Switch.scala 30:53:@8430.4]
  assign valid_26_16 = io_inValid_16 & _T_27712; // @[Switch.scala 30:36:@8431.4]
  assign _T_27715 = io_inAddr_17 == 6'h1a; // @[Switch.scala 30:53:@8433.4]
  assign valid_26_17 = io_inValid_17 & _T_27715; // @[Switch.scala 30:36:@8434.4]
  assign _T_27718 = io_inAddr_18 == 6'h1a; // @[Switch.scala 30:53:@8436.4]
  assign valid_26_18 = io_inValid_18 & _T_27718; // @[Switch.scala 30:36:@8437.4]
  assign _T_27721 = io_inAddr_19 == 6'h1a; // @[Switch.scala 30:53:@8439.4]
  assign valid_26_19 = io_inValid_19 & _T_27721; // @[Switch.scala 30:36:@8440.4]
  assign _T_27724 = io_inAddr_20 == 6'h1a; // @[Switch.scala 30:53:@8442.4]
  assign valid_26_20 = io_inValid_20 & _T_27724; // @[Switch.scala 30:36:@8443.4]
  assign _T_27727 = io_inAddr_21 == 6'h1a; // @[Switch.scala 30:53:@8445.4]
  assign valid_26_21 = io_inValid_21 & _T_27727; // @[Switch.scala 30:36:@8446.4]
  assign _T_27730 = io_inAddr_22 == 6'h1a; // @[Switch.scala 30:53:@8448.4]
  assign valid_26_22 = io_inValid_22 & _T_27730; // @[Switch.scala 30:36:@8449.4]
  assign _T_27733 = io_inAddr_23 == 6'h1a; // @[Switch.scala 30:53:@8451.4]
  assign valid_26_23 = io_inValid_23 & _T_27733; // @[Switch.scala 30:36:@8452.4]
  assign _T_27736 = io_inAddr_24 == 6'h1a; // @[Switch.scala 30:53:@8454.4]
  assign valid_26_24 = io_inValid_24 & _T_27736; // @[Switch.scala 30:36:@8455.4]
  assign _T_27739 = io_inAddr_25 == 6'h1a; // @[Switch.scala 30:53:@8457.4]
  assign valid_26_25 = io_inValid_25 & _T_27739; // @[Switch.scala 30:36:@8458.4]
  assign _T_27742 = io_inAddr_26 == 6'h1a; // @[Switch.scala 30:53:@8460.4]
  assign valid_26_26 = io_inValid_26 & _T_27742; // @[Switch.scala 30:36:@8461.4]
  assign _T_27745 = io_inAddr_27 == 6'h1a; // @[Switch.scala 30:53:@8463.4]
  assign valid_26_27 = io_inValid_27 & _T_27745; // @[Switch.scala 30:36:@8464.4]
  assign _T_27748 = io_inAddr_28 == 6'h1a; // @[Switch.scala 30:53:@8466.4]
  assign valid_26_28 = io_inValid_28 & _T_27748; // @[Switch.scala 30:36:@8467.4]
  assign _T_27751 = io_inAddr_29 == 6'h1a; // @[Switch.scala 30:53:@8469.4]
  assign valid_26_29 = io_inValid_29 & _T_27751; // @[Switch.scala 30:36:@8470.4]
  assign _T_27754 = io_inAddr_30 == 6'h1a; // @[Switch.scala 30:53:@8472.4]
  assign valid_26_30 = io_inValid_30 & _T_27754; // @[Switch.scala 30:36:@8473.4]
  assign _T_27757 = io_inAddr_31 == 6'h1a; // @[Switch.scala 30:53:@8475.4]
  assign valid_26_31 = io_inValid_31 & _T_27757; // @[Switch.scala 30:36:@8476.4]
  assign _T_27760 = io_inAddr_32 == 6'h1a; // @[Switch.scala 30:53:@8478.4]
  assign valid_26_32 = io_inValid_32 & _T_27760; // @[Switch.scala 30:36:@8479.4]
  assign _T_27763 = io_inAddr_33 == 6'h1a; // @[Switch.scala 30:53:@8481.4]
  assign valid_26_33 = io_inValid_33 & _T_27763; // @[Switch.scala 30:36:@8482.4]
  assign _T_27766 = io_inAddr_34 == 6'h1a; // @[Switch.scala 30:53:@8484.4]
  assign valid_26_34 = io_inValid_34 & _T_27766; // @[Switch.scala 30:36:@8485.4]
  assign _T_27769 = io_inAddr_35 == 6'h1a; // @[Switch.scala 30:53:@8487.4]
  assign valid_26_35 = io_inValid_35 & _T_27769; // @[Switch.scala 30:36:@8488.4]
  assign _T_27772 = io_inAddr_36 == 6'h1a; // @[Switch.scala 30:53:@8490.4]
  assign valid_26_36 = io_inValid_36 & _T_27772; // @[Switch.scala 30:36:@8491.4]
  assign _T_27775 = io_inAddr_37 == 6'h1a; // @[Switch.scala 30:53:@8493.4]
  assign valid_26_37 = io_inValid_37 & _T_27775; // @[Switch.scala 30:36:@8494.4]
  assign _T_27778 = io_inAddr_38 == 6'h1a; // @[Switch.scala 30:53:@8496.4]
  assign valid_26_38 = io_inValid_38 & _T_27778; // @[Switch.scala 30:36:@8497.4]
  assign _T_27781 = io_inAddr_39 == 6'h1a; // @[Switch.scala 30:53:@8499.4]
  assign valid_26_39 = io_inValid_39 & _T_27781; // @[Switch.scala 30:36:@8500.4]
  assign _T_27784 = io_inAddr_40 == 6'h1a; // @[Switch.scala 30:53:@8502.4]
  assign valid_26_40 = io_inValid_40 & _T_27784; // @[Switch.scala 30:36:@8503.4]
  assign _T_27787 = io_inAddr_41 == 6'h1a; // @[Switch.scala 30:53:@8505.4]
  assign valid_26_41 = io_inValid_41 & _T_27787; // @[Switch.scala 30:36:@8506.4]
  assign _T_27790 = io_inAddr_42 == 6'h1a; // @[Switch.scala 30:53:@8508.4]
  assign valid_26_42 = io_inValid_42 & _T_27790; // @[Switch.scala 30:36:@8509.4]
  assign _T_27793 = io_inAddr_43 == 6'h1a; // @[Switch.scala 30:53:@8511.4]
  assign valid_26_43 = io_inValid_43 & _T_27793; // @[Switch.scala 30:36:@8512.4]
  assign _T_27796 = io_inAddr_44 == 6'h1a; // @[Switch.scala 30:53:@8514.4]
  assign valid_26_44 = io_inValid_44 & _T_27796; // @[Switch.scala 30:36:@8515.4]
  assign _T_27799 = io_inAddr_45 == 6'h1a; // @[Switch.scala 30:53:@8517.4]
  assign valid_26_45 = io_inValid_45 & _T_27799; // @[Switch.scala 30:36:@8518.4]
  assign _T_27802 = io_inAddr_46 == 6'h1a; // @[Switch.scala 30:53:@8520.4]
  assign valid_26_46 = io_inValid_46 & _T_27802; // @[Switch.scala 30:36:@8521.4]
  assign _T_27805 = io_inAddr_47 == 6'h1a; // @[Switch.scala 30:53:@8523.4]
  assign valid_26_47 = io_inValid_47 & _T_27805; // @[Switch.scala 30:36:@8524.4]
  assign _T_27808 = io_inAddr_48 == 6'h1a; // @[Switch.scala 30:53:@8526.4]
  assign valid_26_48 = io_inValid_48 & _T_27808; // @[Switch.scala 30:36:@8527.4]
  assign _T_27811 = io_inAddr_49 == 6'h1a; // @[Switch.scala 30:53:@8529.4]
  assign valid_26_49 = io_inValid_49 & _T_27811; // @[Switch.scala 30:36:@8530.4]
  assign _T_27814 = io_inAddr_50 == 6'h1a; // @[Switch.scala 30:53:@8532.4]
  assign valid_26_50 = io_inValid_50 & _T_27814; // @[Switch.scala 30:36:@8533.4]
  assign _T_27817 = io_inAddr_51 == 6'h1a; // @[Switch.scala 30:53:@8535.4]
  assign valid_26_51 = io_inValid_51 & _T_27817; // @[Switch.scala 30:36:@8536.4]
  assign _T_27820 = io_inAddr_52 == 6'h1a; // @[Switch.scala 30:53:@8538.4]
  assign valid_26_52 = io_inValid_52 & _T_27820; // @[Switch.scala 30:36:@8539.4]
  assign _T_27823 = io_inAddr_53 == 6'h1a; // @[Switch.scala 30:53:@8541.4]
  assign valid_26_53 = io_inValid_53 & _T_27823; // @[Switch.scala 30:36:@8542.4]
  assign _T_27826 = io_inAddr_54 == 6'h1a; // @[Switch.scala 30:53:@8544.4]
  assign valid_26_54 = io_inValid_54 & _T_27826; // @[Switch.scala 30:36:@8545.4]
  assign _T_27829 = io_inAddr_55 == 6'h1a; // @[Switch.scala 30:53:@8547.4]
  assign valid_26_55 = io_inValid_55 & _T_27829; // @[Switch.scala 30:36:@8548.4]
  assign _T_27832 = io_inAddr_56 == 6'h1a; // @[Switch.scala 30:53:@8550.4]
  assign valid_26_56 = io_inValid_56 & _T_27832; // @[Switch.scala 30:36:@8551.4]
  assign _T_27835 = io_inAddr_57 == 6'h1a; // @[Switch.scala 30:53:@8553.4]
  assign valid_26_57 = io_inValid_57 & _T_27835; // @[Switch.scala 30:36:@8554.4]
  assign _T_27838 = io_inAddr_58 == 6'h1a; // @[Switch.scala 30:53:@8556.4]
  assign valid_26_58 = io_inValid_58 & _T_27838; // @[Switch.scala 30:36:@8557.4]
  assign _T_27841 = io_inAddr_59 == 6'h1a; // @[Switch.scala 30:53:@8559.4]
  assign valid_26_59 = io_inValid_59 & _T_27841; // @[Switch.scala 30:36:@8560.4]
  assign _T_27844 = io_inAddr_60 == 6'h1a; // @[Switch.scala 30:53:@8562.4]
  assign valid_26_60 = io_inValid_60 & _T_27844; // @[Switch.scala 30:36:@8563.4]
  assign _T_27847 = io_inAddr_61 == 6'h1a; // @[Switch.scala 30:53:@8565.4]
  assign valid_26_61 = io_inValid_61 & _T_27847; // @[Switch.scala 30:36:@8566.4]
  assign _T_27850 = io_inAddr_62 == 6'h1a; // @[Switch.scala 30:53:@8568.4]
  assign valid_26_62 = io_inValid_62 & _T_27850; // @[Switch.scala 30:36:@8569.4]
  assign _T_27853 = io_inAddr_63 == 6'h1a; // @[Switch.scala 30:53:@8571.4]
  assign valid_26_63 = io_inValid_63 & _T_27853; // @[Switch.scala 30:36:@8572.4]
  assign _T_27919 = valid_26_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@8574.4]
  assign _T_27920 = valid_26_61 ? 6'h3d : _T_27919; // @[Mux.scala 31:69:@8575.4]
  assign _T_27921 = valid_26_60 ? 6'h3c : _T_27920; // @[Mux.scala 31:69:@8576.4]
  assign _T_27922 = valid_26_59 ? 6'h3b : _T_27921; // @[Mux.scala 31:69:@8577.4]
  assign _T_27923 = valid_26_58 ? 6'h3a : _T_27922; // @[Mux.scala 31:69:@8578.4]
  assign _T_27924 = valid_26_57 ? 6'h39 : _T_27923; // @[Mux.scala 31:69:@8579.4]
  assign _T_27925 = valid_26_56 ? 6'h38 : _T_27924; // @[Mux.scala 31:69:@8580.4]
  assign _T_27926 = valid_26_55 ? 6'h37 : _T_27925; // @[Mux.scala 31:69:@8581.4]
  assign _T_27927 = valid_26_54 ? 6'h36 : _T_27926; // @[Mux.scala 31:69:@8582.4]
  assign _T_27928 = valid_26_53 ? 6'h35 : _T_27927; // @[Mux.scala 31:69:@8583.4]
  assign _T_27929 = valid_26_52 ? 6'h34 : _T_27928; // @[Mux.scala 31:69:@8584.4]
  assign _T_27930 = valid_26_51 ? 6'h33 : _T_27929; // @[Mux.scala 31:69:@8585.4]
  assign _T_27931 = valid_26_50 ? 6'h32 : _T_27930; // @[Mux.scala 31:69:@8586.4]
  assign _T_27932 = valid_26_49 ? 6'h31 : _T_27931; // @[Mux.scala 31:69:@8587.4]
  assign _T_27933 = valid_26_48 ? 6'h30 : _T_27932; // @[Mux.scala 31:69:@8588.4]
  assign _T_27934 = valid_26_47 ? 6'h2f : _T_27933; // @[Mux.scala 31:69:@8589.4]
  assign _T_27935 = valid_26_46 ? 6'h2e : _T_27934; // @[Mux.scala 31:69:@8590.4]
  assign _T_27936 = valid_26_45 ? 6'h2d : _T_27935; // @[Mux.scala 31:69:@8591.4]
  assign _T_27937 = valid_26_44 ? 6'h2c : _T_27936; // @[Mux.scala 31:69:@8592.4]
  assign _T_27938 = valid_26_43 ? 6'h2b : _T_27937; // @[Mux.scala 31:69:@8593.4]
  assign _T_27939 = valid_26_42 ? 6'h2a : _T_27938; // @[Mux.scala 31:69:@8594.4]
  assign _T_27940 = valid_26_41 ? 6'h29 : _T_27939; // @[Mux.scala 31:69:@8595.4]
  assign _T_27941 = valid_26_40 ? 6'h28 : _T_27940; // @[Mux.scala 31:69:@8596.4]
  assign _T_27942 = valid_26_39 ? 6'h27 : _T_27941; // @[Mux.scala 31:69:@8597.4]
  assign _T_27943 = valid_26_38 ? 6'h26 : _T_27942; // @[Mux.scala 31:69:@8598.4]
  assign _T_27944 = valid_26_37 ? 6'h25 : _T_27943; // @[Mux.scala 31:69:@8599.4]
  assign _T_27945 = valid_26_36 ? 6'h24 : _T_27944; // @[Mux.scala 31:69:@8600.4]
  assign _T_27946 = valid_26_35 ? 6'h23 : _T_27945; // @[Mux.scala 31:69:@8601.4]
  assign _T_27947 = valid_26_34 ? 6'h22 : _T_27946; // @[Mux.scala 31:69:@8602.4]
  assign _T_27948 = valid_26_33 ? 6'h21 : _T_27947; // @[Mux.scala 31:69:@8603.4]
  assign _T_27949 = valid_26_32 ? 6'h20 : _T_27948; // @[Mux.scala 31:69:@8604.4]
  assign _T_27950 = valid_26_31 ? 6'h1f : _T_27949; // @[Mux.scala 31:69:@8605.4]
  assign _T_27951 = valid_26_30 ? 6'h1e : _T_27950; // @[Mux.scala 31:69:@8606.4]
  assign _T_27952 = valid_26_29 ? 6'h1d : _T_27951; // @[Mux.scala 31:69:@8607.4]
  assign _T_27953 = valid_26_28 ? 6'h1c : _T_27952; // @[Mux.scala 31:69:@8608.4]
  assign _T_27954 = valid_26_27 ? 6'h1b : _T_27953; // @[Mux.scala 31:69:@8609.4]
  assign _T_27955 = valid_26_26 ? 6'h1a : _T_27954; // @[Mux.scala 31:69:@8610.4]
  assign _T_27956 = valid_26_25 ? 6'h19 : _T_27955; // @[Mux.scala 31:69:@8611.4]
  assign _T_27957 = valid_26_24 ? 6'h18 : _T_27956; // @[Mux.scala 31:69:@8612.4]
  assign _T_27958 = valid_26_23 ? 6'h17 : _T_27957; // @[Mux.scala 31:69:@8613.4]
  assign _T_27959 = valid_26_22 ? 6'h16 : _T_27958; // @[Mux.scala 31:69:@8614.4]
  assign _T_27960 = valid_26_21 ? 6'h15 : _T_27959; // @[Mux.scala 31:69:@8615.4]
  assign _T_27961 = valid_26_20 ? 6'h14 : _T_27960; // @[Mux.scala 31:69:@8616.4]
  assign _T_27962 = valid_26_19 ? 6'h13 : _T_27961; // @[Mux.scala 31:69:@8617.4]
  assign _T_27963 = valid_26_18 ? 6'h12 : _T_27962; // @[Mux.scala 31:69:@8618.4]
  assign _T_27964 = valid_26_17 ? 6'h11 : _T_27963; // @[Mux.scala 31:69:@8619.4]
  assign _T_27965 = valid_26_16 ? 6'h10 : _T_27964; // @[Mux.scala 31:69:@8620.4]
  assign _T_27966 = valid_26_15 ? 6'hf : _T_27965; // @[Mux.scala 31:69:@8621.4]
  assign _T_27967 = valid_26_14 ? 6'he : _T_27966; // @[Mux.scala 31:69:@8622.4]
  assign _T_27968 = valid_26_13 ? 6'hd : _T_27967; // @[Mux.scala 31:69:@8623.4]
  assign _T_27969 = valid_26_12 ? 6'hc : _T_27968; // @[Mux.scala 31:69:@8624.4]
  assign _T_27970 = valid_26_11 ? 6'hb : _T_27969; // @[Mux.scala 31:69:@8625.4]
  assign _T_27971 = valid_26_10 ? 6'ha : _T_27970; // @[Mux.scala 31:69:@8626.4]
  assign _T_27972 = valid_26_9 ? 6'h9 : _T_27971; // @[Mux.scala 31:69:@8627.4]
  assign _T_27973 = valid_26_8 ? 6'h8 : _T_27972; // @[Mux.scala 31:69:@8628.4]
  assign _T_27974 = valid_26_7 ? 6'h7 : _T_27973; // @[Mux.scala 31:69:@8629.4]
  assign _T_27975 = valid_26_6 ? 6'h6 : _T_27974; // @[Mux.scala 31:69:@8630.4]
  assign _T_27976 = valid_26_5 ? 6'h5 : _T_27975; // @[Mux.scala 31:69:@8631.4]
  assign _T_27977 = valid_26_4 ? 6'h4 : _T_27976; // @[Mux.scala 31:69:@8632.4]
  assign _T_27978 = valid_26_3 ? 6'h3 : _T_27977; // @[Mux.scala 31:69:@8633.4]
  assign _T_27979 = valid_26_2 ? 6'h2 : _T_27978; // @[Mux.scala 31:69:@8634.4]
  assign _T_27980 = valid_26_1 ? 6'h1 : _T_27979; // @[Mux.scala 31:69:@8635.4]
  assign select_26 = valid_26_0 ? 6'h0 : _T_27980; // @[Mux.scala 31:69:@8636.4]
  assign _GEN_1665 = 6'h1 == select_26 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1666 = 6'h2 == select_26 ? io_inData_2 : _GEN_1665; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1667 = 6'h3 == select_26 ? io_inData_3 : _GEN_1666; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1668 = 6'h4 == select_26 ? io_inData_4 : _GEN_1667; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1669 = 6'h5 == select_26 ? io_inData_5 : _GEN_1668; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1670 = 6'h6 == select_26 ? io_inData_6 : _GEN_1669; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1671 = 6'h7 == select_26 ? io_inData_7 : _GEN_1670; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1672 = 6'h8 == select_26 ? io_inData_8 : _GEN_1671; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1673 = 6'h9 == select_26 ? io_inData_9 : _GEN_1672; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1674 = 6'ha == select_26 ? io_inData_10 : _GEN_1673; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1675 = 6'hb == select_26 ? io_inData_11 : _GEN_1674; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1676 = 6'hc == select_26 ? io_inData_12 : _GEN_1675; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1677 = 6'hd == select_26 ? io_inData_13 : _GEN_1676; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1678 = 6'he == select_26 ? io_inData_14 : _GEN_1677; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1679 = 6'hf == select_26 ? io_inData_15 : _GEN_1678; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1680 = 6'h10 == select_26 ? io_inData_16 : _GEN_1679; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1681 = 6'h11 == select_26 ? io_inData_17 : _GEN_1680; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1682 = 6'h12 == select_26 ? io_inData_18 : _GEN_1681; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1683 = 6'h13 == select_26 ? io_inData_19 : _GEN_1682; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1684 = 6'h14 == select_26 ? io_inData_20 : _GEN_1683; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1685 = 6'h15 == select_26 ? io_inData_21 : _GEN_1684; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1686 = 6'h16 == select_26 ? io_inData_22 : _GEN_1685; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1687 = 6'h17 == select_26 ? io_inData_23 : _GEN_1686; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1688 = 6'h18 == select_26 ? io_inData_24 : _GEN_1687; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1689 = 6'h19 == select_26 ? io_inData_25 : _GEN_1688; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1690 = 6'h1a == select_26 ? io_inData_26 : _GEN_1689; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1691 = 6'h1b == select_26 ? io_inData_27 : _GEN_1690; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1692 = 6'h1c == select_26 ? io_inData_28 : _GEN_1691; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1693 = 6'h1d == select_26 ? io_inData_29 : _GEN_1692; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1694 = 6'h1e == select_26 ? io_inData_30 : _GEN_1693; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1695 = 6'h1f == select_26 ? io_inData_31 : _GEN_1694; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1696 = 6'h20 == select_26 ? io_inData_32 : _GEN_1695; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1697 = 6'h21 == select_26 ? io_inData_33 : _GEN_1696; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1698 = 6'h22 == select_26 ? io_inData_34 : _GEN_1697; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1699 = 6'h23 == select_26 ? io_inData_35 : _GEN_1698; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1700 = 6'h24 == select_26 ? io_inData_36 : _GEN_1699; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1701 = 6'h25 == select_26 ? io_inData_37 : _GEN_1700; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1702 = 6'h26 == select_26 ? io_inData_38 : _GEN_1701; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1703 = 6'h27 == select_26 ? io_inData_39 : _GEN_1702; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1704 = 6'h28 == select_26 ? io_inData_40 : _GEN_1703; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1705 = 6'h29 == select_26 ? io_inData_41 : _GEN_1704; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1706 = 6'h2a == select_26 ? io_inData_42 : _GEN_1705; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1707 = 6'h2b == select_26 ? io_inData_43 : _GEN_1706; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1708 = 6'h2c == select_26 ? io_inData_44 : _GEN_1707; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1709 = 6'h2d == select_26 ? io_inData_45 : _GEN_1708; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1710 = 6'h2e == select_26 ? io_inData_46 : _GEN_1709; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1711 = 6'h2f == select_26 ? io_inData_47 : _GEN_1710; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1712 = 6'h30 == select_26 ? io_inData_48 : _GEN_1711; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1713 = 6'h31 == select_26 ? io_inData_49 : _GEN_1712; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1714 = 6'h32 == select_26 ? io_inData_50 : _GEN_1713; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1715 = 6'h33 == select_26 ? io_inData_51 : _GEN_1714; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1716 = 6'h34 == select_26 ? io_inData_52 : _GEN_1715; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1717 = 6'h35 == select_26 ? io_inData_53 : _GEN_1716; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1718 = 6'h36 == select_26 ? io_inData_54 : _GEN_1717; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1719 = 6'h37 == select_26 ? io_inData_55 : _GEN_1718; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1720 = 6'h38 == select_26 ? io_inData_56 : _GEN_1719; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1721 = 6'h39 == select_26 ? io_inData_57 : _GEN_1720; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1722 = 6'h3a == select_26 ? io_inData_58 : _GEN_1721; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1723 = 6'h3b == select_26 ? io_inData_59 : _GEN_1722; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1724 = 6'h3c == select_26 ? io_inData_60 : _GEN_1723; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1725 = 6'h3d == select_26 ? io_inData_61 : _GEN_1724; // @[Switch.scala 33:19:@8638.4]
  assign _GEN_1726 = 6'h3e == select_26 ? io_inData_62 : _GEN_1725; // @[Switch.scala 33:19:@8638.4]
  assign _T_27989 = {valid_26_7,valid_26_6,valid_26_5,valid_26_4,valid_26_3,valid_26_2,valid_26_1,valid_26_0}; // @[Switch.scala 34:32:@8645.4]
  assign _T_27997 = {valid_26_15,valid_26_14,valid_26_13,valid_26_12,valid_26_11,valid_26_10,valid_26_9,valid_26_8,_T_27989}; // @[Switch.scala 34:32:@8653.4]
  assign _T_28004 = {valid_26_23,valid_26_22,valid_26_21,valid_26_20,valid_26_19,valid_26_18,valid_26_17,valid_26_16}; // @[Switch.scala 34:32:@8660.4]
  assign _T_28013 = {valid_26_31,valid_26_30,valid_26_29,valid_26_28,valid_26_27,valid_26_26,valid_26_25,valid_26_24,_T_28004,_T_27997}; // @[Switch.scala 34:32:@8669.4]
  assign _T_28020 = {valid_26_39,valid_26_38,valid_26_37,valid_26_36,valid_26_35,valid_26_34,valid_26_33,valid_26_32}; // @[Switch.scala 34:32:@8676.4]
  assign _T_28028 = {valid_26_47,valid_26_46,valid_26_45,valid_26_44,valid_26_43,valid_26_42,valid_26_41,valid_26_40,_T_28020}; // @[Switch.scala 34:32:@8684.4]
  assign _T_28035 = {valid_26_55,valid_26_54,valid_26_53,valid_26_52,valid_26_51,valid_26_50,valid_26_49,valid_26_48}; // @[Switch.scala 34:32:@8691.4]
  assign _T_28044 = {valid_26_63,valid_26_62,valid_26_61,valid_26_60,valid_26_59,valid_26_58,valid_26_57,valid_26_56,_T_28035,_T_28028}; // @[Switch.scala 34:32:@8700.4]
  assign _T_28045 = {_T_28044,_T_28013}; // @[Switch.scala 34:32:@8701.4]
  assign _T_28049 = io_inAddr_0 == 6'h1b; // @[Switch.scala 30:53:@8704.4]
  assign valid_27_0 = io_inValid_0 & _T_28049; // @[Switch.scala 30:36:@8705.4]
  assign _T_28052 = io_inAddr_1 == 6'h1b; // @[Switch.scala 30:53:@8707.4]
  assign valid_27_1 = io_inValid_1 & _T_28052; // @[Switch.scala 30:36:@8708.4]
  assign _T_28055 = io_inAddr_2 == 6'h1b; // @[Switch.scala 30:53:@8710.4]
  assign valid_27_2 = io_inValid_2 & _T_28055; // @[Switch.scala 30:36:@8711.4]
  assign _T_28058 = io_inAddr_3 == 6'h1b; // @[Switch.scala 30:53:@8713.4]
  assign valid_27_3 = io_inValid_3 & _T_28058; // @[Switch.scala 30:36:@8714.4]
  assign _T_28061 = io_inAddr_4 == 6'h1b; // @[Switch.scala 30:53:@8716.4]
  assign valid_27_4 = io_inValid_4 & _T_28061; // @[Switch.scala 30:36:@8717.4]
  assign _T_28064 = io_inAddr_5 == 6'h1b; // @[Switch.scala 30:53:@8719.4]
  assign valid_27_5 = io_inValid_5 & _T_28064; // @[Switch.scala 30:36:@8720.4]
  assign _T_28067 = io_inAddr_6 == 6'h1b; // @[Switch.scala 30:53:@8722.4]
  assign valid_27_6 = io_inValid_6 & _T_28067; // @[Switch.scala 30:36:@8723.4]
  assign _T_28070 = io_inAddr_7 == 6'h1b; // @[Switch.scala 30:53:@8725.4]
  assign valid_27_7 = io_inValid_7 & _T_28070; // @[Switch.scala 30:36:@8726.4]
  assign _T_28073 = io_inAddr_8 == 6'h1b; // @[Switch.scala 30:53:@8728.4]
  assign valid_27_8 = io_inValid_8 & _T_28073; // @[Switch.scala 30:36:@8729.4]
  assign _T_28076 = io_inAddr_9 == 6'h1b; // @[Switch.scala 30:53:@8731.4]
  assign valid_27_9 = io_inValid_9 & _T_28076; // @[Switch.scala 30:36:@8732.4]
  assign _T_28079 = io_inAddr_10 == 6'h1b; // @[Switch.scala 30:53:@8734.4]
  assign valid_27_10 = io_inValid_10 & _T_28079; // @[Switch.scala 30:36:@8735.4]
  assign _T_28082 = io_inAddr_11 == 6'h1b; // @[Switch.scala 30:53:@8737.4]
  assign valid_27_11 = io_inValid_11 & _T_28082; // @[Switch.scala 30:36:@8738.4]
  assign _T_28085 = io_inAddr_12 == 6'h1b; // @[Switch.scala 30:53:@8740.4]
  assign valid_27_12 = io_inValid_12 & _T_28085; // @[Switch.scala 30:36:@8741.4]
  assign _T_28088 = io_inAddr_13 == 6'h1b; // @[Switch.scala 30:53:@8743.4]
  assign valid_27_13 = io_inValid_13 & _T_28088; // @[Switch.scala 30:36:@8744.4]
  assign _T_28091 = io_inAddr_14 == 6'h1b; // @[Switch.scala 30:53:@8746.4]
  assign valid_27_14 = io_inValid_14 & _T_28091; // @[Switch.scala 30:36:@8747.4]
  assign _T_28094 = io_inAddr_15 == 6'h1b; // @[Switch.scala 30:53:@8749.4]
  assign valid_27_15 = io_inValid_15 & _T_28094; // @[Switch.scala 30:36:@8750.4]
  assign _T_28097 = io_inAddr_16 == 6'h1b; // @[Switch.scala 30:53:@8752.4]
  assign valid_27_16 = io_inValid_16 & _T_28097; // @[Switch.scala 30:36:@8753.4]
  assign _T_28100 = io_inAddr_17 == 6'h1b; // @[Switch.scala 30:53:@8755.4]
  assign valid_27_17 = io_inValid_17 & _T_28100; // @[Switch.scala 30:36:@8756.4]
  assign _T_28103 = io_inAddr_18 == 6'h1b; // @[Switch.scala 30:53:@8758.4]
  assign valid_27_18 = io_inValid_18 & _T_28103; // @[Switch.scala 30:36:@8759.4]
  assign _T_28106 = io_inAddr_19 == 6'h1b; // @[Switch.scala 30:53:@8761.4]
  assign valid_27_19 = io_inValid_19 & _T_28106; // @[Switch.scala 30:36:@8762.4]
  assign _T_28109 = io_inAddr_20 == 6'h1b; // @[Switch.scala 30:53:@8764.4]
  assign valid_27_20 = io_inValid_20 & _T_28109; // @[Switch.scala 30:36:@8765.4]
  assign _T_28112 = io_inAddr_21 == 6'h1b; // @[Switch.scala 30:53:@8767.4]
  assign valid_27_21 = io_inValid_21 & _T_28112; // @[Switch.scala 30:36:@8768.4]
  assign _T_28115 = io_inAddr_22 == 6'h1b; // @[Switch.scala 30:53:@8770.4]
  assign valid_27_22 = io_inValid_22 & _T_28115; // @[Switch.scala 30:36:@8771.4]
  assign _T_28118 = io_inAddr_23 == 6'h1b; // @[Switch.scala 30:53:@8773.4]
  assign valid_27_23 = io_inValid_23 & _T_28118; // @[Switch.scala 30:36:@8774.4]
  assign _T_28121 = io_inAddr_24 == 6'h1b; // @[Switch.scala 30:53:@8776.4]
  assign valid_27_24 = io_inValid_24 & _T_28121; // @[Switch.scala 30:36:@8777.4]
  assign _T_28124 = io_inAddr_25 == 6'h1b; // @[Switch.scala 30:53:@8779.4]
  assign valid_27_25 = io_inValid_25 & _T_28124; // @[Switch.scala 30:36:@8780.4]
  assign _T_28127 = io_inAddr_26 == 6'h1b; // @[Switch.scala 30:53:@8782.4]
  assign valid_27_26 = io_inValid_26 & _T_28127; // @[Switch.scala 30:36:@8783.4]
  assign _T_28130 = io_inAddr_27 == 6'h1b; // @[Switch.scala 30:53:@8785.4]
  assign valid_27_27 = io_inValid_27 & _T_28130; // @[Switch.scala 30:36:@8786.4]
  assign _T_28133 = io_inAddr_28 == 6'h1b; // @[Switch.scala 30:53:@8788.4]
  assign valid_27_28 = io_inValid_28 & _T_28133; // @[Switch.scala 30:36:@8789.4]
  assign _T_28136 = io_inAddr_29 == 6'h1b; // @[Switch.scala 30:53:@8791.4]
  assign valid_27_29 = io_inValid_29 & _T_28136; // @[Switch.scala 30:36:@8792.4]
  assign _T_28139 = io_inAddr_30 == 6'h1b; // @[Switch.scala 30:53:@8794.4]
  assign valid_27_30 = io_inValid_30 & _T_28139; // @[Switch.scala 30:36:@8795.4]
  assign _T_28142 = io_inAddr_31 == 6'h1b; // @[Switch.scala 30:53:@8797.4]
  assign valid_27_31 = io_inValid_31 & _T_28142; // @[Switch.scala 30:36:@8798.4]
  assign _T_28145 = io_inAddr_32 == 6'h1b; // @[Switch.scala 30:53:@8800.4]
  assign valid_27_32 = io_inValid_32 & _T_28145; // @[Switch.scala 30:36:@8801.4]
  assign _T_28148 = io_inAddr_33 == 6'h1b; // @[Switch.scala 30:53:@8803.4]
  assign valid_27_33 = io_inValid_33 & _T_28148; // @[Switch.scala 30:36:@8804.4]
  assign _T_28151 = io_inAddr_34 == 6'h1b; // @[Switch.scala 30:53:@8806.4]
  assign valid_27_34 = io_inValid_34 & _T_28151; // @[Switch.scala 30:36:@8807.4]
  assign _T_28154 = io_inAddr_35 == 6'h1b; // @[Switch.scala 30:53:@8809.4]
  assign valid_27_35 = io_inValid_35 & _T_28154; // @[Switch.scala 30:36:@8810.4]
  assign _T_28157 = io_inAddr_36 == 6'h1b; // @[Switch.scala 30:53:@8812.4]
  assign valid_27_36 = io_inValid_36 & _T_28157; // @[Switch.scala 30:36:@8813.4]
  assign _T_28160 = io_inAddr_37 == 6'h1b; // @[Switch.scala 30:53:@8815.4]
  assign valid_27_37 = io_inValid_37 & _T_28160; // @[Switch.scala 30:36:@8816.4]
  assign _T_28163 = io_inAddr_38 == 6'h1b; // @[Switch.scala 30:53:@8818.4]
  assign valid_27_38 = io_inValid_38 & _T_28163; // @[Switch.scala 30:36:@8819.4]
  assign _T_28166 = io_inAddr_39 == 6'h1b; // @[Switch.scala 30:53:@8821.4]
  assign valid_27_39 = io_inValid_39 & _T_28166; // @[Switch.scala 30:36:@8822.4]
  assign _T_28169 = io_inAddr_40 == 6'h1b; // @[Switch.scala 30:53:@8824.4]
  assign valid_27_40 = io_inValid_40 & _T_28169; // @[Switch.scala 30:36:@8825.4]
  assign _T_28172 = io_inAddr_41 == 6'h1b; // @[Switch.scala 30:53:@8827.4]
  assign valid_27_41 = io_inValid_41 & _T_28172; // @[Switch.scala 30:36:@8828.4]
  assign _T_28175 = io_inAddr_42 == 6'h1b; // @[Switch.scala 30:53:@8830.4]
  assign valid_27_42 = io_inValid_42 & _T_28175; // @[Switch.scala 30:36:@8831.4]
  assign _T_28178 = io_inAddr_43 == 6'h1b; // @[Switch.scala 30:53:@8833.4]
  assign valid_27_43 = io_inValid_43 & _T_28178; // @[Switch.scala 30:36:@8834.4]
  assign _T_28181 = io_inAddr_44 == 6'h1b; // @[Switch.scala 30:53:@8836.4]
  assign valid_27_44 = io_inValid_44 & _T_28181; // @[Switch.scala 30:36:@8837.4]
  assign _T_28184 = io_inAddr_45 == 6'h1b; // @[Switch.scala 30:53:@8839.4]
  assign valid_27_45 = io_inValid_45 & _T_28184; // @[Switch.scala 30:36:@8840.4]
  assign _T_28187 = io_inAddr_46 == 6'h1b; // @[Switch.scala 30:53:@8842.4]
  assign valid_27_46 = io_inValid_46 & _T_28187; // @[Switch.scala 30:36:@8843.4]
  assign _T_28190 = io_inAddr_47 == 6'h1b; // @[Switch.scala 30:53:@8845.4]
  assign valid_27_47 = io_inValid_47 & _T_28190; // @[Switch.scala 30:36:@8846.4]
  assign _T_28193 = io_inAddr_48 == 6'h1b; // @[Switch.scala 30:53:@8848.4]
  assign valid_27_48 = io_inValid_48 & _T_28193; // @[Switch.scala 30:36:@8849.4]
  assign _T_28196 = io_inAddr_49 == 6'h1b; // @[Switch.scala 30:53:@8851.4]
  assign valid_27_49 = io_inValid_49 & _T_28196; // @[Switch.scala 30:36:@8852.4]
  assign _T_28199 = io_inAddr_50 == 6'h1b; // @[Switch.scala 30:53:@8854.4]
  assign valid_27_50 = io_inValid_50 & _T_28199; // @[Switch.scala 30:36:@8855.4]
  assign _T_28202 = io_inAddr_51 == 6'h1b; // @[Switch.scala 30:53:@8857.4]
  assign valid_27_51 = io_inValid_51 & _T_28202; // @[Switch.scala 30:36:@8858.4]
  assign _T_28205 = io_inAddr_52 == 6'h1b; // @[Switch.scala 30:53:@8860.4]
  assign valid_27_52 = io_inValid_52 & _T_28205; // @[Switch.scala 30:36:@8861.4]
  assign _T_28208 = io_inAddr_53 == 6'h1b; // @[Switch.scala 30:53:@8863.4]
  assign valid_27_53 = io_inValid_53 & _T_28208; // @[Switch.scala 30:36:@8864.4]
  assign _T_28211 = io_inAddr_54 == 6'h1b; // @[Switch.scala 30:53:@8866.4]
  assign valid_27_54 = io_inValid_54 & _T_28211; // @[Switch.scala 30:36:@8867.4]
  assign _T_28214 = io_inAddr_55 == 6'h1b; // @[Switch.scala 30:53:@8869.4]
  assign valid_27_55 = io_inValid_55 & _T_28214; // @[Switch.scala 30:36:@8870.4]
  assign _T_28217 = io_inAddr_56 == 6'h1b; // @[Switch.scala 30:53:@8872.4]
  assign valid_27_56 = io_inValid_56 & _T_28217; // @[Switch.scala 30:36:@8873.4]
  assign _T_28220 = io_inAddr_57 == 6'h1b; // @[Switch.scala 30:53:@8875.4]
  assign valid_27_57 = io_inValid_57 & _T_28220; // @[Switch.scala 30:36:@8876.4]
  assign _T_28223 = io_inAddr_58 == 6'h1b; // @[Switch.scala 30:53:@8878.4]
  assign valid_27_58 = io_inValid_58 & _T_28223; // @[Switch.scala 30:36:@8879.4]
  assign _T_28226 = io_inAddr_59 == 6'h1b; // @[Switch.scala 30:53:@8881.4]
  assign valid_27_59 = io_inValid_59 & _T_28226; // @[Switch.scala 30:36:@8882.4]
  assign _T_28229 = io_inAddr_60 == 6'h1b; // @[Switch.scala 30:53:@8884.4]
  assign valid_27_60 = io_inValid_60 & _T_28229; // @[Switch.scala 30:36:@8885.4]
  assign _T_28232 = io_inAddr_61 == 6'h1b; // @[Switch.scala 30:53:@8887.4]
  assign valid_27_61 = io_inValid_61 & _T_28232; // @[Switch.scala 30:36:@8888.4]
  assign _T_28235 = io_inAddr_62 == 6'h1b; // @[Switch.scala 30:53:@8890.4]
  assign valid_27_62 = io_inValid_62 & _T_28235; // @[Switch.scala 30:36:@8891.4]
  assign _T_28238 = io_inAddr_63 == 6'h1b; // @[Switch.scala 30:53:@8893.4]
  assign valid_27_63 = io_inValid_63 & _T_28238; // @[Switch.scala 30:36:@8894.4]
  assign _T_28304 = valid_27_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@8896.4]
  assign _T_28305 = valid_27_61 ? 6'h3d : _T_28304; // @[Mux.scala 31:69:@8897.4]
  assign _T_28306 = valid_27_60 ? 6'h3c : _T_28305; // @[Mux.scala 31:69:@8898.4]
  assign _T_28307 = valid_27_59 ? 6'h3b : _T_28306; // @[Mux.scala 31:69:@8899.4]
  assign _T_28308 = valid_27_58 ? 6'h3a : _T_28307; // @[Mux.scala 31:69:@8900.4]
  assign _T_28309 = valid_27_57 ? 6'h39 : _T_28308; // @[Mux.scala 31:69:@8901.4]
  assign _T_28310 = valid_27_56 ? 6'h38 : _T_28309; // @[Mux.scala 31:69:@8902.4]
  assign _T_28311 = valid_27_55 ? 6'h37 : _T_28310; // @[Mux.scala 31:69:@8903.4]
  assign _T_28312 = valid_27_54 ? 6'h36 : _T_28311; // @[Mux.scala 31:69:@8904.4]
  assign _T_28313 = valid_27_53 ? 6'h35 : _T_28312; // @[Mux.scala 31:69:@8905.4]
  assign _T_28314 = valid_27_52 ? 6'h34 : _T_28313; // @[Mux.scala 31:69:@8906.4]
  assign _T_28315 = valid_27_51 ? 6'h33 : _T_28314; // @[Mux.scala 31:69:@8907.4]
  assign _T_28316 = valid_27_50 ? 6'h32 : _T_28315; // @[Mux.scala 31:69:@8908.4]
  assign _T_28317 = valid_27_49 ? 6'h31 : _T_28316; // @[Mux.scala 31:69:@8909.4]
  assign _T_28318 = valid_27_48 ? 6'h30 : _T_28317; // @[Mux.scala 31:69:@8910.4]
  assign _T_28319 = valid_27_47 ? 6'h2f : _T_28318; // @[Mux.scala 31:69:@8911.4]
  assign _T_28320 = valid_27_46 ? 6'h2e : _T_28319; // @[Mux.scala 31:69:@8912.4]
  assign _T_28321 = valid_27_45 ? 6'h2d : _T_28320; // @[Mux.scala 31:69:@8913.4]
  assign _T_28322 = valid_27_44 ? 6'h2c : _T_28321; // @[Mux.scala 31:69:@8914.4]
  assign _T_28323 = valid_27_43 ? 6'h2b : _T_28322; // @[Mux.scala 31:69:@8915.4]
  assign _T_28324 = valid_27_42 ? 6'h2a : _T_28323; // @[Mux.scala 31:69:@8916.4]
  assign _T_28325 = valid_27_41 ? 6'h29 : _T_28324; // @[Mux.scala 31:69:@8917.4]
  assign _T_28326 = valid_27_40 ? 6'h28 : _T_28325; // @[Mux.scala 31:69:@8918.4]
  assign _T_28327 = valid_27_39 ? 6'h27 : _T_28326; // @[Mux.scala 31:69:@8919.4]
  assign _T_28328 = valid_27_38 ? 6'h26 : _T_28327; // @[Mux.scala 31:69:@8920.4]
  assign _T_28329 = valid_27_37 ? 6'h25 : _T_28328; // @[Mux.scala 31:69:@8921.4]
  assign _T_28330 = valid_27_36 ? 6'h24 : _T_28329; // @[Mux.scala 31:69:@8922.4]
  assign _T_28331 = valid_27_35 ? 6'h23 : _T_28330; // @[Mux.scala 31:69:@8923.4]
  assign _T_28332 = valid_27_34 ? 6'h22 : _T_28331; // @[Mux.scala 31:69:@8924.4]
  assign _T_28333 = valid_27_33 ? 6'h21 : _T_28332; // @[Mux.scala 31:69:@8925.4]
  assign _T_28334 = valid_27_32 ? 6'h20 : _T_28333; // @[Mux.scala 31:69:@8926.4]
  assign _T_28335 = valid_27_31 ? 6'h1f : _T_28334; // @[Mux.scala 31:69:@8927.4]
  assign _T_28336 = valid_27_30 ? 6'h1e : _T_28335; // @[Mux.scala 31:69:@8928.4]
  assign _T_28337 = valid_27_29 ? 6'h1d : _T_28336; // @[Mux.scala 31:69:@8929.4]
  assign _T_28338 = valid_27_28 ? 6'h1c : _T_28337; // @[Mux.scala 31:69:@8930.4]
  assign _T_28339 = valid_27_27 ? 6'h1b : _T_28338; // @[Mux.scala 31:69:@8931.4]
  assign _T_28340 = valid_27_26 ? 6'h1a : _T_28339; // @[Mux.scala 31:69:@8932.4]
  assign _T_28341 = valid_27_25 ? 6'h19 : _T_28340; // @[Mux.scala 31:69:@8933.4]
  assign _T_28342 = valid_27_24 ? 6'h18 : _T_28341; // @[Mux.scala 31:69:@8934.4]
  assign _T_28343 = valid_27_23 ? 6'h17 : _T_28342; // @[Mux.scala 31:69:@8935.4]
  assign _T_28344 = valid_27_22 ? 6'h16 : _T_28343; // @[Mux.scala 31:69:@8936.4]
  assign _T_28345 = valid_27_21 ? 6'h15 : _T_28344; // @[Mux.scala 31:69:@8937.4]
  assign _T_28346 = valid_27_20 ? 6'h14 : _T_28345; // @[Mux.scala 31:69:@8938.4]
  assign _T_28347 = valid_27_19 ? 6'h13 : _T_28346; // @[Mux.scala 31:69:@8939.4]
  assign _T_28348 = valid_27_18 ? 6'h12 : _T_28347; // @[Mux.scala 31:69:@8940.4]
  assign _T_28349 = valid_27_17 ? 6'h11 : _T_28348; // @[Mux.scala 31:69:@8941.4]
  assign _T_28350 = valid_27_16 ? 6'h10 : _T_28349; // @[Mux.scala 31:69:@8942.4]
  assign _T_28351 = valid_27_15 ? 6'hf : _T_28350; // @[Mux.scala 31:69:@8943.4]
  assign _T_28352 = valid_27_14 ? 6'he : _T_28351; // @[Mux.scala 31:69:@8944.4]
  assign _T_28353 = valid_27_13 ? 6'hd : _T_28352; // @[Mux.scala 31:69:@8945.4]
  assign _T_28354 = valid_27_12 ? 6'hc : _T_28353; // @[Mux.scala 31:69:@8946.4]
  assign _T_28355 = valid_27_11 ? 6'hb : _T_28354; // @[Mux.scala 31:69:@8947.4]
  assign _T_28356 = valid_27_10 ? 6'ha : _T_28355; // @[Mux.scala 31:69:@8948.4]
  assign _T_28357 = valid_27_9 ? 6'h9 : _T_28356; // @[Mux.scala 31:69:@8949.4]
  assign _T_28358 = valid_27_8 ? 6'h8 : _T_28357; // @[Mux.scala 31:69:@8950.4]
  assign _T_28359 = valid_27_7 ? 6'h7 : _T_28358; // @[Mux.scala 31:69:@8951.4]
  assign _T_28360 = valid_27_6 ? 6'h6 : _T_28359; // @[Mux.scala 31:69:@8952.4]
  assign _T_28361 = valid_27_5 ? 6'h5 : _T_28360; // @[Mux.scala 31:69:@8953.4]
  assign _T_28362 = valid_27_4 ? 6'h4 : _T_28361; // @[Mux.scala 31:69:@8954.4]
  assign _T_28363 = valid_27_3 ? 6'h3 : _T_28362; // @[Mux.scala 31:69:@8955.4]
  assign _T_28364 = valid_27_2 ? 6'h2 : _T_28363; // @[Mux.scala 31:69:@8956.4]
  assign _T_28365 = valid_27_1 ? 6'h1 : _T_28364; // @[Mux.scala 31:69:@8957.4]
  assign select_27 = valid_27_0 ? 6'h0 : _T_28365; // @[Mux.scala 31:69:@8958.4]
  assign _GEN_1729 = 6'h1 == select_27 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1730 = 6'h2 == select_27 ? io_inData_2 : _GEN_1729; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1731 = 6'h3 == select_27 ? io_inData_3 : _GEN_1730; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1732 = 6'h4 == select_27 ? io_inData_4 : _GEN_1731; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1733 = 6'h5 == select_27 ? io_inData_5 : _GEN_1732; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1734 = 6'h6 == select_27 ? io_inData_6 : _GEN_1733; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1735 = 6'h7 == select_27 ? io_inData_7 : _GEN_1734; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1736 = 6'h8 == select_27 ? io_inData_8 : _GEN_1735; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1737 = 6'h9 == select_27 ? io_inData_9 : _GEN_1736; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1738 = 6'ha == select_27 ? io_inData_10 : _GEN_1737; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1739 = 6'hb == select_27 ? io_inData_11 : _GEN_1738; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1740 = 6'hc == select_27 ? io_inData_12 : _GEN_1739; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1741 = 6'hd == select_27 ? io_inData_13 : _GEN_1740; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1742 = 6'he == select_27 ? io_inData_14 : _GEN_1741; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1743 = 6'hf == select_27 ? io_inData_15 : _GEN_1742; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1744 = 6'h10 == select_27 ? io_inData_16 : _GEN_1743; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1745 = 6'h11 == select_27 ? io_inData_17 : _GEN_1744; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1746 = 6'h12 == select_27 ? io_inData_18 : _GEN_1745; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1747 = 6'h13 == select_27 ? io_inData_19 : _GEN_1746; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1748 = 6'h14 == select_27 ? io_inData_20 : _GEN_1747; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1749 = 6'h15 == select_27 ? io_inData_21 : _GEN_1748; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1750 = 6'h16 == select_27 ? io_inData_22 : _GEN_1749; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1751 = 6'h17 == select_27 ? io_inData_23 : _GEN_1750; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1752 = 6'h18 == select_27 ? io_inData_24 : _GEN_1751; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1753 = 6'h19 == select_27 ? io_inData_25 : _GEN_1752; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1754 = 6'h1a == select_27 ? io_inData_26 : _GEN_1753; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1755 = 6'h1b == select_27 ? io_inData_27 : _GEN_1754; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1756 = 6'h1c == select_27 ? io_inData_28 : _GEN_1755; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1757 = 6'h1d == select_27 ? io_inData_29 : _GEN_1756; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1758 = 6'h1e == select_27 ? io_inData_30 : _GEN_1757; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1759 = 6'h1f == select_27 ? io_inData_31 : _GEN_1758; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1760 = 6'h20 == select_27 ? io_inData_32 : _GEN_1759; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1761 = 6'h21 == select_27 ? io_inData_33 : _GEN_1760; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1762 = 6'h22 == select_27 ? io_inData_34 : _GEN_1761; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1763 = 6'h23 == select_27 ? io_inData_35 : _GEN_1762; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1764 = 6'h24 == select_27 ? io_inData_36 : _GEN_1763; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1765 = 6'h25 == select_27 ? io_inData_37 : _GEN_1764; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1766 = 6'h26 == select_27 ? io_inData_38 : _GEN_1765; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1767 = 6'h27 == select_27 ? io_inData_39 : _GEN_1766; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1768 = 6'h28 == select_27 ? io_inData_40 : _GEN_1767; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1769 = 6'h29 == select_27 ? io_inData_41 : _GEN_1768; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1770 = 6'h2a == select_27 ? io_inData_42 : _GEN_1769; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1771 = 6'h2b == select_27 ? io_inData_43 : _GEN_1770; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1772 = 6'h2c == select_27 ? io_inData_44 : _GEN_1771; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1773 = 6'h2d == select_27 ? io_inData_45 : _GEN_1772; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1774 = 6'h2e == select_27 ? io_inData_46 : _GEN_1773; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1775 = 6'h2f == select_27 ? io_inData_47 : _GEN_1774; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1776 = 6'h30 == select_27 ? io_inData_48 : _GEN_1775; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1777 = 6'h31 == select_27 ? io_inData_49 : _GEN_1776; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1778 = 6'h32 == select_27 ? io_inData_50 : _GEN_1777; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1779 = 6'h33 == select_27 ? io_inData_51 : _GEN_1778; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1780 = 6'h34 == select_27 ? io_inData_52 : _GEN_1779; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1781 = 6'h35 == select_27 ? io_inData_53 : _GEN_1780; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1782 = 6'h36 == select_27 ? io_inData_54 : _GEN_1781; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1783 = 6'h37 == select_27 ? io_inData_55 : _GEN_1782; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1784 = 6'h38 == select_27 ? io_inData_56 : _GEN_1783; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1785 = 6'h39 == select_27 ? io_inData_57 : _GEN_1784; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1786 = 6'h3a == select_27 ? io_inData_58 : _GEN_1785; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1787 = 6'h3b == select_27 ? io_inData_59 : _GEN_1786; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1788 = 6'h3c == select_27 ? io_inData_60 : _GEN_1787; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1789 = 6'h3d == select_27 ? io_inData_61 : _GEN_1788; // @[Switch.scala 33:19:@8960.4]
  assign _GEN_1790 = 6'h3e == select_27 ? io_inData_62 : _GEN_1789; // @[Switch.scala 33:19:@8960.4]
  assign _T_28374 = {valid_27_7,valid_27_6,valid_27_5,valid_27_4,valid_27_3,valid_27_2,valid_27_1,valid_27_0}; // @[Switch.scala 34:32:@8967.4]
  assign _T_28382 = {valid_27_15,valid_27_14,valid_27_13,valid_27_12,valid_27_11,valid_27_10,valid_27_9,valid_27_8,_T_28374}; // @[Switch.scala 34:32:@8975.4]
  assign _T_28389 = {valid_27_23,valid_27_22,valid_27_21,valid_27_20,valid_27_19,valid_27_18,valid_27_17,valid_27_16}; // @[Switch.scala 34:32:@8982.4]
  assign _T_28398 = {valid_27_31,valid_27_30,valid_27_29,valid_27_28,valid_27_27,valid_27_26,valid_27_25,valid_27_24,_T_28389,_T_28382}; // @[Switch.scala 34:32:@8991.4]
  assign _T_28405 = {valid_27_39,valid_27_38,valid_27_37,valid_27_36,valid_27_35,valid_27_34,valid_27_33,valid_27_32}; // @[Switch.scala 34:32:@8998.4]
  assign _T_28413 = {valid_27_47,valid_27_46,valid_27_45,valid_27_44,valid_27_43,valid_27_42,valid_27_41,valid_27_40,_T_28405}; // @[Switch.scala 34:32:@9006.4]
  assign _T_28420 = {valid_27_55,valid_27_54,valid_27_53,valid_27_52,valid_27_51,valid_27_50,valid_27_49,valid_27_48}; // @[Switch.scala 34:32:@9013.4]
  assign _T_28429 = {valid_27_63,valid_27_62,valid_27_61,valid_27_60,valid_27_59,valid_27_58,valid_27_57,valid_27_56,_T_28420,_T_28413}; // @[Switch.scala 34:32:@9022.4]
  assign _T_28430 = {_T_28429,_T_28398}; // @[Switch.scala 34:32:@9023.4]
  assign _T_28434 = io_inAddr_0 == 6'h1c; // @[Switch.scala 30:53:@9026.4]
  assign valid_28_0 = io_inValid_0 & _T_28434; // @[Switch.scala 30:36:@9027.4]
  assign _T_28437 = io_inAddr_1 == 6'h1c; // @[Switch.scala 30:53:@9029.4]
  assign valid_28_1 = io_inValid_1 & _T_28437; // @[Switch.scala 30:36:@9030.4]
  assign _T_28440 = io_inAddr_2 == 6'h1c; // @[Switch.scala 30:53:@9032.4]
  assign valid_28_2 = io_inValid_2 & _T_28440; // @[Switch.scala 30:36:@9033.4]
  assign _T_28443 = io_inAddr_3 == 6'h1c; // @[Switch.scala 30:53:@9035.4]
  assign valid_28_3 = io_inValid_3 & _T_28443; // @[Switch.scala 30:36:@9036.4]
  assign _T_28446 = io_inAddr_4 == 6'h1c; // @[Switch.scala 30:53:@9038.4]
  assign valid_28_4 = io_inValid_4 & _T_28446; // @[Switch.scala 30:36:@9039.4]
  assign _T_28449 = io_inAddr_5 == 6'h1c; // @[Switch.scala 30:53:@9041.4]
  assign valid_28_5 = io_inValid_5 & _T_28449; // @[Switch.scala 30:36:@9042.4]
  assign _T_28452 = io_inAddr_6 == 6'h1c; // @[Switch.scala 30:53:@9044.4]
  assign valid_28_6 = io_inValid_6 & _T_28452; // @[Switch.scala 30:36:@9045.4]
  assign _T_28455 = io_inAddr_7 == 6'h1c; // @[Switch.scala 30:53:@9047.4]
  assign valid_28_7 = io_inValid_7 & _T_28455; // @[Switch.scala 30:36:@9048.4]
  assign _T_28458 = io_inAddr_8 == 6'h1c; // @[Switch.scala 30:53:@9050.4]
  assign valid_28_8 = io_inValid_8 & _T_28458; // @[Switch.scala 30:36:@9051.4]
  assign _T_28461 = io_inAddr_9 == 6'h1c; // @[Switch.scala 30:53:@9053.4]
  assign valid_28_9 = io_inValid_9 & _T_28461; // @[Switch.scala 30:36:@9054.4]
  assign _T_28464 = io_inAddr_10 == 6'h1c; // @[Switch.scala 30:53:@9056.4]
  assign valid_28_10 = io_inValid_10 & _T_28464; // @[Switch.scala 30:36:@9057.4]
  assign _T_28467 = io_inAddr_11 == 6'h1c; // @[Switch.scala 30:53:@9059.4]
  assign valid_28_11 = io_inValid_11 & _T_28467; // @[Switch.scala 30:36:@9060.4]
  assign _T_28470 = io_inAddr_12 == 6'h1c; // @[Switch.scala 30:53:@9062.4]
  assign valid_28_12 = io_inValid_12 & _T_28470; // @[Switch.scala 30:36:@9063.4]
  assign _T_28473 = io_inAddr_13 == 6'h1c; // @[Switch.scala 30:53:@9065.4]
  assign valid_28_13 = io_inValid_13 & _T_28473; // @[Switch.scala 30:36:@9066.4]
  assign _T_28476 = io_inAddr_14 == 6'h1c; // @[Switch.scala 30:53:@9068.4]
  assign valid_28_14 = io_inValid_14 & _T_28476; // @[Switch.scala 30:36:@9069.4]
  assign _T_28479 = io_inAddr_15 == 6'h1c; // @[Switch.scala 30:53:@9071.4]
  assign valid_28_15 = io_inValid_15 & _T_28479; // @[Switch.scala 30:36:@9072.4]
  assign _T_28482 = io_inAddr_16 == 6'h1c; // @[Switch.scala 30:53:@9074.4]
  assign valid_28_16 = io_inValid_16 & _T_28482; // @[Switch.scala 30:36:@9075.4]
  assign _T_28485 = io_inAddr_17 == 6'h1c; // @[Switch.scala 30:53:@9077.4]
  assign valid_28_17 = io_inValid_17 & _T_28485; // @[Switch.scala 30:36:@9078.4]
  assign _T_28488 = io_inAddr_18 == 6'h1c; // @[Switch.scala 30:53:@9080.4]
  assign valid_28_18 = io_inValid_18 & _T_28488; // @[Switch.scala 30:36:@9081.4]
  assign _T_28491 = io_inAddr_19 == 6'h1c; // @[Switch.scala 30:53:@9083.4]
  assign valid_28_19 = io_inValid_19 & _T_28491; // @[Switch.scala 30:36:@9084.4]
  assign _T_28494 = io_inAddr_20 == 6'h1c; // @[Switch.scala 30:53:@9086.4]
  assign valid_28_20 = io_inValid_20 & _T_28494; // @[Switch.scala 30:36:@9087.4]
  assign _T_28497 = io_inAddr_21 == 6'h1c; // @[Switch.scala 30:53:@9089.4]
  assign valid_28_21 = io_inValid_21 & _T_28497; // @[Switch.scala 30:36:@9090.4]
  assign _T_28500 = io_inAddr_22 == 6'h1c; // @[Switch.scala 30:53:@9092.4]
  assign valid_28_22 = io_inValid_22 & _T_28500; // @[Switch.scala 30:36:@9093.4]
  assign _T_28503 = io_inAddr_23 == 6'h1c; // @[Switch.scala 30:53:@9095.4]
  assign valid_28_23 = io_inValid_23 & _T_28503; // @[Switch.scala 30:36:@9096.4]
  assign _T_28506 = io_inAddr_24 == 6'h1c; // @[Switch.scala 30:53:@9098.4]
  assign valid_28_24 = io_inValid_24 & _T_28506; // @[Switch.scala 30:36:@9099.4]
  assign _T_28509 = io_inAddr_25 == 6'h1c; // @[Switch.scala 30:53:@9101.4]
  assign valid_28_25 = io_inValid_25 & _T_28509; // @[Switch.scala 30:36:@9102.4]
  assign _T_28512 = io_inAddr_26 == 6'h1c; // @[Switch.scala 30:53:@9104.4]
  assign valid_28_26 = io_inValid_26 & _T_28512; // @[Switch.scala 30:36:@9105.4]
  assign _T_28515 = io_inAddr_27 == 6'h1c; // @[Switch.scala 30:53:@9107.4]
  assign valid_28_27 = io_inValid_27 & _T_28515; // @[Switch.scala 30:36:@9108.4]
  assign _T_28518 = io_inAddr_28 == 6'h1c; // @[Switch.scala 30:53:@9110.4]
  assign valid_28_28 = io_inValid_28 & _T_28518; // @[Switch.scala 30:36:@9111.4]
  assign _T_28521 = io_inAddr_29 == 6'h1c; // @[Switch.scala 30:53:@9113.4]
  assign valid_28_29 = io_inValid_29 & _T_28521; // @[Switch.scala 30:36:@9114.4]
  assign _T_28524 = io_inAddr_30 == 6'h1c; // @[Switch.scala 30:53:@9116.4]
  assign valid_28_30 = io_inValid_30 & _T_28524; // @[Switch.scala 30:36:@9117.4]
  assign _T_28527 = io_inAddr_31 == 6'h1c; // @[Switch.scala 30:53:@9119.4]
  assign valid_28_31 = io_inValid_31 & _T_28527; // @[Switch.scala 30:36:@9120.4]
  assign _T_28530 = io_inAddr_32 == 6'h1c; // @[Switch.scala 30:53:@9122.4]
  assign valid_28_32 = io_inValid_32 & _T_28530; // @[Switch.scala 30:36:@9123.4]
  assign _T_28533 = io_inAddr_33 == 6'h1c; // @[Switch.scala 30:53:@9125.4]
  assign valid_28_33 = io_inValid_33 & _T_28533; // @[Switch.scala 30:36:@9126.4]
  assign _T_28536 = io_inAddr_34 == 6'h1c; // @[Switch.scala 30:53:@9128.4]
  assign valid_28_34 = io_inValid_34 & _T_28536; // @[Switch.scala 30:36:@9129.4]
  assign _T_28539 = io_inAddr_35 == 6'h1c; // @[Switch.scala 30:53:@9131.4]
  assign valid_28_35 = io_inValid_35 & _T_28539; // @[Switch.scala 30:36:@9132.4]
  assign _T_28542 = io_inAddr_36 == 6'h1c; // @[Switch.scala 30:53:@9134.4]
  assign valid_28_36 = io_inValid_36 & _T_28542; // @[Switch.scala 30:36:@9135.4]
  assign _T_28545 = io_inAddr_37 == 6'h1c; // @[Switch.scala 30:53:@9137.4]
  assign valid_28_37 = io_inValid_37 & _T_28545; // @[Switch.scala 30:36:@9138.4]
  assign _T_28548 = io_inAddr_38 == 6'h1c; // @[Switch.scala 30:53:@9140.4]
  assign valid_28_38 = io_inValid_38 & _T_28548; // @[Switch.scala 30:36:@9141.4]
  assign _T_28551 = io_inAddr_39 == 6'h1c; // @[Switch.scala 30:53:@9143.4]
  assign valid_28_39 = io_inValid_39 & _T_28551; // @[Switch.scala 30:36:@9144.4]
  assign _T_28554 = io_inAddr_40 == 6'h1c; // @[Switch.scala 30:53:@9146.4]
  assign valid_28_40 = io_inValid_40 & _T_28554; // @[Switch.scala 30:36:@9147.4]
  assign _T_28557 = io_inAddr_41 == 6'h1c; // @[Switch.scala 30:53:@9149.4]
  assign valid_28_41 = io_inValid_41 & _T_28557; // @[Switch.scala 30:36:@9150.4]
  assign _T_28560 = io_inAddr_42 == 6'h1c; // @[Switch.scala 30:53:@9152.4]
  assign valid_28_42 = io_inValid_42 & _T_28560; // @[Switch.scala 30:36:@9153.4]
  assign _T_28563 = io_inAddr_43 == 6'h1c; // @[Switch.scala 30:53:@9155.4]
  assign valid_28_43 = io_inValid_43 & _T_28563; // @[Switch.scala 30:36:@9156.4]
  assign _T_28566 = io_inAddr_44 == 6'h1c; // @[Switch.scala 30:53:@9158.4]
  assign valid_28_44 = io_inValid_44 & _T_28566; // @[Switch.scala 30:36:@9159.4]
  assign _T_28569 = io_inAddr_45 == 6'h1c; // @[Switch.scala 30:53:@9161.4]
  assign valid_28_45 = io_inValid_45 & _T_28569; // @[Switch.scala 30:36:@9162.4]
  assign _T_28572 = io_inAddr_46 == 6'h1c; // @[Switch.scala 30:53:@9164.4]
  assign valid_28_46 = io_inValid_46 & _T_28572; // @[Switch.scala 30:36:@9165.4]
  assign _T_28575 = io_inAddr_47 == 6'h1c; // @[Switch.scala 30:53:@9167.4]
  assign valid_28_47 = io_inValid_47 & _T_28575; // @[Switch.scala 30:36:@9168.4]
  assign _T_28578 = io_inAddr_48 == 6'h1c; // @[Switch.scala 30:53:@9170.4]
  assign valid_28_48 = io_inValid_48 & _T_28578; // @[Switch.scala 30:36:@9171.4]
  assign _T_28581 = io_inAddr_49 == 6'h1c; // @[Switch.scala 30:53:@9173.4]
  assign valid_28_49 = io_inValid_49 & _T_28581; // @[Switch.scala 30:36:@9174.4]
  assign _T_28584 = io_inAddr_50 == 6'h1c; // @[Switch.scala 30:53:@9176.4]
  assign valid_28_50 = io_inValid_50 & _T_28584; // @[Switch.scala 30:36:@9177.4]
  assign _T_28587 = io_inAddr_51 == 6'h1c; // @[Switch.scala 30:53:@9179.4]
  assign valid_28_51 = io_inValid_51 & _T_28587; // @[Switch.scala 30:36:@9180.4]
  assign _T_28590 = io_inAddr_52 == 6'h1c; // @[Switch.scala 30:53:@9182.4]
  assign valid_28_52 = io_inValid_52 & _T_28590; // @[Switch.scala 30:36:@9183.4]
  assign _T_28593 = io_inAddr_53 == 6'h1c; // @[Switch.scala 30:53:@9185.4]
  assign valid_28_53 = io_inValid_53 & _T_28593; // @[Switch.scala 30:36:@9186.4]
  assign _T_28596 = io_inAddr_54 == 6'h1c; // @[Switch.scala 30:53:@9188.4]
  assign valid_28_54 = io_inValid_54 & _T_28596; // @[Switch.scala 30:36:@9189.4]
  assign _T_28599 = io_inAddr_55 == 6'h1c; // @[Switch.scala 30:53:@9191.4]
  assign valid_28_55 = io_inValid_55 & _T_28599; // @[Switch.scala 30:36:@9192.4]
  assign _T_28602 = io_inAddr_56 == 6'h1c; // @[Switch.scala 30:53:@9194.4]
  assign valid_28_56 = io_inValid_56 & _T_28602; // @[Switch.scala 30:36:@9195.4]
  assign _T_28605 = io_inAddr_57 == 6'h1c; // @[Switch.scala 30:53:@9197.4]
  assign valid_28_57 = io_inValid_57 & _T_28605; // @[Switch.scala 30:36:@9198.4]
  assign _T_28608 = io_inAddr_58 == 6'h1c; // @[Switch.scala 30:53:@9200.4]
  assign valid_28_58 = io_inValid_58 & _T_28608; // @[Switch.scala 30:36:@9201.4]
  assign _T_28611 = io_inAddr_59 == 6'h1c; // @[Switch.scala 30:53:@9203.4]
  assign valid_28_59 = io_inValid_59 & _T_28611; // @[Switch.scala 30:36:@9204.4]
  assign _T_28614 = io_inAddr_60 == 6'h1c; // @[Switch.scala 30:53:@9206.4]
  assign valid_28_60 = io_inValid_60 & _T_28614; // @[Switch.scala 30:36:@9207.4]
  assign _T_28617 = io_inAddr_61 == 6'h1c; // @[Switch.scala 30:53:@9209.4]
  assign valid_28_61 = io_inValid_61 & _T_28617; // @[Switch.scala 30:36:@9210.4]
  assign _T_28620 = io_inAddr_62 == 6'h1c; // @[Switch.scala 30:53:@9212.4]
  assign valid_28_62 = io_inValid_62 & _T_28620; // @[Switch.scala 30:36:@9213.4]
  assign _T_28623 = io_inAddr_63 == 6'h1c; // @[Switch.scala 30:53:@9215.4]
  assign valid_28_63 = io_inValid_63 & _T_28623; // @[Switch.scala 30:36:@9216.4]
  assign _T_28689 = valid_28_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@9218.4]
  assign _T_28690 = valid_28_61 ? 6'h3d : _T_28689; // @[Mux.scala 31:69:@9219.4]
  assign _T_28691 = valid_28_60 ? 6'h3c : _T_28690; // @[Mux.scala 31:69:@9220.4]
  assign _T_28692 = valid_28_59 ? 6'h3b : _T_28691; // @[Mux.scala 31:69:@9221.4]
  assign _T_28693 = valid_28_58 ? 6'h3a : _T_28692; // @[Mux.scala 31:69:@9222.4]
  assign _T_28694 = valid_28_57 ? 6'h39 : _T_28693; // @[Mux.scala 31:69:@9223.4]
  assign _T_28695 = valid_28_56 ? 6'h38 : _T_28694; // @[Mux.scala 31:69:@9224.4]
  assign _T_28696 = valid_28_55 ? 6'h37 : _T_28695; // @[Mux.scala 31:69:@9225.4]
  assign _T_28697 = valid_28_54 ? 6'h36 : _T_28696; // @[Mux.scala 31:69:@9226.4]
  assign _T_28698 = valid_28_53 ? 6'h35 : _T_28697; // @[Mux.scala 31:69:@9227.4]
  assign _T_28699 = valid_28_52 ? 6'h34 : _T_28698; // @[Mux.scala 31:69:@9228.4]
  assign _T_28700 = valid_28_51 ? 6'h33 : _T_28699; // @[Mux.scala 31:69:@9229.4]
  assign _T_28701 = valid_28_50 ? 6'h32 : _T_28700; // @[Mux.scala 31:69:@9230.4]
  assign _T_28702 = valid_28_49 ? 6'h31 : _T_28701; // @[Mux.scala 31:69:@9231.4]
  assign _T_28703 = valid_28_48 ? 6'h30 : _T_28702; // @[Mux.scala 31:69:@9232.4]
  assign _T_28704 = valid_28_47 ? 6'h2f : _T_28703; // @[Mux.scala 31:69:@9233.4]
  assign _T_28705 = valid_28_46 ? 6'h2e : _T_28704; // @[Mux.scala 31:69:@9234.4]
  assign _T_28706 = valid_28_45 ? 6'h2d : _T_28705; // @[Mux.scala 31:69:@9235.4]
  assign _T_28707 = valid_28_44 ? 6'h2c : _T_28706; // @[Mux.scala 31:69:@9236.4]
  assign _T_28708 = valid_28_43 ? 6'h2b : _T_28707; // @[Mux.scala 31:69:@9237.4]
  assign _T_28709 = valid_28_42 ? 6'h2a : _T_28708; // @[Mux.scala 31:69:@9238.4]
  assign _T_28710 = valid_28_41 ? 6'h29 : _T_28709; // @[Mux.scala 31:69:@9239.4]
  assign _T_28711 = valid_28_40 ? 6'h28 : _T_28710; // @[Mux.scala 31:69:@9240.4]
  assign _T_28712 = valid_28_39 ? 6'h27 : _T_28711; // @[Mux.scala 31:69:@9241.4]
  assign _T_28713 = valid_28_38 ? 6'h26 : _T_28712; // @[Mux.scala 31:69:@9242.4]
  assign _T_28714 = valid_28_37 ? 6'h25 : _T_28713; // @[Mux.scala 31:69:@9243.4]
  assign _T_28715 = valid_28_36 ? 6'h24 : _T_28714; // @[Mux.scala 31:69:@9244.4]
  assign _T_28716 = valid_28_35 ? 6'h23 : _T_28715; // @[Mux.scala 31:69:@9245.4]
  assign _T_28717 = valid_28_34 ? 6'h22 : _T_28716; // @[Mux.scala 31:69:@9246.4]
  assign _T_28718 = valid_28_33 ? 6'h21 : _T_28717; // @[Mux.scala 31:69:@9247.4]
  assign _T_28719 = valid_28_32 ? 6'h20 : _T_28718; // @[Mux.scala 31:69:@9248.4]
  assign _T_28720 = valid_28_31 ? 6'h1f : _T_28719; // @[Mux.scala 31:69:@9249.4]
  assign _T_28721 = valid_28_30 ? 6'h1e : _T_28720; // @[Mux.scala 31:69:@9250.4]
  assign _T_28722 = valid_28_29 ? 6'h1d : _T_28721; // @[Mux.scala 31:69:@9251.4]
  assign _T_28723 = valid_28_28 ? 6'h1c : _T_28722; // @[Mux.scala 31:69:@9252.4]
  assign _T_28724 = valid_28_27 ? 6'h1b : _T_28723; // @[Mux.scala 31:69:@9253.4]
  assign _T_28725 = valid_28_26 ? 6'h1a : _T_28724; // @[Mux.scala 31:69:@9254.4]
  assign _T_28726 = valid_28_25 ? 6'h19 : _T_28725; // @[Mux.scala 31:69:@9255.4]
  assign _T_28727 = valid_28_24 ? 6'h18 : _T_28726; // @[Mux.scala 31:69:@9256.4]
  assign _T_28728 = valid_28_23 ? 6'h17 : _T_28727; // @[Mux.scala 31:69:@9257.4]
  assign _T_28729 = valid_28_22 ? 6'h16 : _T_28728; // @[Mux.scala 31:69:@9258.4]
  assign _T_28730 = valid_28_21 ? 6'h15 : _T_28729; // @[Mux.scala 31:69:@9259.4]
  assign _T_28731 = valid_28_20 ? 6'h14 : _T_28730; // @[Mux.scala 31:69:@9260.4]
  assign _T_28732 = valid_28_19 ? 6'h13 : _T_28731; // @[Mux.scala 31:69:@9261.4]
  assign _T_28733 = valid_28_18 ? 6'h12 : _T_28732; // @[Mux.scala 31:69:@9262.4]
  assign _T_28734 = valid_28_17 ? 6'h11 : _T_28733; // @[Mux.scala 31:69:@9263.4]
  assign _T_28735 = valid_28_16 ? 6'h10 : _T_28734; // @[Mux.scala 31:69:@9264.4]
  assign _T_28736 = valid_28_15 ? 6'hf : _T_28735; // @[Mux.scala 31:69:@9265.4]
  assign _T_28737 = valid_28_14 ? 6'he : _T_28736; // @[Mux.scala 31:69:@9266.4]
  assign _T_28738 = valid_28_13 ? 6'hd : _T_28737; // @[Mux.scala 31:69:@9267.4]
  assign _T_28739 = valid_28_12 ? 6'hc : _T_28738; // @[Mux.scala 31:69:@9268.4]
  assign _T_28740 = valid_28_11 ? 6'hb : _T_28739; // @[Mux.scala 31:69:@9269.4]
  assign _T_28741 = valid_28_10 ? 6'ha : _T_28740; // @[Mux.scala 31:69:@9270.4]
  assign _T_28742 = valid_28_9 ? 6'h9 : _T_28741; // @[Mux.scala 31:69:@9271.4]
  assign _T_28743 = valid_28_8 ? 6'h8 : _T_28742; // @[Mux.scala 31:69:@9272.4]
  assign _T_28744 = valid_28_7 ? 6'h7 : _T_28743; // @[Mux.scala 31:69:@9273.4]
  assign _T_28745 = valid_28_6 ? 6'h6 : _T_28744; // @[Mux.scala 31:69:@9274.4]
  assign _T_28746 = valid_28_5 ? 6'h5 : _T_28745; // @[Mux.scala 31:69:@9275.4]
  assign _T_28747 = valid_28_4 ? 6'h4 : _T_28746; // @[Mux.scala 31:69:@9276.4]
  assign _T_28748 = valid_28_3 ? 6'h3 : _T_28747; // @[Mux.scala 31:69:@9277.4]
  assign _T_28749 = valid_28_2 ? 6'h2 : _T_28748; // @[Mux.scala 31:69:@9278.4]
  assign _T_28750 = valid_28_1 ? 6'h1 : _T_28749; // @[Mux.scala 31:69:@9279.4]
  assign select_28 = valid_28_0 ? 6'h0 : _T_28750; // @[Mux.scala 31:69:@9280.4]
  assign _GEN_1793 = 6'h1 == select_28 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1794 = 6'h2 == select_28 ? io_inData_2 : _GEN_1793; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1795 = 6'h3 == select_28 ? io_inData_3 : _GEN_1794; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1796 = 6'h4 == select_28 ? io_inData_4 : _GEN_1795; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1797 = 6'h5 == select_28 ? io_inData_5 : _GEN_1796; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1798 = 6'h6 == select_28 ? io_inData_6 : _GEN_1797; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1799 = 6'h7 == select_28 ? io_inData_7 : _GEN_1798; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1800 = 6'h8 == select_28 ? io_inData_8 : _GEN_1799; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1801 = 6'h9 == select_28 ? io_inData_9 : _GEN_1800; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1802 = 6'ha == select_28 ? io_inData_10 : _GEN_1801; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1803 = 6'hb == select_28 ? io_inData_11 : _GEN_1802; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1804 = 6'hc == select_28 ? io_inData_12 : _GEN_1803; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1805 = 6'hd == select_28 ? io_inData_13 : _GEN_1804; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1806 = 6'he == select_28 ? io_inData_14 : _GEN_1805; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1807 = 6'hf == select_28 ? io_inData_15 : _GEN_1806; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1808 = 6'h10 == select_28 ? io_inData_16 : _GEN_1807; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1809 = 6'h11 == select_28 ? io_inData_17 : _GEN_1808; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1810 = 6'h12 == select_28 ? io_inData_18 : _GEN_1809; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1811 = 6'h13 == select_28 ? io_inData_19 : _GEN_1810; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1812 = 6'h14 == select_28 ? io_inData_20 : _GEN_1811; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1813 = 6'h15 == select_28 ? io_inData_21 : _GEN_1812; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1814 = 6'h16 == select_28 ? io_inData_22 : _GEN_1813; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1815 = 6'h17 == select_28 ? io_inData_23 : _GEN_1814; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1816 = 6'h18 == select_28 ? io_inData_24 : _GEN_1815; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1817 = 6'h19 == select_28 ? io_inData_25 : _GEN_1816; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1818 = 6'h1a == select_28 ? io_inData_26 : _GEN_1817; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1819 = 6'h1b == select_28 ? io_inData_27 : _GEN_1818; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1820 = 6'h1c == select_28 ? io_inData_28 : _GEN_1819; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1821 = 6'h1d == select_28 ? io_inData_29 : _GEN_1820; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1822 = 6'h1e == select_28 ? io_inData_30 : _GEN_1821; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1823 = 6'h1f == select_28 ? io_inData_31 : _GEN_1822; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1824 = 6'h20 == select_28 ? io_inData_32 : _GEN_1823; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1825 = 6'h21 == select_28 ? io_inData_33 : _GEN_1824; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1826 = 6'h22 == select_28 ? io_inData_34 : _GEN_1825; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1827 = 6'h23 == select_28 ? io_inData_35 : _GEN_1826; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1828 = 6'h24 == select_28 ? io_inData_36 : _GEN_1827; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1829 = 6'h25 == select_28 ? io_inData_37 : _GEN_1828; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1830 = 6'h26 == select_28 ? io_inData_38 : _GEN_1829; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1831 = 6'h27 == select_28 ? io_inData_39 : _GEN_1830; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1832 = 6'h28 == select_28 ? io_inData_40 : _GEN_1831; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1833 = 6'h29 == select_28 ? io_inData_41 : _GEN_1832; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1834 = 6'h2a == select_28 ? io_inData_42 : _GEN_1833; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1835 = 6'h2b == select_28 ? io_inData_43 : _GEN_1834; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1836 = 6'h2c == select_28 ? io_inData_44 : _GEN_1835; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1837 = 6'h2d == select_28 ? io_inData_45 : _GEN_1836; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1838 = 6'h2e == select_28 ? io_inData_46 : _GEN_1837; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1839 = 6'h2f == select_28 ? io_inData_47 : _GEN_1838; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1840 = 6'h30 == select_28 ? io_inData_48 : _GEN_1839; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1841 = 6'h31 == select_28 ? io_inData_49 : _GEN_1840; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1842 = 6'h32 == select_28 ? io_inData_50 : _GEN_1841; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1843 = 6'h33 == select_28 ? io_inData_51 : _GEN_1842; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1844 = 6'h34 == select_28 ? io_inData_52 : _GEN_1843; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1845 = 6'h35 == select_28 ? io_inData_53 : _GEN_1844; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1846 = 6'h36 == select_28 ? io_inData_54 : _GEN_1845; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1847 = 6'h37 == select_28 ? io_inData_55 : _GEN_1846; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1848 = 6'h38 == select_28 ? io_inData_56 : _GEN_1847; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1849 = 6'h39 == select_28 ? io_inData_57 : _GEN_1848; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1850 = 6'h3a == select_28 ? io_inData_58 : _GEN_1849; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1851 = 6'h3b == select_28 ? io_inData_59 : _GEN_1850; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1852 = 6'h3c == select_28 ? io_inData_60 : _GEN_1851; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1853 = 6'h3d == select_28 ? io_inData_61 : _GEN_1852; // @[Switch.scala 33:19:@9282.4]
  assign _GEN_1854 = 6'h3e == select_28 ? io_inData_62 : _GEN_1853; // @[Switch.scala 33:19:@9282.4]
  assign _T_28759 = {valid_28_7,valid_28_6,valid_28_5,valid_28_4,valid_28_3,valid_28_2,valid_28_1,valid_28_0}; // @[Switch.scala 34:32:@9289.4]
  assign _T_28767 = {valid_28_15,valid_28_14,valid_28_13,valid_28_12,valid_28_11,valid_28_10,valid_28_9,valid_28_8,_T_28759}; // @[Switch.scala 34:32:@9297.4]
  assign _T_28774 = {valid_28_23,valid_28_22,valid_28_21,valid_28_20,valid_28_19,valid_28_18,valid_28_17,valid_28_16}; // @[Switch.scala 34:32:@9304.4]
  assign _T_28783 = {valid_28_31,valid_28_30,valid_28_29,valid_28_28,valid_28_27,valid_28_26,valid_28_25,valid_28_24,_T_28774,_T_28767}; // @[Switch.scala 34:32:@9313.4]
  assign _T_28790 = {valid_28_39,valid_28_38,valid_28_37,valid_28_36,valid_28_35,valid_28_34,valid_28_33,valid_28_32}; // @[Switch.scala 34:32:@9320.4]
  assign _T_28798 = {valid_28_47,valid_28_46,valid_28_45,valid_28_44,valid_28_43,valid_28_42,valid_28_41,valid_28_40,_T_28790}; // @[Switch.scala 34:32:@9328.4]
  assign _T_28805 = {valid_28_55,valid_28_54,valid_28_53,valid_28_52,valid_28_51,valid_28_50,valid_28_49,valid_28_48}; // @[Switch.scala 34:32:@9335.4]
  assign _T_28814 = {valid_28_63,valid_28_62,valid_28_61,valid_28_60,valid_28_59,valid_28_58,valid_28_57,valid_28_56,_T_28805,_T_28798}; // @[Switch.scala 34:32:@9344.4]
  assign _T_28815 = {_T_28814,_T_28783}; // @[Switch.scala 34:32:@9345.4]
  assign _T_28819 = io_inAddr_0 == 6'h1d; // @[Switch.scala 30:53:@9348.4]
  assign valid_29_0 = io_inValid_0 & _T_28819; // @[Switch.scala 30:36:@9349.4]
  assign _T_28822 = io_inAddr_1 == 6'h1d; // @[Switch.scala 30:53:@9351.4]
  assign valid_29_1 = io_inValid_1 & _T_28822; // @[Switch.scala 30:36:@9352.4]
  assign _T_28825 = io_inAddr_2 == 6'h1d; // @[Switch.scala 30:53:@9354.4]
  assign valid_29_2 = io_inValid_2 & _T_28825; // @[Switch.scala 30:36:@9355.4]
  assign _T_28828 = io_inAddr_3 == 6'h1d; // @[Switch.scala 30:53:@9357.4]
  assign valid_29_3 = io_inValid_3 & _T_28828; // @[Switch.scala 30:36:@9358.4]
  assign _T_28831 = io_inAddr_4 == 6'h1d; // @[Switch.scala 30:53:@9360.4]
  assign valid_29_4 = io_inValid_4 & _T_28831; // @[Switch.scala 30:36:@9361.4]
  assign _T_28834 = io_inAddr_5 == 6'h1d; // @[Switch.scala 30:53:@9363.4]
  assign valid_29_5 = io_inValid_5 & _T_28834; // @[Switch.scala 30:36:@9364.4]
  assign _T_28837 = io_inAddr_6 == 6'h1d; // @[Switch.scala 30:53:@9366.4]
  assign valid_29_6 = io_inValid_6 & _T_28837; // @[Switch.scala 30:36:@9367.4]
  assign _T_28840 = io_inAddr_7 == 6'h1d; // @[Switch.scala 30:53:@9369.4]
  assign valid_29_7 = io_inValid_7 & _T_28840; // @[Switch.scala 30:36:@9370.4]
  assign _T_28843 = io_inAddr_8 == 6'h1d; // @[Switch.scala 30:53:@9372.4]
  assign valid_29_8 = io_inValid_8 & _T_28843; // @[Switch.scala 30:36:@9373.4]
  assign _T_28846 = io_inAddr_9 == 6'h1d; // @[Switch.scala 30:53:@9375.4]
  assign valid_29_9 = io_inValid_9 & _T_28846; // @[Switch.scala 30:36:@9376.4]
  assign _T_28849 = io_inAddr_10 == 6'h1d; // @[Switch.scala 30:53:@9378.4]
  assign valid_29_10 = io_inValid_10 & _T_28849; // @[Switch.scala 30:36:@9379.4]
  assign _T_28852 = io_inAddr_11 == 6'h1d; // @[Switch.scala 30:53:@9381.4]
  assign valid_29_11 = io_inValid_11 & _T_28852; // @[Switch.scala 30:36:@9382.4]
  assign _T_28855 = io_inAddr_12 == 6'h1d; // @[Switch.scala 30:53:@9384.4]
  assign valid_29_12 = io_inValid_12 & _T_28855; // @[Switch.scala 30:36:@9385.4]
  assign _T_28858 = io_inAddr_13 == 6'h1d; // @[Switch.scala 30:53:@9387.4]
  assign valid_29_13 = io_inValid_13 & _T_28858; // @[Switch.scala 30:36:@9388.4]
  assign _T_28861 = io_inAddr_14 == 6'h1d; // @[Switch.scala 30:53:@9390.4]
  assign valid_29_14 = io_inValid_14 & _T_28861; // @[Switch.scala 30:36:@9391.4]
  assign _T_28864 = io_inAddr_15 == 6'h1d; // @[Switch.scala 30:53:@9393.4]
  assign valid_29_15 = io_inValid_15 & _T_28864; // @[Switch.scala 30:36:@9394.4]
  assign _T_28867 = io_inAddr_16 == 6'h1d; // @[Switch.scala 30:53:@9396.4]
  assign valid_29_16 = io_inValid_16 & _T_28867; // @[Switch.scala 30:36:@9397.4]
  assign _T_28870 = io_inAddr_17 == 6'h1d; // @[Switch.scala 30:53:@9399.4]
  assign valid_29_17 = io_inValid_17 & _T_28870; // @[Switch.scala 30:36:@9400.4]
  assign _T_28873 = io_inAddr_18 == 6'h1d; // @[Switch.scala 30:53:@9402.4]
  assign valid_29_18 = io_inValid_18 & _T_28873; // @[Switch.scala 30:36:@9403.4]
  assign _T_28876 = io_inAddr_19 == 6'h1d; // @[Switch.scala 30:53:@9405.4]
  assign valid_29_19 = io_inValid_19 & _T_28876; // @[Switch.scala 30:36:@9406.4]
  assign _T_28879 = io_inAddr_20 == 6'h1d; // @[Switch.scala 30:53:@9408.4]
  assign valid_29_20 = io_inValid_20 & _T_28879; // @[Switch.scala 30:36:@9409.4]
  assign _T_28882 = io_inAddr_21 == 6'h1d; // @[Switch.scala 30:53:@9411.4]
  assign valid_29_21 = io_inValid_21 & _T_28882; // @[Switch.scala 30:36:@9412.4]
  assign _T_28885 = io_inAddr_22 == 6'h1d; // @[Switch.scala 30:53:@9414.4]
  assign valid_29_22 = io_inValid_22 & _T_28885; // @[Switch.scala 30:36:@9415.4]
  assign _T_28888 = io_inAddr_23 == 6'h1d; // @[Switch.scala 30:53:@9417.4]
  assign valid_29_23 = io_inValid_23 & _T_28888; // @[Switch.scala 30:36:@9418.4]
  assign _T_28891 = io_inAddr_24 == 6'h1d; // @[Switch.scala 30:53:@9420.4]
  assign valid_29_24 = io_inValid_24 & _T_28891; // @[Switch.scala 30:36:@9421.4]
  assign _T_28894 = io_inAddr_25 == 6'h1d; // @[Switch.scala 30:53:@9423.4]
  assign valid_29_25 = io_inValid_25 & _T_28894; // @[Switch.scala 30:36:@9424.4]
  assign _T_28897 = io_inAddr_26 == 6'h1d; // @[Switch.scala 30:53:@9426.4]
  assign valid_29_26 = io_inValid_26 & _T_28897; // @[Switch.scala 30:36:@9427.4]
  assign _T_28900 = io_inAddr_27 == 6'h1d; // @[Switch.scala 30:53:@9429.4]
  assign valid_29_27 = io_inValid_27 & _T_28900; // @[Switch.scala 30:36:@9430.4]
  assign _T_28903 = io_inAddr_28 == 6'h1d; // @[Switch.scala 30:53:@9432.4]
  assign valid_29_28 = io_inValid_28 & _T_28903; // @[Switch.scala 30:36:@9433.4]
  assign _T_28906 = io_inAddr_29 == 6'h1d; // @[Switch.scala 30:53:@9435.4]
  assign valid_29_29 = io_inValid_29 & _T_28906; // @[Switch.scala 30:36:@9436.4]
  assign _T_28909 = io_inAddr_30 == 6'h1d; // @[Switch.scala 30:53:@9438.4]
  assign valid_29_30 = io_inValid_30 & _T_28909; // @[Switch.scala 30:36:@9439.4]
  assign _T_28912 = io_inAddr_31 == 6'h1d; // @[Switch.scala 30:53:@9441.4]
  assign valid_29_31 = io_inValid_31 & _T_28912; // @[Switch.scala 30:36:@9442.4]
  assign _T_28915 = io_inAddr_32 == 6'h1d; // @[Switch.scala 30:53:@9444.4]
  assign valid_29_32 = io_inValid_32 & _T_28915; // @[Switch.scala 30:36:@9445.4]
  assign _T_28918 = io_inAddr_33 == 6'h1d; // @[Switch.scala 30:53:@9447.4]
  assign valid_29_33 = io_inValid_33 & _T_28918; // @[Switch.scala 30:36:@9448.4]
  assign _T_28921 = io_inAddr_34 == 6'h1d; // @[Switch.scala 30:53:@9450.4]
  assign valid_29_34 = io_inValid_34 & _T_28921; // @[Switch.scala 30:36:@9451.4]
  assign _T_28924 = io_inAddr_35 == 6'h1d; // @[Switch.scala 30:53:@9453.4]
  assign valid_29_35 = io_inValid_35 & _T_28924; // @[Switch.scala 30:36:@9454.4]
  assign _T_28927 = io_inAddr_36 == 6'h1d; // @[Switch.scala 30:53:@9456.4]
  assign valid_29_36 = io_inValid_36 & _T_28927; // @[Switch.scala 30:36:@9457.4]
  assign _T_28930 = io_inAddr_37 == 6'h1d; // @[Switch.scala 30:53:@9459.4]
  assign valid_29_37 = io_inValid_37 & _T_28930; // @[Switch.scala 30:36:@9460.4]
  assign _T_28933 = io_inAddr_38 == 6'h1d; // @[Switch.scala 30:53:@9462.4]
  assign valid_29_38 = io_inValid_38 & _T_28933; // @[Switch.scala 30:36:@9463.4]
  assign _T_28936 = io_inAddr_39 == 6'h1d; // @[Switch.scala 30:53:@9465.4]
  assign valid_29_39 = io_inValid_39 & _T_28936; // @[Switch.scala 30:36:@9466.4]
  assign _T_28939 = io_inAddr_40 == 6'h1d; // @[Switch.scala 30:53:@9468.4]
  assign valid_29_40 = io_inValid_40 & _T_28939; // @[Switch.scala 30:36:@9469.4]
  assign _T_28942 = io_inAddr_41 == 6'h1d; // @[Switch.scala 30:53:@9471.4]
  assign valid_29_41 = io_inValid_41 & _T_28942; // @[Switch.scala 30:36:@9472.4]
  assign _T_28945 = io_inAddr_42 == 6'h1d; // @[Switch.scala 30:53:@9474.4]
  assign valid_29_42 = io_inValid_42 & _T_28945; // @[Switch.scala 30:36:@9475.4]
  assign _T_28948 = io_inAddr_43 == 6'h1d; // @[Switch.scala 30:53:@9477.4]
  assign valid_29_43 = io_inValid_43 & _T_28948; // @[Switch.scala 30:36:@9478.4]
  assign _T_28951 = io_inAddr_44 == 6'h1d; // @[Switch.scala 30:53:@9480.4]
  assign valid_29_44 = io_inValid_44 & _T_28951; // @[Switch.scala 30:36:@9481.4]
  assign _T_28954 = io_inAddr_45 == 6'h1d; // @[Switch.scala 30:53:@9483.4]
  assign valid_29_45 = io_inValid_45 & _T_28954; // @[Switch.scala 30:36:@9484.4]
  assign _T_28957 = io_inAddr_46 == 6'h1d; // @[Switch.scala 30:53:@9486.4]
  assign valid_29_46 = io_inValid_46 & _T_28957; // @[Switch.scala 30:36:@9487.4]
  assign _T_28960 = io_inAddr_47 == 6'h1d; // @[Switch.scala 30:53:@9489.4]
  assign valid_29_47 = io_inValid_47 & _T_28960; // @[Switch.scala 30:36:@9490.4]
  assign _T_28963 = io_inAddr_48 == 6'h1d; // @[Switch.scala 30:53:@9492.4]
  assign valid_29_48 = io_inValid_48 & _T_28963; // @[Switch.scala 30:36:@9493.4]
  assign _T_28966 = io_inAddr_49 == 6'h1d; // @[Switch.scala 30:53:@9495.4]
  assign valid_29_49 = io_inValid_49 & _T_28966; // @[Switch.scala 30:36:@9496.4]
  assign _T_28969 = io_inAddr_50 == 6'h1d; // @[Switch.scala 30:53:@9498.4]
  assign valid_29_50 = io_inValid_50 & _T_28969; // @[Switch.scala 30:36:@9499.4]
  assign _T_28972 = io_inAddr_51 == 6'h1d; // @[Switch.scala 30:53:@9501.4]
  assign valid_29_51 = io_inValid_51 & _T_28972; // @[Switch.scala 30:36:@9502.4]
  assign _T_28975 = io_inAddr_52 == 6'h1d; // @[Switch.scala 30:53:@9504.4]
  assign valid_29_52 = io_inValid_52 & _T_28975; // @[Switch.scala 30:36:@9505.4]
  assign _T_28978 = io_inAddr_53 == 6'h1d; // @[Switch.scala 30:53:@9507.4]
  assign valid_29_53 = io_inValid_53 & _T_28978; // @[Switch.scala 30:36:@9508.4]
  assign _T_28981 = io_inAddr_54 == 6'h1d; // @[Switch.scala 30:53:@9510.4]
  assign valid_29_54 = io_inValid_54 & _T_28981; // @[Switch.scala 30:36:@9511.4]
  assign _T_28984 = io_inAddr_55 == 6'h1d; // @[Switch.scala 30:53:@9513.4]
  assign valid_29_55 = io_inValid_55 & _T_28984; // @[Switch.scala 30:36:@9514.4]
  assign _T_28987 = io_inAddr_56 == 6'h1d; // @[Switch.scala 30:53:@9516.4]
  assign valid_29_56 = io_inValid_56 & _T_28987; // @[Switch.scala 30:36:@9517.4]
  assign _T_28990 = io_inAddr_57 == 6'h1d; // @[Switch.scala 30:53:@9519.4]
  assign valid_29_57 = io_inValid_57 & _T_28990; // @[Switch.scala 30:36:@9520.4]
  assign _T_28993 = io_inAddr_58 == 6'h1d; // @[Switch.scala 30:53:@9522.4]
  assign valid_29_58 = io_inValid_58 & _T_28993; // @[Switch.scala 30:36:@9523.4]
  assign _T_28996 = io_inAddr_59 == 6'h1d; // @[Switch.scala 30:53:@9525.4]
  assign valid_29_59 = io_inValid_59 & _T_28996; // @[Switch.scala 30:36:@9526.4]
  assign _T_28999 = io_inAddr_60 == 6'h1d; // @[Switch.scala 30:53:@9528.4]
  assign valid_29_60 = io_inValid_60 & _T_28999; // @[Switch.scala 30:36:@9529.4]
  assign _T_29002 = io_inAddr_61 == 6'h1d; // @[Switch.scala 30:53:@9531.4]
  assign valid_29_61 = io_inValid_61 & _T_29002; // @[Switch.scala 30:36:@9532.4]
  assign _T_29005 = io_inAddr_62 == 6'h1d; // @[Switch.scala 30:53:@9534.4]
  assign valid_29_62 = io_inValid_62 & _T_29005; // @[Switch.scala 30:36:@9535.4]
  assign _T_29008 = io_inAddr_63 == 6'h1d; // @[Switch.scala 30:53:@9537.4]
  assign valid_29_63 = io_inValid_63 & _T_29008; // @[Switch.scala 30:36:@9538.4]
  assign _T_29074 = valid_29_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@9540.4]
  assign _T_29075 = valid_29_61 ? 6'h3d : _T_29074; // @[Mux.scala 31:69:@9541.4]
  assign _T_29076 = valid_29_60 ? 6'h3c : _T_29075; // @[Mux.scala 31:69:@9542.4]
  assign _T_29077 = valid_29_59 ? 6'h3b : _T_29076; // @[Mux.scala 31:69:@9543.4]
  assign _T_29078 = valid_29_58 ? 6'h3a : _T_29077; // @[Mux.scala 31:69:@9544.4]
  assign _T_29079 = valid_29_57 ? 6'h39 : _T_29078; // @[Mux.scala 31:69:@9545.4]
  assign _T_29080 = valid_29_56 ? 6'h38 : _T_29079; // @[Mux.scala 31:69:@9546.4]
  assign _T_29081 = valid_29_55 ? 6'h37 : _T_29080; // @[Mux.scala 31:69:@9547.4]
  assign _T_29082 = valid_29_54 ? 6'h36 : _T_29081; // @[Mux.scala 31:69:@9548.4]
  assign _T_29083 = valid_29_53 ? 6'h35 : _T_29082; // @[Mux.scala 31:69:@9549.4]
  assign _T_29084 = valid_29_52 ? 6'h34 : _T_29083; // @[Mux.scala 31:69:@9550.4]
  assign _T_29085 = valid_29_51 ? 6'h33 : _T_29084; // @[Mux.scala 31:69:@9551.4]
  assign _T_29086 = valid_29_50 ? 6'h32 : _T_29085; // @[Mux.scala 31:69:@9552.4]
  assign _T_29087 = valid_29_49 ? 6'h31 : _T_29086; // @[Mux.scala 31:69:@9553.4]
  assign _T_29088 = valid_29_48 ? 6'h30 : _T_29087; // @[Mux.scala 31:69:@9554.4]
  assign _T_29089 = valid_29_47 ? 6'h2f : _T_29088; // @[Mux.scala 31:69:@9555.4]
  assign _T_29090 = valid_29_46 ? 6'h2e : _T_29089; // @[Mux.scala 31:69:@9556.4]
  assign _T_29091 = valid_29_45 ? 6'h2d : _T_29090; // @[Mux.scala 31:69:@9557.4]
  assign _T_29092 = valid_29_44 ? 6'h2c : _T_29091; // @[Mux.scala 31:69:@9558.4]
  assign _T_29093 = valid_29_43 ? 6'h2b : _T_29092; // @[Mux.scala 31:69:@9559.4]
  assign _T_29094 = valid_29_42 ? 6'h2a : _T_29093; // @[Mux.scala 31:69:@9560.4]
  assign _T_29095 = valid_29_41 ? 6'h29 : _T_29094; // @[Mux.scala 31:69:@9561.4]
  assign _T_29096 = valid_29_40 ? 6'h28 : _T_29095; // @[Mux.scala 31:69:@9562.4]
  assign _T_29097 = valid_29_39 ? 6'h27 : _T_29096; // @[Mux.scala 31:69:@9563.4]
  assign _T_29098 = valid_29_38 ? 6'h26 : _T_29097; // @[Mux.scala 31:69:@9564.4]
  assign _T_29099 = valid_29_37 ? 6'h25 : _T_29098; // @[Mux.scala 31:69:@9565.4]
  assign _T_29100 = valid_29_36 ? 6'h24 : _T_29099; // @[Mux.scala 31:69:@9566.4]
  assign _T_29101 = valid_29_35 ? 6'h23 : _T_29100; // @[Mux.scala 31:69:@9567.4]
  assign _T_29102 = valid_29_34 ? 6'h22 : _T_29101; // @[Mux.scala 31:69:@9568.4]
  assign _T_29103 = valid_29_33 ? 6'h21 : _T_29102; // @[Mux.scala 31:69:@9569.4]
  assign _T_29104 = valid_29_32 ? 6'h20 : _T_29103; // @[Mux.scala 31:69:@9570.4]
  assign _T_29105 = valid_29_31 ? 6'h1f : _T_29104; // @[Mux.scala 31:69:@9571.4]
  assign _T_29106 = valid_29_30 ? 6'h1e : _T_29105; // @[Mux.scala 31:69:@9572.4]
  assign _T_29107 = valid_29_29 ? 6'h1d : _T_29106; // @[Mux.scala 31:69:@9573.4]
  assign _T_29108 = valid_29_28 ? 6'h1c : _T_29107; // @[Mux.scala 31:69:@9574.4]
  assign _T_29109 = valid_29_27 ? 6'h1b : _T_29108; // @[Mux.scala 31:69:@9575.4]
  assign _T_29110 = valid_29_26 ? 6'h1a : _T_29109; // @[Mux.scala 31:69:@9576.4]
  assign _T_29111 = valid_29_25 ? 6'h19 : _T_29110; // @[Mux.scala 31:69:@9577.4]
  assign _T_29112 = valid_29_24 ? 6'h18 : _T_29111; // @[Mux.scala 31:69:@9578.4]
  assign _T_29113 = valid_29_23 ? 6'h17 : _T_29112; // @[Mux.scala 31:69:@9579.4]
  assign _T_29114 = valid_29_22 ? 6'h16 : _T_29113; // @[Mux.scala 31:69:@9580.4]
  assign _T_29115 = valid_29_21 ? 6'h15 : _T_29114; // @[Mux.scala 31:69:@9581.4]
  assign _T_29116 = valid_29_20 ? 6'h14 : _T_29115; // @[Mux.scala 31:69:@9582.4]
  assign _T_29117 = valid_29_19 ? 6'h13 : _T_29116; // @[Mux.scala 31:69:@9583.4]
  assign _T_29118 = valid_29_18 ? 6'h12 : _T_29117; // @[Mux.scala 31:69:@9584.4]
  assign _T_29119 = valid_29_17 ? 6'h11 : _T_29118; // @[Mux.scala 31:69:@9585.4]
  assign _T_29120 = valid_29_16 ? 6'h10 : _T_29119; // @[Mux.scala 31:69:@9586.4]
  assign _T_29121 = valid_29_15 ? 6'hf : _T_29120; // @[Mux.scala 31:69:@9587.4]
  assign _T_29122 = valid_29_14 ? 6'he : _T_29121; // @[Mux.scala 31:69:@9588.4]
  assign _T_29123 = valid_29_13 ? 6'hd : _T_29122; // @[Mux.scala 31:69:@9589.4]
  assign _T_29124 = valid_29_12 ? 6'hc : _T_29123; // @[Mux.scala 31:69:@9590.4]
  assign _T_29125 = valid_29_11 ? 6'hb : _T_29124; // @[Mux.scala 31:69:@9591.4]
  assign _T_29126 = valid_29_10 ? 6'ha : _T_29125; // @[Mux.scala 31:69:@9592.4]
  assign _T_29127 = valid_29_9 ? 6'h9 : _T_29126; // @[Mux.scala 31:69:@9593.4]
  assign _T_29128 = valid_29_8 ? 6'h8 : _T_29127; // @[Mux.scala 31:69:@9594.4]
  assign _T_29129 = valid_29_7 ? 6'h7 : _T_29128; // @[Mux.scala 31:69:@9595.4]
  assign _T_29130 = valid_29_6 ? 6'h6 : _T_29129; // @[Mux.scala 31:69:@9596.4]
  assign _T_29131 = valid_29_5 ? 6'h5 : _T_29130; // @[Mux.scala 31:69:@9597.4]
  assign _T_29132 = valid_29_4 ? 6'h4 : _T_29131; // @[Mux.scala 31:69:@9598.4]
  assign _T_29133 = valid_29_3 ? 6'h3 : _T_29132; // @[Mux.scala 31:69:@9599.4]
  assign _T_29134 = valid_29_2 ? 6'h2 : _T_29133; // @[Mux.scala 31:69:@9600.4]
  assign _T_29135 = valid_29_1 ? 6'h1 : _T_29134; // @[Mux.scala 31:69:@9601.4]
  assign select_29 = valid_29_0 ? 6'h0 : _T_29135; // @[Mux.scala 31:69:@9602.4]
  assign _GEN_1857 = 6'h1 == select_29 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1858 = 6'h2 == select_29 ? io_inData_2 : _GEN_1857; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1859 = 6'h3 == select_29 ? io_inData_3 : _GEN_1858; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1860 = 6'h4 == select_29 ? io_inData_4 : _GEN_1859; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1861 = 6'h5 == select_29 ? io_inData_5 : _GEN_1860; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1862 = 6'h6 == select_29 ? io_inData_6 : _GEN_1861; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1863 = 6'h7 == select_29 ? io_inData_7 : _GEN_1862; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1864 = 6'h8 == select_29 ? io_inData_8 : _GEN_1863; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1865 = 6'h9 == select_29 ? io_inData_9 : _GEN_1864; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1866 = 6'ha == select_29 ? io_inData_10 : _GEN_1865; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1867 = 6'hb == select_29 ? io_inData_11 : _GEN_1866; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1868 = 6'hc == select_29 ? io_inData_12 : _GEN_1867; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1869 = 6'hd == select_29 ? io_inData_13 : _GEN_1868; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1870 = 6'he == select_29 ? io_inData_14 : _GEN_1869; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1871 = 6'hf == select_29 ? io_inData_15 : _GEN_1870; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1872 = 6'h10 == select_29 ? io_inData_16 : _GEN_1871; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1873 = 6'h11 == select_29 ? io_inData_17 : _GEN_1872; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1874 = 6'h12 == select_29 ? io_inData_18 : _GEN_1873; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1875 = 6'h13 == select_29 ? io_inData_19 : _GEN_1874; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1876 = 6'h14 == select_29 ? io_inData_20 : _GEN_1875; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1877 = 6'h15 == select_29 ? io_inData_21 : _GEN_1876; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1878 = 6'h16 == select_29 ? io_inData_22 : _GEN_1877; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1879 = 6'h17 == select_29 ? io_inData_23 : _GEN_1878; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1880 = 6'h18 == select_29 ? io_inData_24 : _GEN_1879; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1881 = 6'h19 == select_29 ? io_inData_25 : _GEN_1880; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1882 = 6'h1a == select_29 ? io_inData_26 : _GEN_1881; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1883 = 6'h1b == select_29 ? io_inData_27 : _GEN_1882; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1884 = 6'h1c == select_29 ? io_inData_28 : _GEN_1883; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1885 = 6'h1d == select_29 ? io_inData_29 : _GEN_1884; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1886 = 6'h1e == select_29 ? io_inData_30 : _GEN_1885; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1887 = 6'h1f == select_29 ? io_inData_31 : _GEN_1886; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1888 = 6'h20 == select_29 ? io_inData_32 : _GEN_1887; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1889 = 6'h21 == select_29 ? io_inData_33 : _GEN_1888; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1890 = 6'h22 == select_29 ? io_inData_34 : _GEN_1889; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1891 = 6'h23 == select_29 ? io_inData_35 : _GEN_1890; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1892 = 6'h24 == select_29 ? io_inData_36 : _GEN_1891; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1893 = 6'h25 == select_29 ? io_inData_37 : _GEN_1892; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1894 = 6'h26 == select_29 ? io_inData_38 : _GEN_1893; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1895 = 6'h27 == select_29 ? io_inData_39 : _GEN_1894; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1896 = 6'h28 == select_29 ? io_inData_40 : _GEN_1895; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1897 = 6'h29 == select_29 ? io_inData_41 : _GEN_1896; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1898 = 6'h2a == select_29 ? io_inData_42 : _GEN_1897; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1899 = 6'h2b == select_29 ? io_inData_43 : _GEN_1898; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1900 = 6'h2c == select_29 ? io_inData_44 : _GEN_1899; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1901 = 6'h2d == select_29 ? io_inData_45 : _GEN_1900; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1902 = 6'h2e == select_29 ? io_inData_46 : _GEN_1901; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1903 = 6'h2f == select_29 ? io_inData_47 : _GEN_1902; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1904 = 6'h30 == select_29 ? io_inData_48 : _GEN_1903; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1905 = 6'h31 == select_29 ? io_inData_49 : _GEN_1904; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1906 = 6'h32 == select_29 ? io_inData_50 : _GEN_1905; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1907 = 6'h33 == select_29 ? io_inData_51 : _GEN_1906; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1908 = 6'h34 == select_29 ? io_inData_52 : _GEN_1907; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1909 = 6'h35 == select_29 ? io_inData_53 : _GEN_1908; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1910 = 6'h36 == select_29 ? io_inData_54 : _GEN_1909; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1911 = 6'h37 == select_29 ? io_inData_55 : _GEN_1910; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1912 = 6'h38 == select_29 ? io_inData_56 : _GEN_1911; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1913 = 6'h39 == select_29 ? io_inData_57 : _GEN_1912; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1914 = 6'h3a == select_29 ? io_inData_58 : _GEN_1913; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1915 = 6'h3b == select_29 ? io_inData_59 : _GEN_1914; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1916 = 6'h3c == select_29 ? io_inData_60 : _GEN_1915; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1917 = 6'h3d == select_29 ? io_inData_61 : _GEN_1916; // @[Switch.scala 33:19:@9604.4]
  assign _GEN_1918 = 6'h3e == select_29 ? io_inData_62 : _GEN_1917; // @[Switch.scala 33:19:@9604.4]
  assign _T_29144 = {valid_29_7,valid_29_6,valid_29_5,valid_29_4,valid_29_3,valid_29_2,valid_29_1,valid_29_0}; // @[Switch.scala 34:32:@9611.4]
  assign _T_29152 = {valid_29_15,valid_29_14,valid_29_13,valid_29_12,valid_29_11,valid_29_10,valid_29_9,valid_29_8,_T_29144}; // @[Switch.scala 34:32:@9619.4]
  assign _T_29159 = {valid_29_23,valid_29_22,valid_29_21,valid_29_20,valid_29_19,valid_29_18,valid_29_17,valid_29_16}; // @[Switch.scala 34:32:@9626.4]
  assign _T_29168 = {valid_29_31,valid_29_30,valid_29_29,valid_29_28,valid_29_27,valid_29_26,valid_29_25,valid_29_24,_T_29159,_T_29152}; // @[Switch.scala 34:32:@9635.4]
  assign _T_29175 = {valid_29_39,valid_29_38,valid_29_37,valid_29_36,valid_29_35,valid_29_34,valid_29_33,valid_29_32}; // @[Switch.scala 34:32:@9642.4]
  assign _T_29183 = {valid_29_47,valid_29_46,valid_29_45,valid_29_44,valid_29_43,valid_29_42,valid_29_41,valid_29_40,_T_29175}; // @[Switch.scala 34:32:@9650.4]
  assign _T_29190 = {valid_29_55,valid_29_54,valid_29_53,valid_29_52,valid_29_51,valid_29_50,valid_29_49,valid_29_48}; // @[Switch.scala 34:32:@9657.4]
  assign _T_29199 = {valid_29_63,valid_29_62,valid_29_61,valid_29_60,valid_29_59,valid_29_58,valid_29_57,valid_29_56,_T_29190,_T_29183}; // @[Switch.scala 34:32:@9666.4]
  assign _T_29200 = {_T_29199,_T_29168}; // @[Switch.scala 34:32:@9667.4]
  assign _T_29204 = io_inAddr_0 == 6'h1e; // @[Switch.scala 30:53:@9670.4]
  assign valid_30_0 = io_inValid_0 & _T_29204; // @[Switch.scala 30:36:@9671.4]
  assign _T_29207 = io_inAddr_1 == 6'h1e; // @[Switch.scala 30:53:@9673.4]
  assign valid_30_1 = io_inValid_1 & _T_29207; // @[Switch.scala 30:36:@9674.4]
  assign _T_29210 = io_inAddr_2 == 6'h1e; // @[Switch.scala 30:53:@9676.4]
  assign valid_30_2 = io_inValid_2 & _T_29210; // @[Switch.scala 30:36:@9677.4]
  assign _T_29213 = io_inAddr_3 == 6'h1e; // @[Switch.scala 30:53:@9679.4]
  assign valid_30_3 = io_inValid_3 & _T_29213; // @[Switch.scala 30:36:@9680.4]
  assign _T_29216 = io_inAddr_4 == 6'h1e; // @[Switch.scala 30:53:@9682.4]
  assign valid_30_4 = io_inValid_4 & _T_29216; // @[Switch.scala 30:36:@9683.4]
  assign _T_29219 = io_inAddr_5 == 6'h1e; // @[Switch.scala 30:53:@9685.4]
  assign valid_30_5 = io_inValid_5 & _T_29219; // @[Switch.scala 30:36:@9686.4]
  assign _T_29222 = io_inAddr_6 == 6'h1e; // @[Switch.scala 30:53:@9688.4]
  assign valid_30_6 = io_inValid_6 & _T_29222; // @[Switch.scala 30:36:@9689.4]
  assign _T_29225 = io_inAddr_7 == 6'h1e; // @[Switch.scala 30:53:@9691.4]
  assign valid_30_7 = io_inValid_7 & _T_29225; // @[Switch.scala 30:36:@9692.4]
  assign _T_29228 = io_inAddr_8 == 6'h1e; // @[Switch.scala 30:53:@9694.4]
  assign valid_30_8 = io_inValid_8 & _T_29228; // @[Switch.scala 30:36:@9695.4]
  assign _T_29231 = io_inAddr_9 == 6'h1e; // @[Switch.scala 30:53:@9697.4]
  assign valid_30_9 = io_inValid_9 & _T_29231; // @[Switch.scala 30:36:@9698.4]
  assign _T_29234 = io_inAddr_10 == 6'h1e; // @[Switch.scala 30:53:@9700.4]
  assign valid_30_10 = io_inValid_10 & _T_29234; // @[Switch.scala 30:36:@9701.4]
  assign _T_29237 = io_inAddr_11 == 6'h1e; // @[Switch.scala 30:53:@9703.4]
  assign valid_30_11 = io_inValid_11 & _T_29237; // @[Switch.scala 30:36:@9704.4]
  assign _T_29240 = io_inAddr_12 == 6'h1e; // @[Switch.scala 30:53:@9706.4]
  assign valid_30_12 = io_inValid_12 & _T_29240; // @[Switch.scala 30:36:@9707.4]
  assign _T_29243 = io_inAddr_13 == 6'h1e; // @[Switch.scala 30:53:@9709.4]
  assign valid_30_13 = io_inValid_13 & _T_29243; // @[Switch.scala 30:36:@9710.4]
  assign _T_29246 = io_inAddr_14 == 6'h1e; // @[Switch.scala 30:53:@9712.4]
  assign valid_30_14 = io_inValid_14 & _T_29246; // @[Switch.scala 30:36:@9713.4]
  assign _T_29249 = io_inAddr_15 == 6'h1e; // @[Switch.scala 30:53:@9715.4]
  assign valid_30_15 = io_inValid_15 & _T_29249; // @[Switch.scala 30:36:@9716.4]
  assign _T_29252 = io_inAddr_16 == 6'h1e; // @[Switch.scala 30:53:@9718.4]
  assign valid_30_16 = io_inValid_16 & _T_29252; // @[Switch.scala 30:36:@9719.4]
  assign _T_29255 = io_inAddr_17 == 6'h1e; // @[Switch.scala 30:53:@9721.4]
  assign valid_30_17 = io_inValid_17 & _T_29255; // @[Switch.scala 30:36:@9722.4]
  assign _T_29258 = io_inAddr_18 == 6'h1e; // @[Switch.scala 30:53:@9724.4]
  assign valid_30_18 = io_inValid_18 & _T_29258; // @[Switch.scala 30:36:@9725.4]
  assign _T_29261 = io_inAddr_19 == 6'h1e; // @[Switch.scala 30:53:@9727.4]
  assign valid_30_19 = io_inValid_19 & _T_29261; // @[Switch.scala 30:36:@9728.4]
  assign _T_29264 = io_inAddr_20 == 6'h1e; // @[Switch.scala 30:53:@9730.4]
  assign valid_30_20 = io_inValid_20 & _T_29264; // @[Switch.scala 30:36:@9731.4]
  assign _T_29267 = io_inAddr_21 == 6'h1e; // @[Switch.scala 30:53:@9733.4]
  assign valid_30_21 = io_inValid_21 & _T_29267; // @[Switch.scala 30:36:@9734.4]
  assign _T_29270 = io_inAddr_22 == 6'h1e; // @[Switch.scala 30:53:@9736.4]
  assign valid_30_22 = io_inValid_22 & _T_29270; // @[Switch.scala 30:36:@9737.4]
  assign _T_29273 = io_inAddr_23 == 6'h1e; // @[Switch.scala 30:53:@9739.4]
  assign valid_30_23 = io_inValid_23 & _T_29273; // @[Switch.scala 30:36:@9740.4]
  assign _T_29276 = io_inAddr_24 == 6'h1e; // @[Switch.scala 30:53:@9742.4]
  assign valid_30_24 = io_inValid_24 & _T_29276; // @[Switch.scala 30:36:@9743.4]
  assign _T_29279 = io_inAddr_25 == 6'h1e; // @[Switch.scala 30:53:@9745.4]
  assign valid_30_25 = io_inValid_25 & _T_29279; // @[Switch.scala 30:36:@9746.4]
  assign _T_29282 = io_inAddr_26 == 6'h1e; // @[Switch.scala 30:53:@9748.4]
  assign valid_30_26 = io_inValid_26 & _T_29282; // @[Switch.scala 30:36:@9749.4]
  assign _T_29285 = io_inAddr_27 == 6'h1e; // @[Switch.scala 30:53:@9751.4]
  assign valid_30_27 = io_inValid_27 & _T_29285; // @[Switch.scala 30:36:@9752.4]
  assign _T_29288 = io_inAddr_28 == 6'h1e; // @[Switch.scala 30:53:@9754.4]
  assign valid_30_28 = io_inValid_28 & _T_29288; // @[Switch.scala 30:36:@9755.4]
  assign _T_29291 = io_inAddr_29 == 6'h1e; // @[Switch.scala 30:53:@9757.4]
  assign valid_30_29 = io_inValid_29 & _T_29291; // @[Switch.scala 30:36:@9758.4]
  assign _T_29294 = io_inAddr_30 == 6'h1e; // @[Switch.scala 30:53:@9760.4]
  assign valid_30_30 = io_inValid_30 & _T_29294; // @[Switch.scala 30:36:@9761.4]
  assign _T_29297 = io_inAddr_31 == 6'h1e; // @[Switch.scala 30:53:@9763.4]
  assign valid_30_31 = io_inValid_31 & _T_29297; // @[Switch.scala 30:36:@9764.4]
  assign _T_29300 = io_inAddr_32 == 6'h1e; // @[Switch.scala 30:53:@9766.4]
  assign valid_30_32 = io_inValid_32 & _T_29300; // @[Switch.scala 30:36:@9767.4]
  assign _T_29303 = io_inAddr_33 == 6'h1e; // @[Switch.scala 30:53:@9769.4]
  assign valid_30_33 = io_inValid_33 & _T_29303; // @[Switch.scala 30:36:@9770.4]
  assign _T_29306 = io_inAddr_34 == 6'h1e; // @[Switch.scala 30:53:@9772.4]
  assign valid_30_34 = io_inValid_34 & _T_29306; // @[Switch.scala 30:36:@9773.4]
  assign _T_29309 = io_inAddr_35 == 6'h1e; // @[Switch.scala 30:53:@9775.4]
  assign valid_30_35 = io_inValid_35 & _T_29309; // @[Switch.scala 30:36:@9776.4]
  assign _T_29312 = io_inAddr_36 == 6'h1e; // @[Switch.scala 30:53:@9778.4]
  assign valid_30_36 = io_inValid_36 & _T_29312; // @[Switch.scala 30:36:@9779.4]
  assign _T_29315 = io_inAddr_37 == 6'h1e; // @[Switch.scala 30:53:@9781.4]
  assign valid_30_37 = io_inValid_37 & _T_29315; // @[Switch.scala 30:36:@9782.4]
  assign _T_29318 = io_inAddr_38 == 6'h1e; // @[Switch.scala 30:53:@9784.4]
  assign valid_30_38 = io_inValid_38 & _T_29318; // @[Switch.scala 30:36:@9785.4]
  assign _T_29321 = io_inAddr_39 == 6'h1e; // @[Switch.scala 30:53:@9787.4]
  assign valid_30_39 = io_inValid_39 & _T_29321; // @[Switch.scala 30:36:@9788.4]
  assign _T_29324 = io_inAddr_40 == 6'h1e; // @[Switch.scala 30:53:@9790.4]
  assign valid_30_40 = io_inValid_40 & _T_29324; // @[Switch.scala 30:36:@9791.4]
  assign _T_29327 = io_inAddr_41 == 6'h1e; // @[Switch.scala 30:53:@9793.4]
  assign valid_30_41 = io_inValid_41 & _T_29327; // @[Switch.scala 30:36:@9794.4]
  assign _T_29330 = io_inAddr_42 == 6'h1e; // @[Switch.scala 30:53:@9796.4]
  assign valid_30_42 = io_inValid_42 & _T_29330; // @[Switch.scala 30:36:@9797.4]
  assign _T_29333 = io_inAddr_43 == 6'h1e; // @[Switch.scala 30:53:@9799.4]
  assign valid_30_43 = io_inValid_43 & _T_29333; // @[Switch.scala 30:36:@9800.4]
  assign _T_29336 = io_inAddr_44 == 6'h1e; // @[Switch.scala 30:53:@9802.4]
  assign valid_30_44 = io_inValid_44 & _T_29336; // @[Switch.scala 30:36:@9803.4]
  assign _T_29339 = io_inAddr_45 == 6'h1e; // @[Switch.scala 30:53:@9805.4]
  assign valid_30_45 = io_inValid_45 & _T_29339; // @[Switch.scala 30:36:@9806.4]
  assign _T_29342 = io_inAddr_46 == 6'h1e; // @[Switch.scala 30:53:@9808.4]
  assign valid_30_46 = io_inValid_46 & _T_29342; // @[Switch.scala 30:36:@9809.4]
  assign _T_29345 = io_inAddr_47 == 6'h1e; // @[Switch.scala 30:53:@9811.4]
  assign valid_30_47 = io_inValid_47 & _T_29345; // @[Switch.scala 30:36:@9812.4]
  assign _T_29348 = io_inAddr_48 == 6'h1e; // @[Switch.scala 30:53:@9814.4]
  assign valid_30_48 = io_inValid_48 & _T_29348; // @[Switch.scala 30:36:@9815.4]
  assign _T_29351 = io_inAddr_49 == 6'h1e; // @[Switch.scala 30:53:@9817.4]
  assign valid_30_49 = io_inValid_49 & _T_29351; // @[Switch.scala 30:36:@9818.4]
  assign _T_29354 = io_inAddr_50 == 6'h1e; // @[Switch.scala 30:53:@9820.4]
  assign valid_30_50 = io_inValid_50 & _T_29354; // @[Switch.scala 30:36:@9821.4]
  assign _T_29357 = io_inAddr_51 == 6'h1e; // @[Switch.scala 30:53:@9823.4]
  assign valid_30_51 = io_inValid_51 & _T_29357; // @[Switch.scala 30:36:@9824.4]
  assign _T_29360 = io_inAddr_52 == 6'h1e; // @[Switch.scala 30:53:@9826.4]
  assign valid_30_52 = io_inValid_52 & _T_29360; // @[Switch.scala 30:36:@9827.4]
  assign _T_29363 = io_inAddr_53 == 6'h1e; // @[Switch.scala 30:53:@9829.4]
  assign valid_30_53 = io_inValid_53 & _T_29363; // @[Switch.scala 30:36:@9830.4]
  assign _T_29366 = io_inAddr_54 == 6'h1e; // @[Switch.scala 30:53:@9832.4]
  assign valid_30_54 = io_inValid_54 & _T_29366; // @[Switch.scala 30:36:@9833.4]
  assign _T_29369 = io_inAddr_55 == 6'h1e; // @[Switch.scala 30:53:@9835.4]
  assign valid_30_55 = io_inValid_55 & _T_29369; // @[Switch.scala 30:36:@9836.4]
  assign _T_29372 = io_inAddr_56 == 6'h1e; // @[Switch.scala 30:53:@9838.4]
  assign valid_30_56 = io_inValid_56 & _T_29372; // @[Switch.scala 30:36:@9839.4]
  assign _T_29375 = io_inAddr_57 == 6'h1e; // @[Switch.scala 30:53:@9841.4]
  assign valid_30_57 = io_inValid_57 & _T_29375; // @[Switch.scala 30:36:@9842.4]
  assign _T_29378 = io_inAddr_58 == 6'h1e; // @[Switch.scala 30:53:@9844.4]
  assign valid_30_58 = io_inValid_58 & _T_29378; // @[Switch.scala 30:36:@9845.4]
  assign _T_29381 = io_inAddr_59 == 6'h1e; // @[Switch.scala 30:53:@9847.4]
  assign valid_30_59 = io_inValid_59 & _T_29381; // @[Switch.scala 30:36:@9848.4]
  assign _T_29384 = io_inAddr_60 == 6'h1e; // @[Switch.scala 30:53:@9850.4]
  assign valid_30_60 = io_inValid_60 & _T_29384; // @[Switch.scala 30:36:@9851.4]
  assign _T_29387 = io_inAddr_61 == 6'h1e; // @[Switch.scala 30:53:@9853.4]
  assign valid_30_61 = io_inValid_61 & _T_29387; // @[Switch.scala 30:36:@9854.4]
  assign _T_29390 = io_inAddr_62 == 6'h1e; // @[Switch.scala 30:53:@9856.4]
  assign valid_30_62 = io_inValid_62 & _T_29390; // @[Switch.scala 30:36:@9857.4]
  assign _T_29393 = io_inAddr_63 == 6'h1e; // @[Switch.scala 30:53:@9859.4]
  assign valid_30_63 = io_inValid_63 & _T_29393; // @[Switch.scala 30:36:@9860.4]
  assign _T_29459 = valid_30_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@9862.4]
  assign _T_29460 = valid_30_61 ? 6'h3d : _T_29459; // @[Mux.scala 31:69:@9863.4]
  assign _T_29461 = valid_30_60 ? 6'h3c : _T_29460; // @[Mux.scala 31:69:@9864.4]
  assign _T_29462 = valid_30_59 ? 6'h3b : _T_29461; // @[Mux.scala 31:69:@9865.4]
  assign _T_29463 = valid_30_58 ? 6'h3a : _T_29462; // @[Mux.scala 31:69:@9866.4]
  assign _T_29464 = valid_30_57 ? 6'h39 : _T_29463; // @[Mux.scala 31:69:@9867.4]
  assign _T_29465 = valid_30_56 ? 6'h38 : _T_29464; // @[Mux.scala 31:69:@9868.4]
  assign _T_29466 = valid_30_55 ? 6'h37 : _T_29465; // @[Mux.scala 31:69:@9869.4]
  assign _T_29467 = valid_30_54 ? 6'h36 : _T_29466; // @[Mux.scala 31:69:@9870.4]
  assign _T_29468 = valid_30_53 ? 6'h35 : _T_29467; // @[Mux.scala 31:69:@9871.4]
  assign _T_29469 = valid_30_52 ? 6'h34 : _T_29468; // @[Mux.scala 31:69:@9872.4]
  assign _T_29470 = valid_30_51 ? 6'h33 : _T_29469; // @[Mux.scala 31:69:@9873.4]
  assign _T_29471 = valid_30_50 ? 6'h32 : _T_29470; // @[Mux.scala 31:69:@9874.4]
  assign _T_29472 = valid_30_49 ? 6'h31 : _T_29471; // @[Mux.scala 31:69:@9875.4]
  assign _T_29473 = valid_30_48 ? 6'h30 : _T_29472; // @[Mux.scala 31:69:@9876.4]
  assign _T_29474 = valid_30_47 ? 6'h2f : _T_29473; // @[Mux.scala 31:69:@9877.4]
  assign _T_29475 = valid_30_46 ? 6'h2e : _T_29474; // @[Mux.scala 31:69:@9878.4]
  assign _T_29476 = valid_30_45 ? 6'h2d : _T_29475; // @[Mux.scala 31:69:@9879.4]
  assign _T_29477 = valid_30_44 ? 6'h2c : _T_29476; // @[Mux.scala 31:69:@9880.4]
  assign _T_29478 = valid_30_43 ? 6'h2b : _T_29477; // @[Mux.scala 31:69:@9881.4]
  assign _T_29479 = valid_30_42 ? 6'h2a : _T_29478; // @[Mux.scala 31:69:@9882.4]
  assign _T_29480 = valid_30_41 ? 6'h29 : _T_29479; // @[Mux.scala 31:69:@9883.4]
  assign _T_29481 = valid_30_40 ? 6'h28 : _T_29480; // @[Mux.scala 31:69:@9884.4]
  assign _T_29482 = valid_30_39 ? 6'h27 : _T_29481; // @[Mux.scala 31:69:@9885.4]
  assign _T_29483 = valid_30_38 ? 6'h26 : _T_29482; // @[Mux.scala 31:69:@9886.4]
  assign _T_29484 = valid_30_37 ? 6'h25 : _T_29483; // @[Mux.scala 31:69:@9887.4]
  assign _T_29485 = valid_30_36 ? 6'h24 : _T_29484; // @[Mux.scala 31:69:@9888.4]
  assign _T_29486 = valid_30_35 ? 6'h23 : _T_29485; // @[Mux.scala 31:69:@9889.4]
  assign _T_29487 = valid_30_34 ? 6'h22 : _T_29486; // @[Mux.scala 31:69:@9890.4]
  assign _T_29488 = valid_30_33 ? 6'h21 : _T_29487; // @[Mux.scala 31:69:@9891.4]
  assign _T_29489 = valid_30_32 ? 6'h20 : _T_29488; // @[Mux.scala 31:69:@9892.4]
  assign _T_29490 = valid_30_31 ? 6'h1f : _T_29489; // @[Mux.scala 31:69:@9893.4]
  assign _T_29491 = valid_30_30 ? 6'h1e : _T_29490; // @[Mux.scala 31:69:@9894.4]
  assign _T_29492 = valid_30_29 ? 6'h1d : _T_29491; // @[Mux.scala 31:69:@9895.4]
  assign _T_29493 = valid_30_28 ? 6'h1c : _T_29492; // @[Mux.scala 31:69:@9896.4]
  assign _T_29494 = valid_30_27 ? 6'h1b : _T_29493; // @[Mux.scala 31:69:@9897.4]
  assign _T_29495 = valid_30_26 ? 6'h1a : _T_29494; // @[Mux.scala 31:69:@9898.4]
  assign _T_29496 = valid_30_25 ? 6'h19 : _T_29495; // @[Mux.scala 31:69:@9899.4]
  assign _T_29497 = valid_30_24 ? 6'h18 : _T_29496; // @[Mux.scala 31:69:@9900.4]
  assign _T_29498 = valid_30_23 ? 6'h17 : _T_29497; // @[Mux.scala 31:69:@9901.4]
  assign _T_29499 = valid_30_22 ? 6'h16 : _T_29498; // @[Mux.scala 31:69:@9902.4]
  assign _T_29500 = valid_30_21 ? 6'h15 : _T_29499; // @[Mux.scala 31:69:@9903.4]
  assign _T_29501 = valid_30_20 ? 6'h14 : _T_29500; // @[Mux.scala 31:69:@9904.4]
  assign _T_29502 = valid_30_19 ? 6'h13 : _T_29501; // @[Mux.scala 31:69:@9905.4]
  assign _T_29503 = valid_30_18 ? 6'h12 : _T_29502; // @[Mux.scala 31:69:@9906.4]
  assign _T_29504 = valid_30_17 ? 6'h11 : _T_29503; // @[Mux.scala 31:69:@9907.4]
  assign _T_29505 = valid_30_16 ? 6'h10 : _T_29504; // @[Mux.scala 31:69:@9908.4]
  assign _T_29506 = valid_30_15 ? 6'hf : _T_29505; // @[Mux.scala 31:69:@9909.4]
  assign _T_29507 = valid_30_14 ? 6'he : _T_29506; // @[Mux.scala 31:69:@9910.4]
  assign _T_29508 = valid_30_13 ? 6'hd : _T_29507; // @[Mux.scala 31:69:@9911.4]
  assign _T_29509 = valid_30_12 ? 6'hc : _T_29508; // @[Mux.scala 31:69:@9912.4]
  assign _T_29510 = valid_30_11 ? 6'hb : _T_29509; // @[Mux.scala 31:69:@9913.4]
  assign _T_29511 = valid_30_10 ? 6'ha : _T_29510; // @[Mux.scala 31:69:@9914.4]
  assign _T_29512 = valid_30_9 ? 6'h9 : _T_29511; // @[Mux.scala 31:69:@9915.4]
  assign _T_29513 = valid_30_8 ? 6'h8 : _T_29512; // @[Mux.scala 31:69:@9916.4]
  assign _T_29514 = valid_30_7 ? 6'h7 : _T_29513; // @[Mux.scala 31:69:@9917.4]
  assign _T_29515 = valid_30_6 ? 6'h6 : _T_29514; // @[Mux.scala 31:69:@9918.4]
  assign _T_29516 = valid_30_5 ? 6'h5 : _T_29515; // @[Mux.scala 31:69:@9919.4]
  assign _T_29517 = valid_30_4 ? 6'h4 : _T_29516; // @[Mux.scala 31:69:@9920.4]
  assign _T_29518 = valid_30_3 ? 6'h3 : _T_29517; // @[Mux.scala 31:69:@9921.4]
  assign _T_29519 = valid_30_2 ? 6'h2 : _T_29518; // @[Mux.scala 31:69:@9922.4]
  assign _T_29520 = valid_30_1 ? 6'h1 : _T_29519; // @[Mux.scala 31:69:@9923.4]
  assign select_30 = valid_30_0 ? 6'h0 : _T_29520; // @[Mux.scala 31:69:@9924.4]
  assign _GEN_1921 = 6'h1 == select_30 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1922 = 6'h2 == select_30 ? io_inData_2 : _GEN_1921; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1923 = 6'h3 == select_30 ? io_inData_3 : _GEN_1922; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1924 = 6'h4 == select_30 ? io_inData_4 : _GEN_1923; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1925 = 6'h5 == select_30 ? io_inData_5 : _GEN_1924; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1926 = 6'h6 == select_30 ? io_inData_6 : _GEN_1925; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1927 = 6'h7 == select_30 ? io_inData_7 : _GEN_1926; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1928 = 6'h8 == select_30 ? io_inData_8 : _GEN_1927; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1929 = 6'h9 == select_30 ? io_inData_9 : _GEN_1928; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1930 = 6'ha == select_30 ? io_inData_10 : _GEN_1929; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1931 = 6'hb == select_30 ? io_inData_11 : _GEN_1930; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1932 = 6'hc == select_30 ? io_inData_12 : _GEN_1931; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1933 = 6'hd == select_30 ? io_inData_13 : _GEN_1932; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1934 = 6'he == select_30 ? io_inData_14 : _GEN_1933; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1935 = 6'hf == select_30 ? io_inData_15 : _GEN_1934; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1936 = 6'h10 == select_30 ? io_inData_16 : _GEN_1935; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1937 = 6'h11 == select_30 ? io_inData_17 : _GEN_1936; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1938 = 6'h12 == select_30 ? io_inData_18 : _GEN_1937; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1939 = 6'h13 == select_30 ? io_inData_19 : _GEN_1938; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1940 = 6'h14 == select_30 ? io_inData_20 : _GEN_1939; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1941 = 6'h15 == select_30 ? io_inData_21 : _GEN_1940; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1942 = 6'h16 == select_30 ? io_inData_22 : _GEN_1941; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1943 = 6'h17 == select_30 ? io_inData_23 : _GEN_1942; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1944 = 6'h18 == select_30 ? io_inData_24 : _GEN_1943; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1945 = 6'h19 == select_30 ? io_inData_25 : _GEN_1944; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1946 = 6'h1a == select_30 ? io_inData_26 : _GEN_1945; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1947 = 6'h1b == select_30 ? io_inData_27 : _GEN_1946; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1948 = 6'h1c == select_30 ? io_inData_28 : _GEN_1947; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1949 = 6'h1d == select_30 ? io_inData_29 : _GEN_1948; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1950 = 6'h1e == select_30 ? io_inData_30 : _GEN_1949; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1951 = 6'h1f == select_30 ? io_inData_31 : _GEN_1950; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1952 = 6'h20 == select_30 ? io_inData_32 : _GEN_1951; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1953 = 6'h21 == select_30 ? io_inData_33 : _GEN_1952; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1954 = 6'h22 == select_30 ? io_inData_34 : _GEN_1953; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1955 = 6'h23 == select_30 ? io_inData_35 : _GEN_1954; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1956 = 6'h24 == select_30 ? io_inData_36 : _GEN_1955; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1957 = 6'h25 == select_30 ? io_inData_37 : _GEN_1956; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1958 = 6'h26 == select_30 ? io_inData_38 : _GEN_1957; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1959 = 6'h27 == select_30 ? io_inData_39 : _GEN_1958; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1960 = 6'h28 == select_30 ? io_inData_40 : _GEN_1959; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1961 = 6'h29 == select_30 ? io_inData_41 : _GEN_1960; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1962 = 6'h2a == select_30 ? io_inData_42 : _GEN_1961; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1963 = 6'h2b == select_30 ? io_inData_43 : _GEN_1962; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1964 = 6'h2c == select_30 ? io_inData_44 : _GEN_1963; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1965 = 6'h2d == select_30 ? io_inData_45 : _GEN_1964; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1966 = 6'h2e == select_30 ? io_inData_46 : _GEN_1965; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1967 = 6'h2f == select_30 ? io_inData_47 : _GEN_1966; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1968 = 6'h30 == select_30 ? io_inData_48 : _GEN_1967; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1969 = 6'h31 == select_30 ? io_inData_49 : _GEN_1968; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1970 = 6'h32 == select_30 ? io_inData_50 : _GEN_1969; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1971 = 6'h33 == select_30 ? io_inData_51 : _GEN_1970; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1972 = 6'h34 == select_30 ? io_inData_52 : _GEN_1971; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1973 = 6'h35 == select_30 ? io_inData_53 : _GEN_1972; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1974 = 6'h36 == select_30 ? io_inData_54 : _GEN_1973; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1975 = 6'h37 == select_30 ? io_inData_55 : _GEN_1974; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1976 = 6'h38 == select_30 ? io_inData_56 : _GEN_1975; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1977 = 6'h39 == select_30 ? io_inData_57 : _GEN_1976; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1978 = 6'h3a == select_30 ? io_inData_58 : _GEN_1977; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1979 = 6'h3b == select_30 ? io_inData_59 : _GEN_1978; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1980 = 6'h3c == select_30 ? io_inData_60 : _GEN_1979; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1981 = 6'h3d == select_30 ? io_inData_61 : _GEN_1980; // @[Switch.scala 33:19:@9926.4]
  assign _GEN_1982 = 6'h3e == select_30 ? io_inData_62 : _GEN_1981; // @[Switch.scala 33:19:@9926.4]
  assign _T_29529 = {valid_30_7,valid_30_6,valid_30_5,valid_30_4,valid_30_3,valid_30_2,valid_30_1,valid_30_0}; // @[Switch.scala 34:32:@9933.4]
  assign _T_29537 = {valid_30_15,valid_30_14,valid_30_13,valid_30_12,valid_30_11,valid_30_10,valid_30_9,valid_30_8,_T_29529}; // @[Switch.scala 34:32:@9941.4]
  assign _T_29544 = {valid_30_23,valid_30_22,valid_30_21,valid_30_20,valid_30_19,valid_30_18,valid_30_17,valid_30_16}; // @[Switch.scala 34:32:@9948.4]
  assign _T_29553 = {valid_30_31,valid_30_30,valid_30_29,valid_30_28,valid_30_27,valid_30_26,valid_30_25,valid_30_24,_T_29544,_T_29537}; // @[Switch.scala 34:32:@9957.4]
  assign _T_29560 = {valid_30_39,valid_30_38,valid_30_37,valid_30_36,valid_30_35,valid_30_34,valid_30_33,valid_30_32}; // @[Switch.scala 34:32:@9964.4]
  assign _T_29568 = {valid_30_47,valid_30_46,valid_30_45,valid_30_44,valid_30_43,valid_30_42,valid_30_41,valid_30_40,_T_29560}; // @[Switch.scala 34:32:@9972.4]
  assign _T_29575 = {valid_30_55,valid_30_54,valid_30_53,valid_30_52,valid_30_51,valid_30_50,valid_30_49,valid_30_48}; // @[Switch.scala 34:32:@9979.4]
  assign _T_29584 = {valid_30_63,valid_30_62,valid_30_61,valid_30_60,valid_30_59,valid_30_58,valid_30_57,valid_30_56,_T_29575,_T_29568}; // @[Switch.scala 34:32:@9988.4]
  assign _T_29585 = {_T_29584,_T_29553}; // @[Switch.scala 34:32:@9989.4]
  assign _T_29589 = io_inAddr_0 == 6'h1f; // @[Switch.scala 30:53:@9992.4]
  assign valid_31_0 = io_inValid_0 & _T_29589; // @[Switch.scala 30:36:@9993.4]
  assign _T_29592 = io_inAddr_1 == 6'h1f; // @[Switch.scala 30:53:@9995.4]
  assign valid_31_1 = io_inValid_1 & _T_29592; // @[Switch.scala 30:36:@9996.4]
  assign _T_29595 = io_inAddr_2 == 6'h1f; // @[Switch.scala 30:53:@9998.4]
  assign valid_31_2 = io_inValid_2 & _T_29595; // @[Switch.scala 30:36:@9999.4]
  assign _T_29598 = io_inAddr_3 == 6'h1f; // @[Switch.scala 30:53:@10001.4]
  assign valid_31_3 = io_inValid_3 & _T_29598; // @[Switch.scala 30:36:@10002.4]
  assign _T_29601 = io_inAddr_4 == 6'h1f; // @[Switch.scala 30:53:@10004.4]
  assign valid_31_4 = io_inValid_4 & _T_29601; // @[Switch.scala 30:36:@10005.4]
  assign _T_29604 = io_inAddr_5 == 6'h1f; // @[Switch.scala 30:53:@10007.4]
  assign valid_31_5 = io_inValid_5 & _T_29604; // @[Switch.scala 30:36:@10008.4]
  assign _T_29607 = io_inAddr_6 == 6'h1f; // @[Switch.scala 30:53:@10010.4]
  assign valid_31_6 = io_inValid_6 & _T_29607; // @[Switch.scala 30:36:@10011.4]
  assign _T_29610 = io_inAddr_7 == 6'h1f; // @[Switch.scala 30:53:@10013.4]
  assign valid_31_7 = io_inValid_7 & _T_29610; // @[Switch.scala 30:36:@10014.4]
  assign _T_29613 = io_inAddr_8 == 6'h1f; // @[Switch.scala 30:53:@10016.4]
  assign valid_31_8 = io_inValid_8 & _T_29613; // @[Switch.scala 30:36:@10017.4]
  assign _T_29616 = io_inAddr_9 == 6'h1f; // @[Switch.scala 30:53:@10019.4]
  assign valid_31_9 = io_inValid_9 & _T_29616; // @[Switch.scala 30:36:@10020.4]
  assign _T_29619 = io_inAddr_10 == 6'h1f; // @[Switch.scala 30:53:@10022.4]
  assign valid_31_10 = io_inValid_10 & _T_29619; // @[Switch.scala 30:36:@10023.4]
  assign _T_29622 = io_inAddr_11 == 6'h1f; // @[Switch.scala 30:53:@10025.4]
  assign valid_31_11 = io_inValid_11 & _T_29622; // @[Switch.scala 30:36:@10026.4]
  assign _T_29625 = io_inAddr_12 == 6'h1f; // @[Switch.scala 30:53:@10028.4]
  assign valid_31_12 = io_inValid_12 & _T_29625; // @[Switch.scala 30:36:@10029.4]
  assign _T_29628 = io_inAddr_13 == 6'h1f; // @[Switch.scala 30:53:@10031.4]
  assign valid_31_13 = io_inValid_13 & _T_29628; // @[Switch.scala 30:36:@10032.4]
  assign _T_29631 = io_inAddr_14 == 6'h1f; // @[Switch.scala 30:53:@10034.4]
  assign valid_31_14 = io_inValid_14 & _T_29631; // @[Switch.scala 30:36:@10035.4]
  assign _T_29634 = io_inAddr_15 == 6'h1f; // @[Switch.scala 30:53:@10037.4]
  assign valid_31_15 = io_inValid_15 & _T_29634; // @[Switch.scala 30:36:@10038.4]
  assign _T_29637 = io_inAddr_16 == 6'h1f; // @[Switch.scala 30:53:@10040.4]
  assign valid_31_16 = io_inValid_16 & _T_29637; // @[Switch.scala 30:36:@10041.4]
  assign _T_29640 = io_inAddr_17 == 6'h1f; // @[Switch.scala 30:53:@10043.4]
  assign valid_31_17 = io_inValid_17 & _T_29640; // @[Switch.scala 30:36:@10044.4]
  assign _T_29643 = io_inAddr_18 == 6'h1f; // @[Switch.scala 30:53:@10046.4]
  assign valid_31_18 = io_inValid_18 & _T_29643; // @[Switch.scala 30:36:@10047.4]
  assign _T_29646 = io_inAddr_19 == 6'h1f; // @[Switch.scala 30:53:@10049.4]
  assign valid_31_19 = io_inValid_19 & _T_29646; // @[Switch.scala 30:36:@10050.4]
  assign _T_29649 = io_inAddr_20 == 6'h1f; // @[Switch.scala 30:53:@10052.4]
  assign valid_31_20 = io_inValid_20 & _T_29649; // @[Switch.scala 30:36:@10053.4]
  assign _T_29652 = io_inAddr_21 == 6'h1f; // @[Switch.scala 30:53:@10055.4]
  assign valid_31_21 = io_inValid_21 & _T_29652; // @[Switch.scala 30:36:@10056.4]
  assign _T_29655 = io_inAddr_22 == 6'h1f; // @[Switch.scala 30:53:@10058.4]
  assign valid_31_22 = io_inValid_22 & _T_29655; // @[Switch.scala 30:36:@10059.4]
  assign _T_29658 = io_inAddr_23 == 6'h1f; // @[Switch.scala 30:53:@10061.4]
  assign valid_31_23 = io_inValid_23 & _T_29658; // @[Switch.scala 30:36:@10062.4]
  assign _T_29661 = io_inAddr_24 == 6'h1f; // @[Switch.scala 30:53:@10064.4]
  assign valid_31_24 = io_inValid_24 & _T_29661; // @[Switch.scala 30:36:@10065.4]
  assign _T_29664 = io_inAddr_25 == 6'h1f; // @[Switch.scala 30:53:@10067.4]
  assign valid_31_25 = io_inValid_25 & _T_29664; // @[Switch.scala 30:36:@10068.4]
  assign _T_29667 = io_inAddr_26 == 6'h1f; // @[Switch.scala 30:53:@10070.4]
  assign valid_31_26 = io_inValid_26 & _T_29667; // @[Switch.scala 30:36:@10071.4]
  assign _T_29670 = io_inAddr_27 == 6'h1f; // @[Switch.scala 30:53:@10073.4]
  assign valid_31_27 = io_inValid_27 & _T_29670; // @[Switch.scala 30:36:@10074.4]
  assign _T_29673 = io_inAddr_28 == 6'h1f; // @[Switch.scala 30:53:@10076.4]
  assign valid_31_28 = io_inValid_28 & _T_29673; // @[Switch.scala 30:36:@10077.4]
  assign _T_29676 = io_inAddr_29 == 6'h1f; // @[Switch.scala 30:53:@10079.4]
  assign valid_31_29 = io_inValid_29 & _T_29676; // @[Switch.scala 30:36:@10080.4]
  assign _T_29679 = io_inAddr_30 == 6'h1f; // @[Switch.scala 30:53:@10082.4]
  assign valid_31_30 = io_inValid_30 & _T_29679; // @[Switch.scala 30:36:@10083.4]
  assign _T_29682 = io_inAddr_31 == 6'h1f; // @[Switch.scala 30:53:@10085.4]
  assign valid_31_31 = io_inValid_31 & _T_29682; // @[Switch.scala 30:36:@10086.4]
  assign _T_29685 = io_inAddr_32 == 6'h1f; // @[Switch.scala 30:53:@10088.4]
  assign valid_31_32 = io_inValid_32 & _T_29685; // @[Switch.scala 30:36:@10089.4]
  assign _T_29688 = io_inAddr_33 == 6'h1f; // @[Switch.scala 30:53:@10091.4]
  assign valid_31_33 = io_inValid_33 & _T_29688; // @[Switch.scala 30:36:@10092.4]
  assign _T_29691 = io_inAddr_34 == 6'h1f; // @[Switch.scala 30:53:@10094.4]
  assign valid_31_34 = io_inValid_34 & _T_29691; // @[Switch.scala 30:36:@10095.4]
  assign _T_29694 = io_inAddr_35 == 6'h1f; // @[Switch.scala 30:53:@10097.4]
  assign valid_31_35 = io_inValid_35 & _T_29694; // @[Switch.scala 30:36:@10098.4]
  assign _T_29697 = io_inAddr_36 == 6'h1f; // @[Switch.scala 30:53:@10100.4]
  assign valid_31_36 = io_inValid_36 & _T_29697; // @[Switch.scala 30:36:@10101.4]
  assign _T_29700 = io_inAddr_37 == 6'h1f; // @[Switch.scala 30:53:@10103.4]
  assign valid_31_37 = io_inValid_37 & _T_29700; // @[Switch.scala 30:36:@10104.4]
  assign _T_29703 = io_inAddr_38 == 6'h1f; // @[Switch.scala 30:53:@10106.4]
  assign valid_31_38 = io_inValid_38 & _T_29703; // @[Switch.scala 30:36:@10107.4]
  assign _T_29706 = io_inAddr_39 == 6'h1f; // @[Switch.scala 30:53:@10109.4]
  assign valid_31_39 = io_inValid_39 & _T_29706; // @[Switch.scala 30:36:@10110.4]
  assign _T_29709 = io_inAddr_40 == 6'h1f; // @[Switch.scala 30:53:@10112.4]
  assign valid_31_40 = io_inValid_40 & _T_29709; // @[Switch.scala 30:36:@10113.4]
  assign _T_29712 = io_inAddr_41 == 6'h1f; // @[Switch.scala 30:53:@10115.4]
  assign valid_31_41 = io_inValid_41 & _T_29712; // @[Switch.scala 30:36:@10116.4]
  assign _T_29715 = io_inAddr_42 == 6'h1f; // @[Switch.scala 30:53:@10118.4]
  assign valid_31_42 = io_inValid_42 & _T_29715; // @[Switch.scala 30:36:@10119.4]
  assign _T_29718 = io_inAddr_43 == 6'h1f; // @[Switch.scala 30:53:@10121.4]
  assign valid_31_43 = io_inValid_43 & _T_29718; // @[Switch.scala 30:36:@10122.4]
  assign _T_29721 = io_inAddr_44 == 6'h1f; // @[Switch.scala 30:53:@10124.4]
  assign valid_31_44 = io_inValid_44 & _T_29721; // @[Switch.scala 30:36:@10125.4]
  assign _T_29724 = io_inAddr_45 == 6'h1f; // @[Switch.scala 30:53:@10127.4]
  assign valid_31_45 = io_inValid_45 & _T_29724; // @[Switch.scala 30:36:@10128.4]
  assign _T_29727 = io_inAddr_46 == 6'h1f; // @[Switch.scala 30:53:@10130.4]
  assign valid_31_46 = io_inValid_46 & _T_29727; // @[Switch.scala 30:36:@10131.4]
  assign _T_29730 = io_inAddr_47 == 6'h1f; // @[Switch.scala 30:53:@10133.4]
  assign valid_31_47 = io_inValid_47 & _T_29730; // @[Switch.scala 30:36:@10134.4]
  assign _T_29733 = io_inAddr_48 == 6'h1f; // @[Switch.scala 30:53:@10136.4]
  assign valid_31_48 = io_inValid_48 & _T_29733; // @[Switch.scala 30:36:@10137.4]
  assign _T_29736 = io_inAddr_49 == 6'h1f; // @[Switch.scala 30:53:@10139.4]
  assign valid_31_49 = io_inValid_49 & _T_29736; // @[Switch.scala 30:36:@10140.4]
  assign _T_29739 = io_inAddr_50 == 6'h1f; // @[Switch.scala 30:53:@10142.4]
  assign valid_31_50 = io_inValid_50 & _T_29739; // @[Switch.scala 30:36:@10143.4]
  assign _T_29742 = io_inAddr_51 == 6'h1f; // @[Switch.scala 30:53:@10145.4]
  assign valid_31_51 = io_inValid_51 & _T_29742; // @[Switch.scala 30:36:@10146.4]
  assign _T_29745 = io_inAddr_52 == 6'h1f; // @[Switch.scala 30:53:@10148.4]
  assign valid_31_52 = io_inValid_52 & _T_29745; // @[Switch.scala 30:36:@10149.4]
  assign _T_29748 = io_inAddr_53 == 6'h1f; // @[Switch.scala 30:53:@10151.4]
  assign valid_31_53 = io_inValid_53 & _T_29748; // @[Switch.scala 30:36:@10152.4]
  assign _T_29751 = io_inAddr_54 == 6'h1f; // @[Switch.scala 30:53:@10154.4]
  assign valid_31_54 = io_inValid_54 & _T_29751; // @[Switch.scala 30:36:@10155.4]
  assign _T_29754 = io_inAddr_55 == 6'h1f; // @[Switch.scala 30:53:@10157.4]
  assign valid_31_55 = io_inValid_55 & _T_29754; // @[Switch.scala 30:36:@10158.4]
  assign _T_29757 = io_inAddr_56 == 6'h1f; // @[Switch.scala 30:53:@10160.4]
  assign valid_31_56 = io_inValid_56 & _T_29757; // @[Switch.scala 30:36:@10161.4]
  assign _T_29760 = io_inAddr_57 == 6'h1f; // @[Switch.scala 30:53:@10163.4]
  assign valid_31_57 = io_inValid_57 & _T_29760; // @[Switch.scala 30:36:@10164.4]
  assign _T_29763 = io_inAddr_58 == 6'h1f; // @[Switch.scala 30:53:@10166.4]
  assign valid_31_58 = io_inValid_58 & _T_29763; // @[Switch.scala 30:36:@10167.4]
  assign _T_29766 = io_inAddr_59 == 6'h1f; // @[Switch.scala 30:53:@10169.4]
  assign valid_31_59 = io_inValid_59 & _T_29766; // @[Switch.scala 30:36:@10170.4]
  assign _T_29769 = io_inAddr_60 == 6'h1f; // @[Switch.scala 30:53:@10172.4]
  assign valid_31_60 = io_inValid_60 & _T_29769; // @[Switch.scala 30:36:@10173.4]
  assign _T_29772 = io_inAddr_61 == 6'h1f; // @[Switch.scala 30:53:@10175.4]
  assign valid_31_61 = io_inValid_61 & _T_29772; // @[Switch.scala 30:36:@10176.4]
  assign _T_29775 = io_inAddr_62 == 6'h1f; // @[Switch.scala 30:53:@10178.4]
  assign valid_31_62 = io_inValid_62 & _T_29775; // @[Switch.scala 30:36:@10179.4]
  assign _T_29778 = io_inAddr_63 == 6'h1f; // @[Switch.scala 30:53:@10181.4]
  assign valid_31_63 = io_inValid_63 & _T_29778; // @[Switch.scala 30:36:@10182.4]
  assign _T_29844 = valid_31_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@10184.4]
  assign _T_29845 = valid_31_61 ? 6'h3d : _T_29844; // @[Mux.scala 31:69:@10185.4]
  assign _T_29846 = valid_31_60 ? 6'h3c : _T_29845; // @[Mux.scala 31:69:@10186.4]
  assign _T_29847 = valid_31_59 ? 6'h3b : _T_29846; // @[Mux.scala 31:69:@10187.4]
  assign _T_29848 = valid_31_58 ? 6'h3a : _T_29847; // @[Mux.scala 31:69:@10188.4]
  assign _T_29849 = valid_31_57 ? 6'h39 : _T_29848; // @[Mux.scala 31:69:@10189.4]
  assign _T_29850 = valid_31_56 ? 6'h38 : _T_29849; // @[Mux.scala 31:69:@10190.4]
  assign _T_29851 = valid_31_55 ? 6'h37 : _T_29850; // @[Mux.scala 31:69:@10191.4]
  assign _T_29852 = valid_31_54 ? 6'h36 : _T_29851; // @[Mux.scala 31:69:@10192.4]
  assign _T_29853 = valid_31_53 ? 6'h35 : _T_29852; // @[Mux.scala 31:69:@10193.4]
  assign _T_29854 = valid_31_52 ? 6'h34 : _T_29853; // @[Mux.scala 31:69:@10194.4]
  assign _T_29855 = valid_31_51 ? 6'h33 : _T_29854; // @[Mux.scala 31:69:@10195.4]
  assign _T_29856 = valid_31_50 ? 6'h32 : _T_29855; // @[Mux.scala 31:69:@10196.4]
  assign _T_29857 = valid_31_49 ? 6'h31 : _T_29856; // @[Mux.scala 31:69:@10197.4]
  assign _T_29858 = valid_31_48 ? 6'h30 : _T_29857; // @[Mux.scala 31:69:@10198.4]
  assign _T_29859 = valid_31_47 ? 6'h2f : _T_29858; // @[Mux.scala 31:69:@10199.4]
  assign _T_29860 = valid_31_46 ? 6'h2e : _T_29859; // @[Mux.scala 31:69:@10200.4]
  assign _T_29861 = valid_31_45 ? 6'h2d : _T_29860; // @[Mux.scala 31:69:@10201.4]
  assign _T_29862 = valid_31_44 ? 6'h2c : _T_29861; // @[Mux.scala 31:69:@10202.4]
  assign _T_29863 = valid_31_43 ? 6'h2b : _T_29862; // @[Mux.scala 31:69:@10203.4]
  assign _T_29864 = valid_31_42 ? 6'h2a : _T_29863; // @[Mux.scala 31:69:@10204.4]
  assign _T_29865 = valid_31_41 ? 6'h29 : _T_29864; // @[Mux.scala 31:69:@10205.4]
  assign _T_29866 = valid_31_40 ? 6'h28 : _T_29865; // @[Mux.scala 31:69:@10206.4]
  assign _T_29867 = valid_31_39 ? 6'h27 : _T_29866; // @[Mux.scala 31:69:@10207.4]
  assign _T_29868 = valid_31_38 ? 6'h26 : _T_29867; // @[Mux.scala 31:69:@10208.4]
  assign _T_29869 = valid_31_37 ? 6'h25 : _T_29868; // @[Mux.scala 31:69:@10209.4]
  assign _T_29870 = valid_31_36 ? 6'h24 : _T_29869; // @[Mux.scala 31:69:@10210.4]
  assign _T_29871 = valid_31_35 ? 6'h23 : _T_29870; // @[Mux.scala 31:69:@10211.4]
  assign _T_29872 = valid_31_34 ? 6'h22 : _T_29871; // @[Mux.scala 31:69:@10212.4]
  assign _T_29873 = valid_31_33 ? 6'h21 : _T_29872; // @[Mux.scala 31:69:@10213.4]
  assign _T_29874 = valid_31_32 ? 6'h20 : _T_29873; // @[Mux.scala 31:69:@10214.4]
  assign _T_29875 = valid_31_31 ? 6'h1f : _T_29874; // @[Mux.scala 31:69:@10215.4]
  assign _T_29876 = valid_31_30 ? 6'h1e : _T_29875; // @[Mux.scala 31:69:@10216.4]
  assign _T_29877 = valid_31_29 ? 6'h1d : _T_29876; // @[Mux.scala 31:69:@10217.4]
  assign _T_29878 = valid_31_28 ? 6'h1c : _T_29877; // @[Mux.scala 31:69:@10218.4]
  assign _T_29879 = valid_31_27 ? 6'h1b : _T_29878; // @[Mux.scala 31:69:@10219.4]
  assign _T_29880 = valid_31_26 ? 6'h1a : _T_29879; // @[Mux.scala 31:69:@10220.4]
  assign _T_29881 = valid_31_25 ? 6'h19 : _T_29880; // @[Mux.scala 31:69:@10221.4]
  assign _T_29882 = valid_31_24 ? 6'h18 : _T_29881; // @[Mux.scala 31:69:@10222.4]
  assign _T_29883 = valid_31_23 ? 6'h17 : _T_29882; // @[Mux.scala 31:69:@10223.4]
  assign _T_29884 = valid_31_22 ? 6'h16 : _T_29883; // @[Mux.scala 31:69:@10224.4]
  assign _T_29885 = valid_31_21 ? 6'h15 : _T_29884; // @[Mux.scala 31:69:@10225.4]
  assign _T_29886 = valid_31_20 ? 6'h14 : _T_29885; // @[Mux.scala 31:69:@10226.4]
  assign _T_29887 = valid_31_19 ? 6'h13 : _T_29886; // @[Mux.scala 31:69:@10227.4]
  assign _T_29888 = valid_31_18 ? 6'h12 : _T_29887; // @[Mux.scala 31:69:@10228.4]
  assign _T_29889 = valid_31_17 ? 6'h11 : _T_29888; // @[Mux.scala 31:69:@10229.4]
  assign _T_29890 = valid_31_16 ? 6'h10 : _T_29889; // @[Mux.scala 31:69:@10230.4]
  assign _T_29891 = valid_31_15 ? 6'hf : _T_29890; // @[Mux.scala 31:69:@10231.4]
  assign _T_29892 = valid_31_14 ? 6'he : _T_29891; // @[Mux.scala 31:69:@10232.4]
  assign _T_29893 = valid_31_13 ? 6'hd : _T_29892; // @[Mux.scala 31:69:@10233.4]
  assign _T_29894 = valid_31_12 ? 6'hc : _T_29893; // @[Mux.scala 31:69:@10234.4]
  assign _T_29895 = valid_31_11 ? 6'hb : _T_29894; // @[Mux.scala 31:69:@10235.4]
  assign _T_29896 = valid_31_10 ? 6'ha : _T_29895; // @[Mux.scala 31:69:@10236.4]
  assign _T_29897 = valid_31_9 ? 6'h9 : _T_29896; // @[Mux.scala 31:69:@10237.4]
  assign _T_29898 = valid_31_8 ? 6'h8 : _T_29897; // @[Mux.scala 31:69:@10238.4]
  assign _T_29899 = valid_31_7 ? 6'h7 : _T_29898; // @[Mux.scala 31:69:@10239.4]
  assign _T_29900 = valid_31_6 ? 6'h6 : _T_29899; // @[Mux.scala 31:69:@10240.4]
  assign _T_29901 = valid_31_5 ? 6'h5 : _T_29900; // @[Mux.scala 31:69:@10241.4]
  assign _T_29902 = valid_31_4 ? 6'h4 : _T_29901; // @[Mux.scala 31:69:@10242.4]
  assign _T_29903 = valid_31_3 ? 6'h3 : _T_29902; // @[Mux.scala 31:69:@10243.4]
  assign _T_29904 = valid_31_2 ? 6'h2 : _T_29903; // @[Mux.scala 31:69:@10244.4]
  assign _T_29905 = valid_31_1 ? 6'h1 : _T_29904; // @[Mux.scala 31:69:@10245.4]
  assign select_31 = valid_31_0 ? 6'h0 : _T_29905; // @[Mux.scala 31:69:@10246.4]
  assign _GEN_1985 = 6'h1 == select_31 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_1986 = 6'h2 == select_31 ? io_inData_2 : _GEN_1985; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_1987 = 6'h3 == select_31 ? io_inData_3 : _GEN_1986; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_1988 = 6'h4 == select_31 ? io_inData_4 : _GEN_1987; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_1989 = 6'h5 == select_31 ? io_inData_5 : _GEN_1988; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_1990 = 6'h6 == select_31 ? io_inData_6 : _GEN_1989; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_1991 = 6'h7 == select_31 ? io_inData_7 : _GEN_1990; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_1992 = 6'h8 == select_31 ? io_inData_8 : _GEN_1991; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_1993 = 6'h9 == select_31 ? io_inData_9 : _GEN_1992; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_1994 = 6'ha == select_31 ? io_inData_10 : _GEN_1993; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_1995 = 6'hb == select_31 ? io_inData_11 : _GEN_1994; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_1996 = 6'hc == select_31 ? io_inData_12 : _GEN_1995; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_1997 = 6'hd == select_31 ? io_inData_13 : _GEN_1996; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_1998 = 6'he == select_31 ? io_inData_14 : _GEN_1997; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_1999 = 6'hf == select_31 ? io_inData_15 : _GEN_1998; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2000 = 6'h10 == select_31 ? io_inData_16 : _GEN_1999; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2001 = 6'h11 == select_31 ? io_inData_17 : _GEN_2000; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2002 = 6'h12 == select_31 ? io_inData_18 : _GEN_2001; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2003 = 6'h13 == select_31 ? io_inData_19 : _GEN_2002; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2004 = 6'h14 == select_31 ? io_inData_20 : _GEN_2003; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2005 = 6'h15 == select_31 ? io_inData_21 : _GEN_2004; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2006 = 6'h16 == select_31 ? io_inData_22 : _GEN_2005; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2007 = 6'h17 == select_31 ? io_inData_23 : _GEN_2006; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2008 = 6'h18 == select_31 ? io_inData_24 : _GEN_2007; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2009 = 6'h19 == select_31 ? io_inData_25 : _GEN_2008; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2010 = 6'h1a == select_31 ? io_inData_26 : _GEN_2009; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2011 = 6'h1b == select_31 ? io_inData_27 : _GEN_2010; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2012 = 6'h1c == select_31 ? io_inData_28 : _GEN_2011; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2013 = 6'h1d == select_31 ? io_inData_29 : _GEN_2012; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2014 = 6'h1e == select_31 ? io_inData_30 : _GEN_2013; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2015 = 6'h1f == select_31 ? io_inData_31 : _GEN_2014; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2016 = 6'h20 == select_31 ? io_inData_32 : _GEN_2015; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2017 = 6'h21 == select_31 ? io_inData_33 : _GEN_2016; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2018 = 6'h22 == select_31 ? io_inData_34 : _GEN_2017; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2019 = 6'h23 == select_31 ? io_inData_35 : _GEN_2018; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2020 = 6'h24 == select_31 ? io_inData_36 : _GEN_2019; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2021 = 6'h25 == select_31 ? io_inData_37 : _GEN_2020; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2022 = 6'h26 == select_31 ? io_inData_38 : _GEN_2021; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2023 = 6'h27 == select_31 ? io_inData_39 : _GEN_2022; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2024 = 6'h28 == select_31 ? io_inData_40 : _GEN_2023; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2025 = 6'h29 == select_31 ? io_inData_41 : _GEN_2024; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2026 = 6'h2a == select_31 ? io_inData_42 : _GEN_2025; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2027 = 6'h2b == select_31 ? io_inData_43 : _GEN_2026; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2028 = 6'h2c == select_31 ? io_inData_44 : _GEN_2027; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2029 = 6'h2d == select_31 ? io_inData_45 : _GEN_2028; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2030 = 6'h2e == select_31 ? io_inData_46 : _GEN_2029; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2031 = 6'h2f == select_31 ? io_inData_47 : _GEN_2030; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2032 = 6'h30 == select_31 ? io_inData_48 : _GEN_2031; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2033 = 6'h31 == select_31 ? io_inData_49 : _GEN_2032; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2034 = 6'h32 == select_31 ? io_inData_50 : _GEN_2033; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2035 = 6'h33 == select_31 ? io_inData_51 : _GEN_2034; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2036 = 6'h34 == select_31 ? io_inData_52 : _GEN_2035; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2037 = 6'h35 == select_31 ? io_inData_53 : _GEN_2036; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2038 = 6'h36 == select_31 ? io_inData_54 : _GEN_2037; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2039 = 6'h37 == select_31 ? io_inData_55 : _GEN_2038; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2040 = 6'h38 == select_31 ? io_inData_56 : _GEN_2039; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2041 = 6'h39 == select_31 ? io_inData_57 : _GEN_2040; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2042 = 6'h3a == select_31 ? io_inData_58 : _GEN_2041; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2043 = 6'h3b == select_31 ? io_inData_59 : _GEN_2042; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2044 = 6'h3c == select_31 ? io_inData_60 : _GEN_2043; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2045 = 6'h3d == select_31 ? io_inData_61 : _GEN_2044; // @[Switch.scala 33:19:@10248.4]
  assign _GEN_2046 = 6'h3e == select_31 ? io_inData_62 : _GEN_2045; // @[Switch.scala 33:19:@10248.4]
  assign _T_29914 = {valid_31_7,valid_31_6,valid_31_5,valid_31_4,valid_31_3,valid_31_2,valid_31_1,valid_31_0}; // @[Switch.scala 34:32:@10255.4]
  assign _T_29922 = {valid_31_15,valid_31_14,valid_31_13,valid_31_12,valid_31_11,valid_31_10,valid_31_9,valid_31_8,_T_29914}; // @[Switch.scala 34:32:@10263.4]
  assign _T_29929 = {valid_31_23,valid_31_22,valid_31_21,valid_31_20,valid_31_19,valid_31_18,valid_31_17,valid_31_16}; // @[Switch.scala 34:32:@10270.4]
  assign _T_29938 = {valid_31_31,valid_31_30,valid_31_29,valid_31_28,valid_31_27,valid_31_26,valid_31_25,valid_31_24,_T_29929,_T_29922}; // @[Switch.scala 34:32:@10279.4]
  assign _T_29945 = {valid_31_39,valid_31_38,valid_31_37,valid_31_36,valid_31_35,valid_31_34,valid_31_33,valid_31_32}; // @[Switch.scala 34:32:@10286.4]
  assign _T_29953 = {valid_31_47,valid_31_46,valid_31_45,valid_31_44,valid_31_43,valid_31_42,valid_31_41,valid_31_40,_T_29945}; // @[Switch.scala 34:32:@10294.4]
  assign _T_29960 = {valid_31_55,valid_31_54,valid_31_53,valid_31_52,valid_31_51,valid_31_50,valid_31_49,valid_31_48}; // @[Switch.scala 34:32:@10301.4]
  assign _T_29969 = {valid_31_63,valid_31_62,valid_31_61,valid_31_60,valid_31_59,valid_31_58,valid_31_57,valid_31_56,_T_29960,_T_29953}; // @[Switch.scala 34:32:@10310.4]
  assign _T_29970 = {_T_29969,_T_29938}; // @[Switch.scala 34:32:@10311.4]
  assign _T_29974 = io_inAddr_0 == 6'h20; // @[Switch.scala 30:53:@10314.4]
  assign valid_32_0 = io_inValid_0 & _T_29974; // @[Switch.scala 30:36:@10315.4]
  assign _T_29977 = io_inAddr_1 == 6'h20; // @[Switch.scala 30:53:@10317.4]
  assign valid_32_1 = io_inValid_1 & _T_29977; // @[Switch.scala 30:36:@10318.4]
  assign _T_29980 = io_inAddr_2 == 6'h20; // @[Switch.scala 30:53:@10320.4]
  assign valid_32_2 = io_inValid_2 & _T_29980; // @[Switch.scala 30:36:@10321.4]
  assign _T_29983 = io_inAddr_3 == 6'h20; // @[Switch.scala 30:53:@10323.4]
  assign valid_32_3 = io_inValid_3 & _T_29983; // @[Switch.scala 30:36:@10324.4]
  assign _T_29986 = io_inAddr_4 == 6'h20; // @[Switch.scala 30:53:@10326.4]
  assign valid_32_4 = io_inValid_4 & _T_29986; // @[Switch.scala 30:36:@10327.4]
  assign _T_29989 = io_inAddr_5 == 6'h20; // @[Switch.scala 30:53:@10329.4]
  assign valid_32_5 = io_inValid_5 & _T_29989; // @[Switch.scala 30:36:@10330.4]
  assign _T_29992 = io_inAddr_6 == 6'h20; // @[Switch.scala 30:53:@10332.4]
  assign valid_32_6 = io_inValid_6 & _T_29992; // @[Switch.scala 30:36:@10333.4]
  assign _T_29995 = io_inAddr_7 == 6'h20; // @[Switch.scala 30:53:@10335.4]
  assign valid_32_7 = io_inValid_7 & _T_29995; // @[Switch.scala 30:36:@10336.4]
  assign _T_29998 = io_inAddr_8 == 6'h20; // @[Switch.scala 30:53:@10338.4]
  assign valid_32_8 = io_inValid_8 & _T_29998; // @[Switch.scala 30:36:@10339.4]
  assign _T_30001 = io_inAddr_9 == 6'h20; // @[Switch.scala 30:53:@10341.4]
  assign valid_32_9 = io_inValid_9 & _T_30001; // @[Switch.scala 30:36:@10342.4]
  assign _T_30004 = io_inAddr_10 == 6'h20; // @[Switch.scala 30:53:@10344.4]
  assign valid_32_10 = io_inValid_10 & _T_30004; // @[Switch.scala 30:36:@10345.4]
  assign _T_30007 = io_inAddr_11 == 6'h20; // @[Switch.scala 30:53:@10347.4]
  assign valid_32_11 = io_inValid_11 & _T_30007; // @[Switch.scala 30:36:@10348.4]
  assign _T_30010 = io_inAddr_12 == 6'h20; // @[Switch.scala 30:53:@10350.4]
  assign valid_32_12 = io_inValid_12 & _T_30010; // @[Switch.scala 30:36:@10351.4]
  assign _T_30013 = io_inAddr_13 == 6'h20; // @[Switch.scala 30:53:@10353.4]
  assign valid_32_13 = io_inValid_13 & _T_30013; // @[Switch.scala 30:36:@10354.4]
  assign _T_30016 = io_inAddr_14 == 6'h20; // @[Switch.scala 30:53:@10356.4]
  assign valid_32_14 = io_inValid_14 & _T_30016; // @[Switch.scala 30:36:@10357.4]
  assign _T_30019 = io_inAddr_15 == 6'h20; // @[Switch.scala 30:53:@10359.4]
  assign valid_32_15 = io_inValid_15 & _T_30019; // @[Switch.scala 30:36:@10360.4]
  assign _T_30022 = io_inAddr_16 == 6'h20; // @[Switch.scala 30:53:@10362.4]
  assign valid_32_16 = io_inValid_16 & _T_30022; // @[Switch.scala 30:36:@10363.4]
  assign _T_30025 = io_inAddr_17 == 6'h20; // @[Switch.scala 30:53:@10365.4]
  assign valid_32_17 = io_inValid_17 & _T_30025; // @[Switch.scala 30:36:@10366.4]
  assign _T_30028 = io_inAddr_18 == 6'h20; // @[Switch.scala 30:53:@10368.4]
  assign valid_32_18 = io_inValid_18 & _T_30028; // @[Switch.scala 30:36:@10369.4]
  assign _T_30031 = io_inAddr_19 == 6'h20; // @[Switch.scala 30:53:@10371.4]
  assign valid_32_19 = io_inValid_19 & _T_30031; // @[Switch.scala 30:36:@10372.4]
  assign _T_30034 = io_inAddr_20 == 6'h20; // @[Switch.scala 30:53:@10374.4]
  assign valid_32_20 = io_inValid_20 & _T_30034; // @[Switch.scala 30:36:@10375.4]
  assign _T_30037 = io_inAddr_21 == 6'h20; // @[Switch.scala 30:53:@10377.4]
  assign valid_32_21 = io_inValid_21 & _T_30037; // @[Switch.scala 30:36:@10378.4]
  assign _T_30040 = io_inAddr_22 == 6'h20; // @[Switch.scala 30:53:@10380.4]
  assign valid_32_22 = io_inValid_22 & _T_30040; // @[Switch.scala 30:36:@10381.4]
  assign _T_30043 = io_inAddr_23 == 6'h20; // @[Switch.scala 30:53:@10383.4]
  assign valid_32_23 = io_inValid_23 & _T_30043; // @[Switch.scala 30:36:@10384.4]
  assign _T_30046 = io_inAddr_24 == 6'h20; // @[Switch.scala 30:53:@10386.4]
  assign valid_32_24 = io_inValid_24 & _T_30046; // @[Switch.scala 30:36:@10387.4]
  assign _T_30049 = io_inAddr_25 == 6'h20; // @[Switch.scala 30:53:@10389.4]
  assign valid_32_25 = io_inValid_25 & _T_30049; // @[Switch.scala 30:36:@10390.4]
  assign _T_30052 = io_inAddr_26 == 6'h20; // @[Switch.scala 30:53:@10392.4]
  assign valid_32_26 = io_inValid_26 & _T_30052; // @[Switch.scala 30:36:@10393.4]
  assign _T_30055 = io_inAddr_27 == 6'h20; // @[Switch.scala 30:53:@10395.4]
  assign valid_32_27 = io_inValid_27 & _T_30055; // @[Switch.scala 30:36:@10396.4]
  assign _T_30058 = io_inAddr_28 == 6'h20; // @[Switch.scala 30:53:@10398.4]
  assign valid_32_28 = io_inValid_28 & _T_30058; // @[Switch.scala 30:36:@10399.4]
  assign _T_30061 = io_inAddr_29 == 6'h20; // @[Switch.scala 30:53:@10401.4]
  assign valid_32_29 = io_inValid_29 & _T_30061; // @[Switch.scala 30:36:@10402.4]
  assign _T_30064 = io_inAddr_30 == 6'h20; // @[Switch.scala 30:53:@10404.4]
  assign valid_32_30 = io_inValid_30 & _T_30064; // @[Switch.scala 30:36:@10405.4]
  assign _T_30067 = io_inAddr_31 == 6'h20; // @[Switch.scala 30:53:@10407.4]
  assign valid_32_31 = io_inValid_31 & _T_30067; // @[Switch.scala 30:36:@10408.4]
  assign _T_30070 = io_inAddr_32 == 6'h20; // @[Switch.scala 30:53:@10410.4]
  assign valid_32_32 = io_inValid_32 & _T_30070; // @[Switch.scala 30:36:@10411.4]
  assign _T_30073 = io_inAddr_33 == 6'h20; // @[Switch.scala 30:53:@10413.4]
  assign valid_32_33 = io_inValid_33 & _T_30073; // @[Switch.scala 30:36:@10414.4]
  assign _T_30076 = io_inAddr_34 == 6'h20; // @[Switch.scala 30:53:@10416.4]
  assign valid_32_34 = io_inValid_34 & _T_30076; // @[Switch.scala 30:36:@10417.4]
  assign _T_30079 = io_inAddr_35 == 6'h20; // @[Switch.scala 30:53:@10419.4]
  assign valid_32_35 = io_inValid_35 & _T_30079; // @[Switch.scala 30:36:@10420.4]
  assign _T_30082 = io_inAddr_36 == 6'h20; // @[Switch.scala 30:53:@10422.4]
  assign valid_32_36 = io_inValid_36 & _T_30082; // @[Switch.scala 30:36:@10423.4]
  assign _T_30085 = io_inAddr_37 == 6'h20; // @[Switch.scala 30:53:@10425.4]
  assign valid_32_37 = io_inValid_37 & _T_30085; // @[Switch.scala 30:36:@10426.4]
  assign _T_30088 = io_inAddr_38 == 6'h20; // @[Switch.scala 30:53:@10428.4]
  assign valid_32_38 = io_inValid_38 & _T_30088; // @[Switch.scala 30:36:@10429.4]
  assign _T_30091 = io_inAddr_39 == 6'h20; // @[Switch.scala 30:53:@10431.4]
  assign valid_32_39 = io_inValid_39 & _T_30091; // @[Switch.scala 30:36:@10432.4]
  assign _T_30094 = io_inAddr_40 == 6'h20; // @[Switch.scala 30:53:@10434.4]
  assign valid_32_40 = io_inValid_40 & _T_30094; // @[Switch.scala 30:36:@10435.4]
  assign _T_30097 = io_inAddr_41 == 6'h20; // @[Switch.scala 30:53:@10437.4]
  assign valid_32_41 = io_inValid_41 & _T_30097; // @[Switch.scala 30:36:@10438.4]
  assign _T_30100 = io_inAddr_42 == 6'h20; // @[Switch.scala 30:53:@10440.4]
  assign valid_32_42 = io_inValid_42 & _T_30100; // @[Switch.scala 30:36:@10441.4]
  assign _T_30103 = io_inAddr_43 == 6'h20; // @[Switch.scala 30:53:@10443.4]
  assign valid_32_43 = io_inValid_43 & _T_30103; // @[Switch.scala 30:36:@10444.4]
  assign _T_30106 = io_inAddr_44 == 6'h20; // @[Switch.scala 30:53:@10446.4]
  assign valid_32_44 = io_inValid_44 & _T_30106; // @[Switch.scala 30:36:@10447.4]
  assign _T_30109 = io_inAddr_45 == 6'h20; // @[Switch.scala 30:53:@10449.4]
  assign valid_32_45 = io_inValid_45 & _T_30109; // @[Switch.scala 30:36:@10450.4]
  assign _T_30112 = io_inAddr_46 == 6'h20; // @[Switch.scala 30:53:@10452.4]
  assign valid_32_46 = io_inValid_46 & _T_30112; // @[Switch.scala 30:36:@10453.4]
  assign _T_30115 = io_inAddr_47 == 6'h20; // @[Switch.scala 30:53:@10455.4]
  assign valid_32_47 = io_inValid_47 & _T_30115; // @[Switch.scala 30:36:@10456.4]
  assign _T_30118 = io_inAddr_48 == 6'h20; // @[Switch.scala 30:53:@10458.4]
  assign valid_32_48 = io_inValid_48 & _T_30118; // @[Switch.scala 30:36:@10459.4]
  assign _T_30121 = io_inAddr_49 == 6'h20; // @[Switch.scala 30:53:@10461.4]
  assign valid_32_49 = io_inValid_49 & _T_30121; // @[Switch.scala 30:36:@10462.4]
  assign _T_30124 = io_inAddr_50 == 6'h20; // @[Switch.scala 30:53:@10464.4]
  assign valid_32_50 = io_inValid_50 & _T_30124; // @[Switch.scala 30:36:@10465.4]
  assign _T_30127 = io_inAddr_51 == 6'h20; // @[Switch.scala 30:53:@10467.4]
  assign valid_32_51 = io_inValid_51 & _T_30127; // @[Switch.scala 30:36:@10468.4]
  assign _T_30130 = io_inAddr_52 == 6'h20; // @[Switch.scala 30:53:@10470.4]
  assign valid_32_52 = io_inValid_52 & _T_30130; // @[Switch.scala 30:36:@10471.4]
  assign _T_30133 = io_inAddr_53 == 6'h20; // @[Switch.scala 30:53:@10473.4]
  assign valid_32_53 = io_inValid_53 & _T_30133; // @[Switch.scala 30:36:@10474.4]
  assign _T_30136 = io_inAddr_54 == 6'h20; // @[Switch.scala 30:53:@10476.4]
  assign valid_32_54 = io_inValid_54 & _T_30136; // @[Switch.scala 30:36:@10477.4]
  assign _T_30139 = io_inAddr_55 == 6'h20; // @[Switch.scala 30:53:@10479.4]
  assign valid_32_55 = io_inValid_55 & _T_30139; // @[Switch.scala 30:36:@10480.4]
  assign _T_30142 = io_inAddr_56 == 6'h20; // @[Switch.scala 30:53:@10482.4]
  assign valid_32_56 = io_inValid_56 & _T_30142; // @[Switch.scala 30:36:@10483.4]
  assign _T_30145 = io_inAddr_57 == 6'h20; // @[Switch.scala 30:53:@10485.4]
  assign valid_32_57 = io_inValid_57 & _T_30145; // @[Switch.scala 30:36:@10486.4]
  assign _T_30148 = io_inAddr_58 == 6'h20; // @[Switch.scala 30:53:@10488.4]
  assign valid_32_58 = io_inValid_58 & _T_30148; // @[Switch.scala 30:36:@10489.4]
  assign _T_30151 = io_inAddr_59 == 6'h20; // @[Switch.scala 30:53:@10491.4]
  assign valid_32_59 = io_inValid_59 & _T_30151; // @[Switch.scala 30:36:@10492.4]
  assign _T_30154 = io_inAddr_60 == 6'h20; // @[Switch.scala 30:53:@10494.4]
  assign valid_32_60 = io_inValid_60 & _T_30154; // @[Switch.scala 30:36:@10495.4]
  assign _T_30157 = io_inAddr_61 == 6'h20; // @[Switch.scala 30:53:@10497.4]
  assign valid_32_61 = io_inValid_61 & _T_30157; // @[Switch.scala 30:36:@10498.4]
  assign _T_30160 = io_inAddr_62 == 6'h20; // @[Switch.scala 30:53:@10500.4]
  assign valid_32_62 = io_inValid_62 & _T_30160; // @[Switch.scala 30:36:@10501.4]
  assign _T_30163 = io_inAddr_63 == 6'h20; // @[Switch.scala 30:53:@10503.4]
  assign valid_32_63 = io_inValid_63 & _T_30163; // @[Switch.scala 30:36:@10504.4]
  assign _T_30229 = valid_32_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@10506.4]
  assign _T_30230 = valid_32_61 ? 6'h3d : _T_30229; // @[Mux.scala 31:69:@10507.4]
  assign _T_30231 = valid_32_60 ? 6'h3c : _T_30230; // @[Mux.scala 31:69:@10508.4]
  assign _T_30232 = valid_32_59 ? 6'h3b : _T_30231; // @[Mux.scala 31:69:@10509.4]
  assign _T_30233 = valid_32_58 ? 6'h3a : _T_30232; // @[Mux.scala 31:69:@10510.4]
  assign _T_30234 = valid_32_57 ? 6'h39 : _T_30233; // @[Mux.scala 31:69:@10511.4]
  assign _T_30235 = valid_32_56 ? 6'h38 : _T_30234; // @[Mux.scala 31:69:@10512.4]
  assign _T_30236 = valid_32_55 ? 6'h37 : _T_30235; // @[Mux.scala 31:69:@10513.4]
  assign _T_30237 = valid_32_54 ? 6'h36 : _T_30236; // @[Mux.scala 31:69:@10514.4]
  assign _T_30238 = valid_32_53 ? 6'h35 : _T_30237; // @[Mux.scala 31:69:@10515.4]
  assign _T_30239 = valid_32_52 ? 6'h34 : _T_30238; // @[Mux.scala 31:69:@10516.4]
  assign _T_30240 = valid_32_51 ? 6'h33 : _T_30239; // @[Mux.scala 31:69:@10517.4]
  assign _T_30241 = valid_32_50 ? 6'h32 : _T_30240; // @[Mux.scala 31:69:@10518.4]
  assign _T_30242 = valid_32_49 ? 6'h31 : _T_30241; // @[Mux.scala 31:69:@10519.4]
  assign _T_30243 = valid_32_48 ? 6'h30 : _T_30242; // @[Mux.scala 31:69:@10520.4]
  assign _T_30244 = valid_32_47 ? 6'h2f : _T_30243; // @[Mux.scala 31:69:@10521.4]
  assign _T_30245 = valid_32_46 ? 6'h2e : _T_30244; // @[Mux.scala 31:69:@10522.4]
  assign _T_30246 = valid_32_45 ? 6'h2d : _T_30245; // @[Mux.scala 31:69:@10523.4]
  assign _T_30247 = valid_32_44 ? 6'h2c : _T_30246; // @[Mux.scala 31:69:@10524.4]
  assign _T_30248 = valid_32_43 ? 6'h2b : _T_30247; // @[Mux.scala 31:69:@10525.4]
  assign _T_30249 = valid_32_42 ? 6'h2a : _T_30248; // @[Mux.scala 31:69:@10526.4]
  assign _T_30250 = valid_32_41 ? 6'h29 : _T_30249; // @[Mux.scala 31:69:@10527.4]
  assign _T_30251 = valid_32_40 ? 6'h28 : _T_30250; // @[Mux.scala 31:69:@10528.4]
  assign _T_30252 = valid_32_39 ? 6'h27 : _T_30251; // @[Mux.scala 31:69:@10529.4]
  assign _T_30253 = valid_32_38 ? 6'h26 : _T_30252; // @[Mux.scala 31:69:@10530.4]
  assign _T_30254 = valid_32_37 ? 6'h25 : _T_30253; // @[Mux.scala 31:69:@10531.4]
  assign _T_30255 = valid_32_36 ? 6'h24 : _T_30254; // @[Mux.scala 31:69:@10532.4]
  assign _T_30256 = valid_32_35 ? 6'h23 : _T_30255; // @[Mux.scala 31:69:@10533.4]
  assign _T_30257 = valid_32_34 ? 6'h22 : _T_30256; // @[Mux.scala 31:69:@10534.4]
  assign _T_30258 = valid_32_33 ? 6'h21 : _T_30257; // @[Mux.scala 31:69:@10535.4]
  assign _T_30259 = valid_32_32 ? 6'h20 : _T_30258; // @[Mux.scala 31:69:@10536.4]
  assign _T_30260 = valid_32_31 ? 6'h1f : _T_30259; // @[Mux.scala 31:69:@10537.4]
  assign _T_30261 = valid_32_30 ? 6'h1e : _T_30260; // @[Mux.scala 31:69:@10538.4]
  assign _T_30262 = valid_32_29 ? 6'h1d : _T_30261; // @[Mux.scala 31:69:@10539.4]
  assign _T_30263 = valid_32_28 ? 6'h1c : _T_30262; // @[Mux.scala 31:69:@10540.4]
  assign _T_30264 = valid_32_27 ? 6'h1b : _T_30263; // @[Mux.scala 31:69:@10541.4]
  assign _T_30265 = valid_32_26 ? 6'h1a : _T_30264; // @[Mux.scala 31:69:@10542.4]
  assign _T_30266 = valid_32_25 ? 6'h19 : _T_30265; // @[Mux.scala 31:69:@10543.4]
  assign _T_30267 = valid_32_24 ? 6'h18 : _T_30266; // @[Mux.scala 31:69:@10544.4]
  assign _T_30268 = valid_32_23 ? 6'h17 : _T_30267; // @[Mux.scala 31:69:@10545.4]
  assign _T_30269 = valid_32_22 ? 6'h16 : _T_30268; // @[Mux.scala 31:69:@10546.4]
  assign _T_30270 = valid_32_21 ? 6'h15 : _T_30269; // @[Mux.scala 31:69:@10547.4]
  assign _T_30271 = valid_32_20 ? 6'h14 : _T_30270; // @[Mux.scala 31:69:@10548.4]
  assign _T_30272 = valid_32_19 ? 6'h13 : _T_30271; // @[Mux.scala 31:69:@10549.4]
  assign _T_30273 = valid_32_18 ? 6'h12 : _T_30272; // @[Mux.scala 31:69:@10550.4]
  assign _T_30274 = valid_32_17 ? 6'h11 : _T_30273; // @[Mux.scala 31:69:@10551.4]
  assign _T_30275 = valid_32_16 ? 6'h10 : _T_30274; // @[Mux.scala 31:69:@10552.4]
  assign _T_30276 = valid_32_15 ? 6'hf : _T_30275; // @[Mux.scala 31:69:@10553.4]
  assign _T_30277 = valid_32_14 ? 6'he : _T_30276; // @[Mux.scala 31:69:@10554.4]
  assign _T_30278 = valid_32_13 ? 6'hd : _T_30277; // @[Mux.scala 31:69:@10555.4]
  assign _T_30279 = valid_32_12 ? 6'hc : _T_30278; // @[Mux.scala 31:69:@10556.4]
  assign _T_30280 = valid_32_11 ? 6'hb : _T_30279; // @[Mux.scala 31:69:@10557.4]
  assign _T_30281 = valid_32_10 ? 6'ha : _T_30280; // @[Mux.scala 31:69:@10558.4]
  assign _T_30282 = valid_32_9 ? 6'h9 : _T_30281; // @[Mux.scala 31:69:@10559.4]
  assign _T_30283 = valid_32_8 ? 6'h8 : _T_30282; // @[Mux.scala 31:69:@10560.4]
  assign _T_30284 = valid_32_7 ? 6'h7 : _T_30283; // @[Mux.scala 31:69:@10561.4]
  assign _T_30285 = valid_32_6 ? 6'h6 : _T_30284; // @[Mux.scala 31:69:@10562.4]
  assign _T_30286 = valid_32_5 ? 6'h5 : _T_30285; // @[Mux.scala 31:69:@10563.4]
  assign _T_30287 = valid_32_4 ? 6'h4 : _T_30286; // @[Mux.scala 31:69:@10564.4]
  assign _T_30288 = valid_32_3 ? 6'h3 : _T_30287; // @[Mux.scala 31:69:@10565.4]
  assign _T_30289 = valid_32_2 ? 6'h2 : _T_30288; // @[Mux.scala 31:69:@10566.4]
  assign _T_30290 = valid_32_1 ? 6'h1 : _T_30289; // @[Mux.scala 31:69:@10567.4]
  assign select_32 = valid_32_0 ? 6'h0 : _T_30290; // @[Mux.scala 31:69:@10568.4]
  assign _GEN_2049 = 6'h1 == select_32 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2050 = 6'h2 == select_32 ? io_inData_2 : _GEN_2049; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2051 = 6'h3 == select_32 ? io_inData_3 : _GEN_2050; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2052 = 6'h4 == select_32 ? io_inData_4 : _GEN_2051; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2053 = 6'h5 == select_32 ? io_inData_5 : _GEN_2052; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2054 = 6'h6 == select_32 ? io_inData_6 : _GEN_2053; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2055 = 6'h7 == select_32 ? io_inData_7 : _GEN_2054; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2056 = 6'h8 == select_32 ? io_inData_8 : _GEN_2055; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2057 = 6'h9 == select_32 ? io_inData_9 : _GEN_2056; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2058 = 6'ha == select_32 ? io_inData_10 : _GEN_2057; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2059 = 6'hb == select_32 ? io_inData_11 : _GEN_2058; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2060 = 6'hc == select_32 ? io_inData_12 : _GEN_2059; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2061 = 6'hd == select_32 ? io_inData_13 : _GEN_2060; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2062 = 6'he == select_32 ? io_inData_14 : _GEN_2061; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2063 = 6'hf == select_32 ? io_inData_15 : _GEN_2062; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2064 = 6'h10 == select_32 ? io_inData_16 : _GEN_2063; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2065 = 6'h11 == select_32 ? io_inData_17 : _GEN_2064; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2066 = 6'h12 == select_32 ? io_inData_18 : _GEN_2065; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2067 = 6'h13 == select_32 ? io_inData_19 : _GEN_2066; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2068 = 6'h14 == select_32 ? io_inData_20 : _GEN_2067; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2069 = 6'h15 == select_32 ? io_inData_21 : _GEN_2068; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2070 = 6'h16 == select_32 ? io_inData_22 : _GEN_2069; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2071 = 6'h17 == select_32 ? io_inData_23 : _GEN_2070; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2072 = 6'h18 == select_32 ? io_inData_24 : _GEN_2071; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2073 = 6'h19 == select_32 ? io_inData_25 : _GEN_2072; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2074 = 6'h1a == select_32 ? io_inData_26 : _GEN_2073; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2075 = 6'h1b == select_32 ? io_inData_27 : _GEN_2074; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2076 = 6'h1c == select_32 ? io_inData_28 : _GEN_2075; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2077 = 6'h1d == select_32 ? io_inData_29 : _GEN_2076; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2078 = 6'h1e == select_32 ? io_inData_30 : _GEN_2077; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2079 = 6'h1f == select_32 ? io_inData_31 : _GEN_2078; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2080 = 6'h20 == select_32 ? io_inData_32 : _GEN_2079; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2081 = 6'h21 == select_32 ? io_inData_33 : _GEN_2080; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2082 = 6'h22 == select_32 ? io_inData_34 : _GEN_2081; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2083 = 6'h23 == select_32 ? io_inData_35 : _GEN_2082; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2084 = 6'h24 == select_32 ? io_inData_36 : _GEN_2083; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2085 = 6'h25 == select_32 ? io_inData_37 : _GEN_2084; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2086 = 6'h26 == select_32 ? io_inData_38 : _GEN_2085; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2087 = 6'h27 == select_32 ? io_inData_39 : _GEN_2086; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2088 = 6'h28 == select_32 ? io_inData_40 : _GEN_2087; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2089 = 6'h29 == select_32 ? io_inData_41 : _GEN_2088; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2090 = 6'h2a == select_32 ? io_inData_42 : _GEN_2089; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2091 = 6'h2b == select_32 ? io_inData_43 : _GEN_2090; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2092 = 6'h2c == select_32 ? io_inData_44 : _GEN_2091; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2093 = 6'h2d == select_32 ? io_inData_45 : _GEN_2092; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2094 = 6'h2e == select_32 ? io_inData_46 : _GEN_2093; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2095 = 6'h2f == select_32 ? io_inData_47 : _GEN_2094; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2096 = 6'h30 == select_32 ? io_inData_48 : _GEN_2095; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2097 = 6'h31 == select_32 ? io_inData_49 : _GEN_2096; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2098 = 6'h32 == select_32 ? io_inData_50 : _GEN_2097; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2099 = 6'h33 == select_32 ? io_inData_51 : _GEN_2098; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2100 = 6'h34 == select_32 ? io_inData_52 : _GEN_2099; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2101 = 6'h35 == select_32 ? io_inData_53 : _GEN_2100; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2102 = 6'h36 == select_32 ? io_inData_54 : _GEN_2101; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2103 = 6'h37 == select_32 ? io_inData_55 : _GEN_2102; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2104 = 6'h38 == select_32 ? io_inData_56 : _GEN_2103; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2105 = 6'h39 == select_32 ? io_inData_57 : _GEN_2104; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2106 = 6'h3a == select_32 ? io_inData_58 : _GEN_2105; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2107 = 6'h3b == select_32 ? io_inData_59 : _GEN_2106; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2108 = 6'h3c == select_32 ? io_inData_60 : _GEN_2107; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2109 = 6'h3d == select_32 ? io_inData_61 : _GEN_2108; // @[Switch.scala 33:19:@10570.4]
  assign _GEN_2110 = 6'h3e == select_32 ? io_inData_62 : _GEN_2109; // @[Switch.scala 33:19:@10570.4]
  assign _T_30299 = {valid_32_7,valid_32_6,valid_32_5,valid_32_4,valid_32_3,valid_32_2,valid_32_1,valid_32_0}; // @[Switch.scala 34:32:@10577.4]
  assign _T_30307 = {valid_32_15,valid_32_14,valid_32_13,valid_32_12,valid_32_11,valid_32_10,valid_32_9,valid_32_8,_T_30299}; // @[Switch.scala 34:32:@10585.4]
  assign _T_30314 = {valid_32_23,valid_32_22,valid_32_21,valid_32_20,valid_32_19,valid_32_18,valid_32_17,valid_32_16}; // @[Switch.scala 34:32:@10592.4]
  assign _T_30323 = {valid_32_31,valid_32_30,valid_32_29,valid_32_28,valid_32_27,valid_32_26,valid_32_25,valid_32_24,_T_30314,_T_30307}; // @[Switch.scala 34:32:@10601.4]
  assign _T_30330 = {valid_32_39,valid_32_38,valid_32_37,valid_32_36,valid_32_35,valid_32_34,valid_32_33,valid_32_32}; // @[Switch.scala 34:32:@10608.4]
  assign _T_30338 = {valid_32_47,valid_32_46,valid_32_45,valid_32_44,valid_32_43,valid_32_42,valid_32_41,valid_32_40,_T_30330}; // @[Switch.scala 34:32:@10616.4]
  assign _T_30345 = {valid_32_55,valid_32_54,valid_32_53,valid_32_52,valid_32_51,valid_32_50,valid_32_49,valid_32_48}; // @[Switch.scala 34:32:@10623.4]
  assign _T_30354 = {valid_32_63,valid_32_62,valid_32_61,valid_32_60,valid_32_59,valid_32_58,valid_32_57,valid_32_56,_T_30345,_T_30338}; // @[Switch.scala 34:32:@10632.4]
  assign _T_30355 = {_T_30354,_T_30323}; // @[Switch.scala 34:32:@10633.4]
  assign _T_30359 = io_inAddr_0 == 6'h21; // @[Switch.scala 30:53:@10636.4]
  assign valid_33_0 = io_inValid_0 & _T_30359; // @[Switch.scala 30:36:@10637.4]
  assign _T_30362 = io_inAddr_1 == 6'h21; // @[Switch.scala 30:53:@10639.4]
  assign valid_33_1 = io_inValid_1 & _T_30362; // @[Switch.scala 30:36:@10640.4]
  assign _T_30365 = io_inAddr_2 == 6'h21; // @[Switch.scala 30:53:@10642.4]
  assign valid_33_2 = io_inValid_2 & _T_30365; // @[Switch.scala 30:36:@10643.4]
  assign _T_30368 = io_inAddr_3 == 6'h21; // @[Switch.scala 30:53:@10645.4]
  assign valid_33_3 = io_inValid_3 & _T_30368; // @[Switch.scala 30:36:@10646.4]
  assign _T_30371 = io_inAddr_4 == 6'h21; // @[Switch.scala 30:53:@10648.4]
  assign valid_33_4 = io_inValid_4 & _T_30371; // @[Switch.scala 30:36:@10649.4]
  assign _T_30374 = io_inAddr_5 == 6'h21; // @[Switch.scala 30:53:@10651.4]
  assign valid_33_5 = io_inValid_5 & _T_30374; // @[Switch.scala 30:36:@10652.4]
  assign _T_30377 = io_inAddr_6 == 6'h21; // @[Switch.scala 30:53:@10654.4]
  assign valid_33_6 = io_inValid_6 & _T_30377; // @[Switch.scala 30:36:@10655.4]
  assign _T_30380 = io_inAddr_7 == 6'h21; // @[Switch.scala 30:53:@10657.4]
  assign valid_33_7 = io_inValid_7 & _T_30380; // @[Switch.scala 30:36:@10658.4]
  assign _T_30383 = io_inAddr_8 == 6'h21; // @[Switch.scala 30:53:@10660.4]
  assign valid_33_8 = io_inValid_8 & _T_30383; // @[Switch.scala 30:36:@10661.4]
  assign _T_30386 = io_inAddr_9 == 6'h21; // @[Switch.scala 30:53:@10663.4]
  assign valid_33_9 = io_inValid_9 & _T_30386; // @[Switch.scala 30:36:@10664.4]
  assign _T_30389 = io_inAddr_10 == 6'h21; // @[Switch.scala 30:53:@10666.4]
  assign valid_33_10 = io_inValid_10 & _T_30389; // @[Switch.scala 30:36:@10667.4]
  assign _T_30392 = io_inAddr_11 == 6'h21; // @[Switch.scala 30:53:@10669.4]
  assign valid_33_11 = io_inValid_11 & _T_30392; // @[Switch.scala 30:36:@10670.4]
  assign _T_30395 = io_inAddr_12 == 6'h21; // @[Switch.scala 30:53:@10672.4]
  assign valid_33_12 = io_inValid_12 & _T_30395; // @[Switch.scala 30:36:@10673.4]
  assign _T_30398 = io_inAddr_13 == 6'h21; // @[Switch.scala 30:53:@10675.4]
  assign valid_33_13 = io_inValid_13 & _T_30398; // @[Switch.scala 30:36:@10676.4]
  assign _T_30401 = io_inAddr_14 == 6'h21; // @[Switch.scala 30:53:@10678.4]
  assign valid_33_14 = io_inValid_14 & _T_30401; // @[Switch.scala 30:36:@10679.4]
  assign _T_30404 = io_inAddr_15 == 6'h21; // @[Switch.scala 30:53:@10681.4]
  assign valid_33_15 = io_inValid_15 & _T_30404; // @[Switch.scala 30:36:@10682.4]
  assign _T_30407 = io_inAddr_16 == 6'h21; // @[Switch.scala 30:53:@10684.4]
  assign valid_33_16 = io_inValid_16 & _T_30407; // @[Switch.scala 30:36:@10685.4]
  assign _T_30410 = io_inAddr_17 == 6'h21; // @[Switch.scala 30:53:@10687.4]
  assign valid_33_17 = io_inValid_17 & _T_30410; // @[Switch.scala 30:36:@10688.4]
  assign _T_30413 = io_inAddr_18 == 6'h21; // @[Switch.scala 30:53:@10690.4]
  assign valid_33_18 = io_inValid_18 & _T_30413; // @[Switch.scala 30:36:@10691.4]
  assign _T_30416 = io_inAddr_19 == 6'h21; // @[Switch.scala 30:53:@10693.4]
  assign valid_33_19 = io_inValid_19 & _T_30416; // @[Switch.scala 30:36:@10694.4]
  assign _T_30419 = io_inAddr_20 == 6'h21; // @[Switch.scala 30:53:@10696.4]
  assign valid_33_20 = io_inValid_20 & _T_30419; // @[Switch.scala 30:36:@10697.4]
  assign _T_30422 = io_inAddr_21 == 6'h21; // @[Switch.scala 30:53:@10699.4]
  assign valid_33_21 = io_inValid_21 & _T_30422; // @[Switch.scala 30:36:@10700.4]
  assign _T_30425 = io_inAddr_22 == 6'h21; // @[Switch.scala 30:53:@10702.4]
  assign valid_33_22 = io_inValid_22 & _T_30425; // @[Switch.scala 30:36:@10703.4]
  assign _T_30428 = io_inAddr_23 == 6'h21; // @[Switch.scala 30:53:@10705.4]
  assign valid_33_23 = io_inValid_23 & _T_30428; // @[Switch.scala 30:36:@10706.4]
  assign _T_30431 = io_inAddr_24 == 6'h21; // @[Switch.scala 30:53:@10708.4]
  assign valid_33_24 = io_inValid_24 & _T_30431; // @[Switch.scala 30:36:@10709.4]
  assign _T_30434 = io_inAddr_25 == 6'h21; // @[Switch.scala 30:53:@10711.4]
  assign valid_33_25 = io_inValid_25 & _T_30434; // @[Switch.scala 30:36:@10712.4]
  assign _T_30437 = io_inAddr_26 == 6'h21; // @[Switch.scala 30:53:@10714.4]
  assign valid_33_26 = io_inValid_26 & _T_30437; // @[Switch.scala 30:36:@10715.4]
  assign _T_30440 = io_inAddr_27 == 6'h21; // @[Switch.scala 30:53:@10717.4]
  assign valid_33_27 = io_inValid_27 & _T_30440; // @[Switch.scala 30:36:@10718.4]
  assign _T_30443 = io_inAddr_28 == 6'h21; // @[Switch.scala 30:53:@10720.4]
  assign valid_33_28 = io_inValid_28 & _T_30443; // @[Switch.scala 30:36:@10721.4]
  assign _T_30446 = io_inAddr_29 == 6'h21; // @[Switch.scala 30:53:@10723.4]
  assign valid_33_29 = io_inValid_29 & _T_30446; // @[Switch.scala 30:36:@10724.4]
  assign _T_30449 = io_inAddr_30 == 6'h21; // @[Switch.scala 30:53:@10726.4]
  assign valid_33_30 = io_inValid_30 & _T_30449; // @[Switch.scala 30:36:@10727.4]
  assign _T_30452 = io_inAddr_31 == 6'h21; // @[Switch.scala 30:53:@10729.4]
  assign valid_33_31 = io_inValid_31 & _T_30452; // @[Switch.scala 30:36:@10730.4]
  assign _T_30455 = io_inAddr_32 == 6'h21; // @[Switch.scala 30:53:@10732.4]
  assign valid_33_32 = io_inValid_32 & _T_30455; // @[Switch.scala 30:36:@10733.4]
  assign _T_30458 = io_inAddr_33 == 6'h21; // @[Switch.scala 30:53:@10735.4]
  assign valid_33_33 = io_inValid_33 & _T_30458; // @[Switch.scala 30:36:@10736.4]
  assign _T_30461 = io_inAddr_34 == 6'h21; // @[Switch.scala 30:53:@10738.4]
  assign valid_33_34 = io_inValid_34 & _T_30461; // @[Switch.scala 30:36:@10739.4]
  assign _T_30464 = io_inAddr_35 == 6'h21; // @[Switch.scala 30:53:@10741.4]
  assign valid_33_35 = io_inValid_35 & _T_30464; // @[Switch.scala 30:36:@10742.4]
  assign _T_30467 = io_inAddr_36 == 6'h21; // @[Switch.scala 30:53:@10744.4]
  assign valid_33_36 = io_inValid_36 & _T_30467; // @[Switch.scala 30:36:@10745.4]
  assign _T_30470 = io_inAddr_37 == 6'h21; // @[Switch.scala 30:53:@10747.4]
  assign valid_33_37 = io_inValid_37 & _T_30470; // @[Switch.scala 30:36:@10748.4]
  assign _T_30473 = io_inAddr_38 == 6'h21; // @[Switch.scala 30:53:@10750.4]
  assign valid_33_38 = io_inValid_38 & _T_30473; // @[Switch.scala 30:36:@10751.4]
  assign _T_30476 = io_inAddr_39 == 6'h21; // @[Switch.scala 30:53:@10753.4]
  assign valid_33_39 = io_inValid_39 & _T_30476; // @[Switch.scala 30:36:@10754.4]
  assign _T_30479 = io_inAddr_40 == 6'h21; // @[Switch.scala 30:53:@10756.4]
  assign valid_33_40 = io_inValid_40 & _T_30479; // @[Switch.scala 30:36:@10757.4]
  assign _T_30482 = io_inAddr_41 == 6'h21; // @[Switch.scala 30:53:@10759.4]
  assign valid_33_41 = io_inValid_41 & _T_30482; // @[Switch.scala 30:36:@10760.4]
  assign _T_30485 = io_inAddr_42 == 6'h21; // @[Switch.scala 30:53:@10762.4]
  assign valid_33_42 = io_inValid_42 & _T_30485; // @[Switch.scala 30:36:@10763.4]
  assign _T_30488 = io_inAddr_43 == 6'h21; // @[Switch.scala 30:53:@10765.4]
  assign valid_33_43 = io_inValid_43 & _T_30488; // @[Switch.scala 30:36:@10766.4]
  assign _T_30491 = io_inAddr_44 == 6'h21; // @[Switch.scala 30:53:@10768.4]
  assign valid_33_44 = io_inValid_44 & _T_30491; // @[Switch.scala 30:36:@10769.4]
  assign _T_30494 = io_inAddr_45 == 6'h21; // @[Switch.scala 30:53:@10771.4]
  assign valid_33_45 = io_inValid_45 & _T_30494; // @[Switch.scala 30:36:@10772.4]
  assign _T_30497 = io_inAddr_46 == 6'h21; // @[Switch.scala 30:53:@10774.4]
  assign valid_33_46 = io_inValid_46 & _T_30497; // @[Switch.scala 30:36:@10775.4]
  assign _T_30500 = io_inAddr_47 == 6'h21; // @[Switch.scala 30:53:@10777.4]
  assign valid_33_47 = io_inValid_47 & _T_30500; // @[Switch.scala 30:36:@10778.4]
  assign _T_30503 = io_inAddr_48 == 6'h21; // @[Switch.scala 30:53:@10780.4]
  assign valid_33_48 = io_inValid_48 & _T_30503; // @[Switch.scala 30:36:@10781.4]
  assign _T_30506 = io_inAddr_49 == 6'h21; // @[Switch.scala 30:53:@10783.4]
  assign valid_33_49 = io_inValid_49 & _T_30506; // @[Switch.scala 30:36:@10784.4]
  assign _T_30509 = io_inAddr_50 == 6'h21; // @[Switch.scala 30:53:@10786.4]
  assign valid_33_50 = io_inValid_50 & _T_30509; // @[Switch.scala 30:36:@10787.4]
  assign _T_30512 = io_inAddr_51 == 6'h21; // @[Switch.scala 30:53:@10789.4]
  assign valid_33_51 = io_inValid_51 & _T_30512; // @[Switch.scala 30:36:@10790.4]
  assign _T_30515 = io_inAddr_52 == 6'h21; // @[Switch.scala 30:53:@10792.4]
  assign valid_33_52 = io_inValid_52 & _T_30515; // @[Switch.scala 30:36:@10793.4]
  assign _T_30518 = io_inAddr_53 == 6'h21; // @[Switch.scala 30:53:@10795.4]
  assign valid_33_53 = io_inValid_53 & _T_30518; // @[Switch.scala 30:36:@10796.4]
  assign _T_30521 = io_inAddr_54 == 6'h21; // @[Switch.scala 30:53:@10798.4]
  assign valid_33_54 = io_inValid_54 & _T_30521; // @[Switch.scala 30:36:@10799.4]
  assign _T_30524 = io_inAddr_55 == 6'h21; // @[Switch.scala 30:53:@10801.4]
  assign valid_33_55 = io_inValid_55 & _T_30524; // @[Switch.scala 30:36:@10802.4]
  assign _T_30527 = io_inAddr_56 == 6'h21; // @[Switch.scala 30:53:@10804.4]
  assign valid_33_56 = io_inValid_56 & _T_30527; // @[Switch.scala 30:36:@10805.4]
  assign _T_30530 = io_inAddr_57 == 6'h21; // @[Switch.scala 30:53:@10807.4]
  assign valid_33_57 = io_inValid_57 & _T_30530; // @[Switch.scala 30:36:@10808.4]
  assign _T_30533 = io_inAddr_58 == 6'h21; // @[Switch.scala 30:53:@10810.4]
  assign valid_33_58 = io_inValid_58 & _T_30533; // @[Switch.scala 30:36:@10811.4]
  assign _T_30536 = io_inAddr_59 == 6'h21; // @[Switch.scala 30:53:@10813.4]
  assign valid_33_59 = io_inValid_59 & _T_30536; // @[Switch.scala 30:36:@10814.4]
  assign _T_30539 = io_inAddr_60 == 6'h21; // @[Switch.scala 30:53:@10816.4]
  assign valid_33_60 = io_inValid_60 & _T_30539; // @[Switch.scala 30:36:@10817.4]
  assign _T_30542 = io_inAddr_61 == 6'h21; // @[Switch.scala 30:53:@10819.4]
  assign valid_33_61 = io_inValid_61 & _T_30542; // @[Switch.scala 30:36:@10820.4]
  assign _T_30545 = io_inAddr_62 == 6'h21; // @[Switch.scala 30:53:@10822.4]
  assign valid_33_62 = io_inValid_62 & _T_30545; // @[Switch.scala 30:36:@10823.4]
  assign _T_30548 = io_inAddr_63 == 6'h21; // @[Switch.scala 30:53:@10825.4]
  assign valid_33_63 = io_inValid_63 & _T_30548; // @[Switch.scala 30:36:@10826.4]
  assign _T_30614 = valid_33_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@10828.4]
  assign _T_30615 = valid_33_61 ? 6'h3d : _T_30614; // @[Mux.scala 31:69:@10829.4]
  assign _T_30616 = valid_33_60 ? 6'h3c : _T_30615; // @[Mux.scala 31:69:@10830.4]
  assign _T_30617 = valid_33_59 ? 6'h3b : _T_30616; // @[Mux.scala 31:69:@10831.4]
  assign _T_30618 = valid_33_58 ? 6'h3a : _T_30617; // @[Mux.scala 31:69:@10832.4]
  assign _T_30619 = valid_33_57 ? 6'h39 : _T_30618; // @[Mux.scala 31:69:@10833.4]
  assign _T_30620 = valid_33_56 ? 6'h38 : _T_30619; // @[Mux.scala 31:69:@10834.4]
  assign _T_30621 = valid_33_55 ? 6'h37 : _T_30620; // @[Mux.scala 31:69:@10835.4]
  assign _T_30622 = valid_33_54 ? 6'h36 : _T_30621; // @[Mux.scala 31:69:@10836.4]
  assign _T_30623 = valid_33_53 ? 6'h35 : _T_30622; // @[Mux.scala 31:69:@10837.4]
  assign _T_30624 = valid_33_52 ? 6'h34 : _T_30623; // @[Mux.scala 31:69:@10838.4]
  assign _T_30625 = valid_33_51 ? 6'h33 : _T_30624; // @[Mux.scala 31:69:@10839.4]
  assign _T_30626 = valid_33_50 ? 6'h32 : _T_30625; // @[Mux.scala 31:69:@10840.4]
  assign _T_30627 = valid_33_49 ? 6'h31 : _T_30626; // @[Mux.scala 31:69:@10841.4]
  assign _T_30628 = valid_33_48 ? 6'h30 : _T_30627; // @[Mux.scala 31:69:@10842.4]
  assign _T_30629 = valid_33_47 ? 6'h2f : _T_30628; // @[Mux.scala 31:69:@10843.4]
  assign _T_30630 = valid_33_46 ? 6'h2e : _T_30629; // @[Mux.scala 31:69:@10844.4]
  assign _T_30631 = valid_33_45 ? 6'h2d : _T_30630; // @[Mux.scala 31:69:@10845.4]
  assign _T_30632 = valid_33_44 ? 6'h2c : _T_30631; // @[Mux.scala 31:69:@10846.4]
  assign _T_30633 = valid_33_43 ? 6'h2b : _T_30632; // @[Mux.scala 31:69:@10847.4]
  assign _T_30634 = valid_33_42 ? 6'h2a : _T_30633; // @[Mux.scala 31:69:@10848.4]
  assign _T_30635 = valid_33_41 ? 6'h29 : _T_30634; // @[Mux.scala 31:69:@10849.4]
  assign _T_30636 = valid_33_40 ? 6'h28 : _T_30635; // @[Mux.scala 31:69:@10850.4]
  assign _T_30637 = valid_33_39 ? 6'h27 : _T_30636; // @[Mux.scala 31:69:@10851.4]
  assign _T_30638 = valid_33_38 ? 6'h26 : _T_30637; // @[Mux.scala 31:69:@10852.4]
  assign _T_30639 = valid_33_37 ? 6'h25 : _T_30638; // @[Mux.scala 31:69:@10853.4]
  assign _T_30640 = valid_33_36 ? 6'h24 : _T_30639; // @[Mux.scala 31:69:@10854.4]
  assign _T_30641 = valid_33_35 ? 6'h23 : _T_30640; // @[Mux.scala 31:69:@10855.4]
  assign _T_30642 = valid_33_34 ? 6'h22 : _T_30641; // @[Mux.scala 31:69:@10856.4]
  assign _T_30643 = valid_33_33 ? 6'h21 : _T_30642; // @[Mux.scala 31:69:@10857.4]
  assign _T_30644 = valid_33_32 ? 6'h20 : _T_30643; // @[Mux.scala 31:69:@10858.4]
  assign _T_30645 = valid_33_31 ? 6'h1f : _T_30644; // @[Mux.scala 31:69:@10859.4]
  assign _T_30646 = valid_33_30 ? 6'h1e : _T_30645; // @[Mux.scala 31:69:@10860.4]
  assign _T_30647 = valid_33_29 ? 6'h1d : _T_30646; // @[Mux.scala 31:69:@10861.4]
  assign _T_30648 = valid_33_28 ? 6'h1c : _T_30647; // @[Mux.scala 31:69:@10862.4]
  assign _T_30649 = valid_33_27 ? 6'h1b : _T_30648; // @[Mux.scala 31:69:@10863.4]
  assign _T_30650 = valid_33_26 ? 6'h1a : _T_30649; // @[Mux.scala 31:69:@10864.4]
  assign _T_30651 = valid_33_25 ? 6'h19 : _T_30650; // @[Mux.scala 31:69:@10865.4]
  assign _T_30652 = valid_33_24 ? 6'h18 : _T_30651; // @[Mux.scala 31:69:@10866.4]
  assign _T_30653 = valid_33_23 ? 6'h17 : _T_30652; // @[Mux.scala 31:69:@10867.4]
  assign _T_30654 = valid_33_22 ? 6'h16 : _T_30653; // @[Mux.scala 31:69:@10868.4]
  assign _T_30655 = valid_33_21 ? 6'h15 : _T_30654; // @[Mux.scala 31:69:@10869.4]
  assign _T_30656 = valid_33_20 ? 6'h14 : _T_30655; // @[Mux.scala 31:69:@10870.4]
  assign _T_30657 = valid_33_19 ? 6'h13 : _T_30656; // @[Mux.scala 31:69:@10871.4]
  assign _T_30658 = valid_33_18 ? 6'h12 : _T_30657; // @[Mux.scala 31:69:@10872.4]
  assign _T_30659 = valid_33_17 ? 6'h11 : _T_30658; // @[Mux.scala 31:69:@10873.4]
  assign _T_30660 = valid_33_16 ? 6'h10 : _T_30659; // @[Mux.scala 31:69:@10874.4]
  assign _T_30661 = valid_33_15 ? 6'hf : _T_30660; // @[Mux.scala 31:69:@10875.4]
  assign _T_30662 = valid_33_14 ? 6'he : _T_30661; // @[Mux.scala 31:69:@10876.4]
  assign _T_30663 = valid_33_13 ? 6'hd : _T_30662; // @[Mux.scala 31:69:@10877.4]
  assign _T_30664 = valid_33_12 ? 6'hc : _T_30663; // @[Mux.scala 31:69:@10878.4]
  assign _T_30665 = valid_33_11 ? 6'hb : _T_30664; // @[Mux.scala 31:69:@10879.4]
  assign _T_30666 = valid_33_10 ? 6'ha : _T_30665; // @[Mux.scala 31:69:@10880.4]
  assign _T_30667 = valid_33_9 ? 6'h9 : _T_30666; // @[Mux.scala 31:69:@10881.4]
  assign _T_30668 = valid_33_8 ? 6'h8 : _T_30667; // @[Mux.scala 31:69:@10882.4]
  assign _T_30669 = valid_33_7 ? 6'h7 : _T_30668; // @[Mux.scala 31:69:@10883.4]
  assign _T_30670 = valid_33_6 ? 6'h6 : _T_30669; // @[Mux.scala 31:69:@10884.4]
  assign _T_30671 = valid_33_5 ? 6'h5 : _T_30670; // @[Mux.scala 31:69:@10885.4]
  assign _T_30672 = valid_33_4 ? 6'h4 : _T_30671; // @[Mux.scala 31:69:@10886.4]
  assign _T_30673 = valid_33_3 ? 6'h3 : _T_30672; // @[Mux.scala 31:69:@10887.4]
  assign _T_30674 = valid_33_2 ? 6'h2 : _T_30673; // @[Mux.scala 31:69:@10888.4]
  assign _T_30675 = valid_33_1 ? 6'h1 : _T_30674; // @[Mux.scala 31:69:@10889.4]
  assign select_33 = valid_33_0 ? 6'h0 : _T_30675; // @[Mux.scala 31:69:@10890.4]
  assign _GEN_2113 = 6'h1 == select_33 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2114 = 6'h2 == select_33 ? io_inData_2 : _GEN_2113; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2115 = 6'h3 == select_33 ? io_inData_3 : _GEN_2114; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2116 = 6'h4 == select_33 ? io_inData_4 : _GEN_2115; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2117 = 6'h5 == select_33 ? io_inData_5 : _GEN_2116; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2118 = 6'h6 == select_33 ? io_inData_6 : _GEN_2117; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2119 = 6'h7 == select_33 ? io_inData_7 : _GEN_2118; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2120 = 6'h8 == select_33 ? io_inData_8 : _GEN_2119; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2121 = 6'h9 == select_33 ? io_inData_9 : _GEN_2120; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2122 = 6'ha == select_33 ? io_inData_10 : _GEN_2121; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2123 = 6'hb == select_33 ? io_inData_11 : _GEN_2122; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2124 = 6'hc == select_33 ? io_inData_12 : _GEN_2123; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2125 = 6'hd == select_33 ? io_inData_13 : _GEN_2124; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2126 = 6'he == select_33 ? io_inData_14 : _GEN_2125; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2127 = 6'hf == select_33 ? io_inData_15 : _GEN_2126; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2128 = 6'h10 == select_33 ? io_inData_16 : _GEN_2127; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2129 = 6'h11 == select_33 ? io_inData_17 : _GEN_2128; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2130 = 6'h12 == select_33 ? io_inData_18 : _GEN_2129; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2131 = 6'h13 == select_33 ? io_inData_19 : _GEN_2130; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2132 = 6'h14 == select_33 ? io_inData_20 : _GEN_2131; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2133 = 6'h15 == select_33 ? io_inData_21 : _GEN_2132; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2134 = 6'h16 == select_33 ? io_inData_22 : _GEN_2133; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2135 = 6'h17 == select_33 ? io_inData_23 : _GEN_2134; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2136 = 6'h18 == select_33 ? io_inData_24 : _GEN_2135; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2137 = 6'h19 == select_33 ? io_inData_25 : _GEN_2136; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2138 = 6'h1a == select_33 ? io_inData_26 : _GEN_2137; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2139 = 6'h1b == select_33 ? io_inData_27 : _GEN_2138; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2140 = 6'h1c == select_33 ? io_inData_28 : _GEN_2139; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2141 = 6'h1d == select_33 ? io_inData_29 : _GEN_2140; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2142 = 6'h1e == select_33 ? io_inData_30 : _GEN_2141; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2143 = 6'h1f == select_33 ? io_inData_31 : _GEN_2142; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2144 = 6'h20 == select_33 ? io_inData_32 : _GEN_2143; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2145 = 6'h21 == select_33 ? io_inData_33 : _GEN_2144; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2146 = 6'h22 == select_33 ? io_inData_34 : _GEN_2145; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2147 = 6'h23 == select_33 ? io_inData_35 : _GEN_2146; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2148 = 6'h24 == select_33 ? io_inData_36 : _GEN_2147; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2149 = 6'h25 == select_33 ? io_inData_37 : _GEN_2148; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2150 = 6'h26 == select_33 ? io_inData_38 : _GEN_2149; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2151 = 6'h27 == select_33 ? io_inData_39 : _GEN_2150; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2152 = 6'h28 == select_33 ? io_inData_40 : _GEN_2151; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2153 = 6'h29 == select_33 ? io_inData_41 : _GEN_2152; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2154 = 6'h2a == select_33 ? io_inData_42 : _GEN_2153; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2155 = 6'h2b == select_33 ? io_inData_43 : _GEN_2154; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2156 = 6'h2c == select_33 ? io_inData_44 : _GEN_2155; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2157 = 6'h2d == select_33 ? io_inData_45 : _GEN_2156; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2158 = 6'h2e == select_33 ? io_inData_46 : _GEN_2157; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2159 = 6'h2f == select_33 ? io_inData_47 : _GEN_2158; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2160 = 6'h30 == select_33 ? io_inData_48 : _GEN_2159; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2161 = 6'h31 == select_33 ? io_inData_49 : _GEN_2160; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2162 = 6'h32 == select_33 ? io_inData_50 : _GEN_2161; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2163 = 6'h33 == select_33 ? io_inData_51 : _GEN_2162; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2164 = 6'h34 == select_33 ? io_inData_52 : _GEN_2163; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2165 = 6'h35 == select_33 ? io_inData_53 : _GEN_2164; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2166 = 6'h36 == select_33 ? io_inData_54 : _GEN_2165; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2167 = 6'h37 == select_33 ? io_inData_55 : _GEN_2166; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2168 = 6'h38 == select_33 ? io_inData_56 : _GEN_2167; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2169 = 6'h39 == select_33 ? io_inData_57 : _GEN_2168; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2170 = 6'h3a == select_33 ? io_inData_58 : _GEN_2169; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2171 = 6'h3b == select_33 ? io_inData_59 : _GEN_2170; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2172 = 6'h3c == select_33 ? io_inData_60 : _GEN_2171; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2173 = 6'h3d == select_33 ? io_inData_61 : _GEN_2172; // @[Switch.scala 33:19:@10892.4]
  assign _GEN_2174 = 6'h3e == select_33 ? io_inData_62 : _GEN_2173; // @[Switch.scala 33:19:@10892.4]
  assign _T_30684 = {valid_33_7,valid_33_6,valid_33_5,valid_33_4,valid_33_3,valid_33_2,valid_33_1,valid_33_0}; // @[Switch.scala 34:32:@10899.4]
  assign _T_30692 = {valid_33_15,valid_33_14,valid_33_13,valid_33_12,valid_33_11,valid_33_10,valid_33_9,valid_33_8,_T_30684}; // @[Switch.scala 34:32:@10907.4]
  assign _T_30699 = {valid_33_23,valid_33_22,valid_33_21,valid_33_20,valid_33_19,valid_33_18,valid_33_17,valid_33_16}; // @[Switch.scala 34:32:@10914.4]
  assign _T_30708 = {valid_33_31,valid_33_30,valid_33_29,valid_33_28,valid_33_27,valid_33_26,valid_33_25,valid_33_24,_T_30699,_T_30692}; // @[Switch.scala 34:32:@10923.4]
  assign _T_30715 = {valid_33_39,valid_33_38,valid_33_37,valid_33_36,valid_33_35,valid_33_34,valid_33_33,valid_33_32}; // @[Switch.scala 34:32:@10930.4]
  assign _T_30723 = {valid_33_47,valid_33_46,valid_33_45,valid_33_44,valid_33_43,valid_33_42,valid_33_41,valid_33_40,_T_30715}; // @[Switch.scala 34:32:@10938.4]
  assign _T_30730 = {valid_33_55,valid_33_54,valid_33_53,valid_33_52,valid_33_51,valid_33_50,valid_33_49,valid_33_48}; // @[Switch.scala 34:32:@10945.4]
  assign _T_30739 = {valid_33_63,valid_33_62,valid_33_61,valid_33_60,valid_33_59,valid_33_58,valid_33_57,valid_33_56,_T_30730,_T_30723}; // @[Switch.scala 34:32:@10954.4]
  assign _T_30740 = {_T_30739,_T_30708}; // @[Switch.scala 34:32:@10955.4]
  assign _T_30744 = io_inAddr_0 == 6'h22; // @[Switch.scala 30:53:@10958.4]
  assign valid_34_0 = io_inValid_0 & _T_30744; // @[Switch.scala 30:36:@10959.4]
  assign _T_30747 = io_inAddr_1 == 6'h22; // @[Switch.scala 30:53:@10961.4]
  assign valid_34_1 = io_inValid_1 & _T_30747; // @[Switch.scala 30:36:@10962.4]
  assign _T_30750 = io_inAddr_2 == 6'h22; // @[Switch.scala 30:53:@10964.4]
  assign valid_34_2 = io_inValid_2 & _T_30750; // @[Switch.scala 30:36:@10965.4]
  assign _T_30753 = io_inAddr_3 == 6'h22; // @[Switch.scala 30:53:@10967.4]
  assign valid_34_3 = io_inValid_3 & _T_30753; // @[Switch.scala 30:36:@10968.4]
  assign _T_30756 = io_inAddr_4 == 6'h22; // @[Switch.scala 30:53:@10970.4]
  assign valid_34_4 = io_inValid_4 & _T_30756; // @[Switch.scala 30:36:@10971.4]
  assign _T_30759 = io_inAddr_5 == 6'h22; // @[Switch.scala 30:53:@10973.4]
  assign valid_34_5 = io_inValid_5 & _T_30759; // @[Switch.scala 30:36:@10974.4]
  assign _T_30762 = io_inAddr_6 == 6'h22; // @[Switch.scala 30:53:@10976.4]
  assign valid_34_6 = io_inValid_6 & _T_30762; // @[Switch.scala 30:36:@10977.4]
  assign _T_30765 = io_inAddr_7 == 6'h22; // @[Switch.scala 30:53:@10979.4]
  assign valid_34_7 = io_inValid_7 & _T_30765; // @[Switch.scala 30:36:@10980.4]
  assign _T_30768 = io_inAddr_8 == 6'h22; // @[Switch.scala 30:53:@10982.4]
  assign valid_34_8 = io_inValid_8 & _T_30768; // @[Switch.scala 30:36:@10983.4]
  assign _T_30771 = io_inAddr_9 == 6'h22; // @[Switch.scala 30:53:@10985.4]
  assign valid_34_9 = io_inValid_9 & _T_30771; // @[Switch.scala 30:36:@10986.4]
  assign _T_30774 = io_inAddr_10 == 6'h22; // @[Switch.scala 30:53:@10988.4]
  assign valid_34_10 = io_inValid_10 & _T_30774; // @[Switch.scala 30:36:@10989.4]
  assign _T_30777 = io_inAddr_11 == 6'h22; // @[Switch.scala 30:53:@10991.4]
  assign valid_34_11 = io_inValid_11 & _T_30777; // @[Switch.scala 30:36:@10992.4]
  assign _T_30780 = io_inAddr_12 == 6'h22; // @[Switch.scala 30:53:@10994.4]
  assign valid_34_12 = io_inValid_12 & _T_30780; // @[Switch.scala 30:36:@10995.4]
  assign _T_30783 = io_inAddr_13 == 6'h22; // @[Switch.scala 30:53:@10997.4]
  assign valid_34_13 = io_inValid_13 & _T_30783; // @[Switch.scala 30:36:@10998.4]
  assign _T_30786 = io_inAddr_14 == 6'h22; // @[Switch.scala 30:53:@11000.4]
  assign valid_34_14 = io_inValid_14 & _T_30786; // @[Switch.scala 30:36:@11001.4]
  assign _T_30789 = io_inAddr_15 == 6'h22; // @[Switch.scala 30:53:@11003.4]
  assign valid_34_15 = io_inValid_15 & _T_30789; // @[Switch.scala 30:36:@11004.4]
  assign _T_30792 = io_inAddr_16 == 6'h22; // @[Switch.scala 30:53:@11006.4]
  assign valid_34_16 = io_inValid_16 & _T_30792; // @[Switch.scala 30:36:@11007.4]
  assign _T_30795 = io_inAddr_17 == 6'h22; // @[Switch.scala 30:53:@11009.4]
  assign valid_34_17 = io_inValid_17 & _T_30795; // @[Switch.scala 30:36:@11010.4]
  assign _T_30798 = io_inAddr_18 == 6'h22; // @[Switch.scala 30:53:@11012.4]
  assign valid_34_18 = io_inValid_18 & _T_30798; // @[Switch.scala 30:36:@11013.4]
  assign _T_30801 = io_inAddr_19 == 6'h22; // @[Switch.scala 30:53:@11015.4]
  assign valid_34_19 = io_inValid_19 & _T_30801; // @[Switch.scala 30:36:@11016.4]
  assign _T_30804 = io_inAddr_20 == 6'h22; // @[Switch.scala 30:53:@11018.4]
  assign valid_34_20 = io_inValid_20 & _T_30804; // @[Switch.scala 30:36:@11019.4]
  assign _T_30807 = io_inAddr_21 == 6'h22; // @[Switch.scala 30:53:@11021.4]
  assign valid_34_21 = io_inValid_21 & _T_30807; // @[Switch.scala 30:36:@11022.4]
  assign _T_30810 = io_inAddr_22 == 6'h22; // @[Switch.scala 30:53:@11024.4]
  assign valid_34_22 = io_inValid_22 & _T_30810; // @[Switch.scala 30:36:@11025.4]
  assign _T_30813 = io_inAddr_23 == 6'h22; // @[Switch.scala 30:53:@11027.4]
  assign valid_34_23 = io_inValid_23 & _T_30813; // @[Switch.scala 30:36:@11028.4]
  assign _T_30816 = io_inAddr_24 == 6'h22; // @[Switch.scala 30:53:@11030.4]
  assign valid_34_24 = io_inValid_24 & _T_30816; // @[Switch.scala 30:36:@11031.4]
  assign _T_30819 = io_inAddr_25 == 6'h22; // @[Switch.scala 30:53:@11033.4]
  assign valid_34_25 = io_inValid_25 & _T_30819; // @[Switch.scala 30:36:@11034.4]
  assign _T_30822 = io_inAddr_26 == 6'h22; // @[Switch.scala 30:53:@11036.4]
  assign valid_34_26 = io_inValid_26 & _T_30822; // @[Switch.scala 30:36:@11037.4]
  assign _T_30825 = io_inAddr_27 == 6'h22; // @[Switch.scala 30:53:@11039.4]
  assign valid_34_27 = io_inValid_27 & _T_30825; // @[Switch.scala 30:36:@11040.4]
  assign _T_30828 = io_inAddr_28 == 6'h22; // @[Switch.scala 30:53:@11042.4]
  assign valid_34_28 = io_inValid_28 & _T_30828; // @[Switch.scala 30:36:@11043.4]
  assign _T_30831 = io_inAddr_29 == 6'h22; // @[Switch.scala 30:53:@11045.4]
  assign valid_34_29 = io_inValid_29 & _T_30831; // @[Switch.scala 30:36:@11046.4]
  assign _T_30834 = io_inAddr_30 == 6'h22; // @[Switch.scala 30:53:@11048.4]
  assign valid_34_30 = io_inValid_30 & _T_30834; // @[Switch.scala 30:36:@11049.4]
  assign _T_30837 = io_inAddr_31 == 6'h22; // @[Switch.scala 30:53:@11051.4]
  assign valid_34_31 = io_inValid_31 & _T_30837; // @[Switch.scala 30:36:@11052.4]
  assign _T_30840 = io_inAddr_32 == 6'h22; // @[Switch.scala 30:53:@11054.4]
  assign valid_34_32 = io_inValid_32 & _T_30840; // @[Switch.scala 30:36:@11055.4]
  assign _T_30843 = io_inAddr_33 == 6'h22; // @[Switch.scala 30:53:@11057.4]
  assign valid_34_33 = io_inValid_33 & _T_30843; // @[Switch.scala 30:36:@11058.4]
  assign _T_30846 = io_inAddr_34 == 6'h22; // @[Switch.scala 30:53:@11060.4]
  assign valid_34_34 = io_inValid_34 & _T_30846; // @[Switch.scala 30:36:@11061.4]
  assign _T_30849 = io_inAddr_35 == 6'h22; // @[Switch.scala 30:53:@11063.4]
  assign valid_34_35 = io_inValid_35 & _T_30849; // @[Switch.scala 30:36:@11064.4]
  assign _T_30852 = io_inAddr_36 == 6'h22; // @[Switch.scala 30:53:@11066.4]
  assign valid_34_36 = io_inValid_36 & _T_30852; // @[Switch.scala 30:36:@11067.4]
  assign _T_30855 = io_inAddr_37 == 6'h22; // @[Switch.scala 30:53:@11069.4]
  assign valid_34_37 = io_inValid_37 & _T_30855; // @[Switch.scala 30:36:@11070.4]
  assign _T_30858 = io_inAddr_38 == 6'h22; // @[Switch.scala 30:53:@11072.4]
  assign valid_34_38 = io_inValid_38 & _T_30858; // @[Switch.scala 30:36:@11073.4]
  assign _T_30861 = io_inAddr_39 == 6'h22; // @[Switch.scala 30:53:@11075.4]
  assign valid_34_39 = io_inValid_39 & _T_30861; // @[Switch.scala 30:36:@11076.4]
  assign _T_30864 = io_inAddr_40 == 6'h22; // @[Switch.scala 30:53:@11078.4]
  assign valid_34_40 = io_inValid_40 & _T_30864; // @[Switch.scala 30:36:@11079.4]
  assign _T_30867 = io_inAddr_41 == 6'h22; // @[Switch.scala 30:53:@11081.4]
  assign valid_34_41 = io_inValid_41 & _T_30867; // @[Switch.scala 30:36:@11082.4]
  assign _T_30870 = io_inAddr_42 == 6'h22; // @[Switch.scala 30:53:@11084.4]
  assign valid_34_42 = io_inValid_42 & _T_30870; // @[Switch.scala 30:36:@11085.4]
  assign _T_30873 = io_inAddr_43 == 6'h22; // @[Switch.scala 30:53:@11087.4]
  assign valid_34_43 = io_inValid_43 & _T_30873; // @[Switch.scala 30:36:@11088.4]
  assign _T_30876 = io_inAddr_44 == 6'h22; // @[Switch.scala 30:53:@11090.4]
  assign valid_34_44 = io_inValid_44 & _T_30876; // @[Switch.scala 30:36:@11091.4]
  assign _T_30879 = io_inAddr_45 == 6'h22; // @[Switch.scala 30:53:@11093.4]
  assign valid_34_45 = io_inValid_45 & _T_30879; // @[Switch.scala 30:36:@11094.4]
  assign _T_30882 = io_inAddr_46 == 6'h22; // @[Switch.scala 30:53:@11096.4]
  assign valid_34_46 = io_inValid_46 & _T_30882; // @[Switch.scala 30:36:@11097.4]
  assign _T_30885 = io_inAddr_47 == 6'h22; // @[Switch.scala 30:53:@11099.4]
  assign valid_34_47 = io_inValid_47 & _T_30885; // @[Switch.scala 30:36:@11100.4]
  assign _T_30888 = io_inAddr_48 == 6'h22; // @[Switch.scala 30:53:@11102.4]
  assign valid_34_48 = io_inValid_48 & _T_30888; // @[Switch.scala 30:36:@11103.4]
  assign _T_30891 = io_inAddr_49 == 6'h22; // @[Switch.scala 30:53:@11105.4]
  assign valid_34_49 = io_inValid_49 & _T_30891; // @[Switch.scala 30:36:@11106.4]
  assign _T_30894 = io_inAddr_50 == 6'h22; // @[Switch.scala 30:53:@11108.4]
  assign valid_34_50 = io_inValid_50 & _T_30894; // @[Switch.scala 30:36:@11109.4]
  assign _T_30897 = io_inAddr_51 == 6'h22; // @[Switch.scala 30:53:@11111.4]
  assign valid_34_51 = io_inValid_51 & _T_30897; // @[Switch.scala 30:36:@11112.4]
  assign _T_30900 = io_inAddr_52 == 6'h22; // @[Switch.scala 30:53:@11114.4]
  assign valid_34_52 = io_inValid_52 & _T_30900; // @[Switch.scala 30:36:@11115.4]
  assign _T_30903 = io_inAddr_53 == 6'h22; // @[Switch.scala 30:53:@11117.4]
  assign valid_34_53 = io_inValid_53 & _T_30903; // @[Switch.scala 30:36:@11118.4]
  assign _T_30906 = io_inAddr_54 == 6'h22; // @[Switch.scala 30:53:@11120.4]
  assign valid_34_54 = io_inValid_54 & _T_30906; // @[Switch.scala 30:36:@11121.4]
  assign _T_30909 = io_inAddr_55 == 6'h22; // @[Switch.scala 30:53:@11123.4]
  assign valid_34_55 = io_inValid_55 & _T_30909; // @[Switch.scala 30:36:@11124.4]
  assign _T_30912 = io_inAddr_56 == 6'h22; // @[Switch.scala 30:53:@11126.4]
  assign valid_34_56 = io_inValid_56 & _T_30912; // @[Switch.scala 30:36:@11127.4]
  assign _T_30915 = io_inAddr_57 == 6'h22; // @[Switch.scala 30:53:@11129.4]
  assign valid_34_57 = io_inValid_57 & _T_30915; // @[Switch.scala 30:36:@11130.4]
  assign _T_30918 = io_inAddr_58 == 6'h22; // @[Switch.scala 30:53:@11132.4]
  assign valid_34_58 = io_inValid_58 & _T_30918; // @[Switch.scala 30:36:@11133.4]
  assign _T_30921 = io_inAddr_59 == 6'h22; // @[Switch.scala 30:53:@11135.4]
  assign valid_34_59 = io_inValid_59 & _T_30921; // @[Switch.scala 30:36:@11136.4]
  assign _T_30924 = io_inAddr_60 == 6'h22; // @[Switch.scala 30:53:@11138.4]
  assign valid_34_60 = io_inValid_60 & _T_30924; // @[Switch.scala 30:36:@11139.4]
  assign _T_30927 = io_inAddr_61 == 6'h22; // @[Switch.scala 30:53:@11141.4]
  assign valid_34_61 = io_inValid_61 & _T_30927; // @[Switch.scala 30:36:@11142.4]
  assign _T_30930 = io_inAddr_62 == 6'h22; // @[Switch.scala 30:53:@11144.4]
  assign valid_34_62 = io_inValid_62 & _T_30930; // @[Switch.scala 30:36:@11145.4]
  assign _T_30933 = io_inAddr_63 == 6'h22; // @[Switch.scala 30:53:@11147.4]
  assign valid_34_63 = io_inValid_63 & _T_30933; // @[Switch.scala 30:36:@11148.4]
  assign _T_30999 = valid_34_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@11150.4]
  assign _T_31000 = valid_34_61 ? 6'h3d : _T_30999; // @[Mux.scala 31:69:@11151.4]
  assign _T_31001 = valid_34_60 ? 6'h3c : _T_31000; // @[Mux.scala 31:69:@11152.4]
  assign _T_31002 = valid_34_59 ? 6'h3b : _T_31001; // @[Mux.scala 31:69:@11153.4]
  assign _T_31003 = valid_34_58 ? 6'h3a : _T_31002; // @[Mux.scala 31:69:@11154.4]
  assign _T_31004 = valid_34_57 ? 6'h39 : _T_31003; // @[Mux.scala 31:69:@11155.4]
  assign _T_31005 = valid_34_56 ? 6'h38 : _T_31004; // @[Mux.scala 31:69:@11156.4]
  assign _T_31006 = valid_34_55 ? 6'h37 : _T_31005; // @[Mux.scala 31:69:@11157.4]
  assign _T_31007 = valid_34_54 ? 6'h36 : _T_31006; // @[Mux.scala 31:69:@11158.4]
  assign _T_31008 = valid_34_53 ? 6'h35 : _T_31007; // @[Mux.scala 31:69:@11159.4]
  assign _T_31009 = valid_34_52 ? 6'h34 : _T_31008; // @[Mux.scala 31:69:@11160.4]
  assign _T_31010 = valid_34_51 ? 6'h33 : _T_31009; // @[Mux.scala 31:69:@11161.4]
  assign _T_31011 = valid_34_50 ? 6'h32 : _T_31010; // @[Mux.scala 31:69:@11162.4]
  assign _T_31012 = valid_34_49 ? 6'h31 : _T_31011; // @[Mux.scala 31:69:@11163.4]
  assign _T_31013 = valid_34_48 ? 6'h30 : _T_31012; // @[Mux.scala 31:69:@11164.4]
  assign _T_31014 = valid_34_47 ? 6'h2f : _T_31013; // @[Mux.scala 31:69:@11165.4]
  assign _T_31015 = valid_34_46 ? 6'h2e : _T_31014; // @[Mux.scala 31:69:@11166.4]
  assign _T_31016 = valid_34_45 ? 6'h2d : _T_31015; // @[Mux.scala 31:69:@11167.4]
  assign _T_31017 = valid_34_44 ? 6'h2c : _T_31016; // @[Mux.scala 31:69:@11168.4]
  assign _T_31018 = valid_34_43 ? 6'h2b : _T_31017; // @[Mux.scala 31:69:@11169.4]
  assign _T_31019 = valid_34_42 ? 6'h2a : _T_31018; // @[Mux.scala 31:69:@11170.4]
  assign _T_31020 = valid_34_41 ? 6'h29 : _T_31019; // @[Mux.scala 31:69:@11171.4]
  assign _T_31021 = valid_34_40 ? 6'h28 : _T_31020; // @[Mux.scala 31:69:@11172.4]
  assign _T_31022 = valid_34_39 ? 6'h27 : _T_31021; // @[Mux.scala 31:69:@11173.4]
  assign _T_31023 = valid_34_38 ? 6'h26 : _T_31022; // @[Mux.scala 31:69:@11174.4]
  assign _T_31024 = valid_34_37 ? 6'h25 : _T_31023; // @[Mux.scala 31:69:@11175.4]
  assign _T_31025 = valid_34_36 ? 6'h24 : _T_31024; // @[Mux.scala 31:69:@11176.4]
  assign _T_31026 = valid_34_35 ? 6'h23 : _T_31025; // @[Mux.scala 31:69:@11177.4]
  assign _T_31027 = valid_34_34 ? 6'h22 : _T_31026; // @[Mux.scala 31:69:@11178.4]
  assign _T_31028 = valid_34_33 ? 6'h21 : _T_31027; // @[Mux.scala 31:69:@11179.4]
  assign _T_31029 = valid_34_32 ? 6'h20 : _T_31028; // @[Mux.scala 31:69:@11180.4]
  assign _T_31030 = valid_34_31 ? 6'h1f : _T_31029; // @[Mux.scala 31:69:@11181.4]
  assign _T_31031 = valid_34_30 ? 6'h1e : _T_31030; // @[Mux.scala 31:69:@11182.4]
  assign _T_31032 = valid_34_29 ? 6'h1d : _T_31031; // @[Mux.scala 31:69:@11183.4]
  assign _T_31033 = valid_34_28 ? 6'h1c : _T_31032; // @[Mux.scala 31:69:@11184.4]
  assign _T_31034 = valid_34_27 ? 6'h1b : _T_31033; // @[Mux.scala 31:69:@11185.4]
  assign _T_31035 = valid_34_26 ? 6'h1a : _T_31034; // @[Mux.scala 31:69:@11186.4]
  assign _T_31036 = valid_34_25 ? 6'h19 : _T_31035; // @[Mux.scala 31:69:@11187.4]
  assign _T_31037 = valid_34_24 ? 6'h18 : _T_31036; // @[Mux.scala 31:69:@11188.4]
  assign _T_31038 = valid_34_23 ? 6'h17 : _T_31037; // @[Mux.scala 31:69:@11189.4]
  assign _T_31039 = valid_34_22 ? 6'h16 : _T_31038; // @[Mux.scala 31:69:@11190.4]
  assign _T_31040 = valid_34_21 ? 6'h15 : _T_31039; // @[Mux.scala 31:69:@11191.4]
  assign _T_31041 = valid_34_20 ? 6'h14 : _T_31040; // @[Mux.scala 31:69:@11192.4]
  assign _T_31042 = valid_34_19 ? 6'h13 : _T_31041; // @[Mux.scala 31:69:@11193.4]
  assign _T_31043 = valid_34_18 ? 6'h12 : _T_31042; // @[Mux.scala 31:69:@11194.4]
  assign _T_31044 = valid_34_17 ? 6'h11 : _T_31043; // @[Mux.scala 31:69:@11195.4]
  assign _T_31045 = valid_34_16 ? 6'h10 : _T_31044; // @[Mux.scala 31:69:@11196.4]
  assign _T_31046 = valid_34_15 ? 6'hf : _T_31045; // @[Mux.scala 31:69:@11197.4]
  assign _T_31047 = valid_34_14 ? 6'he : _T_31046; // @[Mux.scala 31:69:@11198.4]
  assign _T_31048 = valid_34_13 ? 6'hd : _T_31047; // @[Mux.scala 31:69:@11199.4]
  assign _T_31049 = valid_34_12 ? 6'hc : _T_31048; // @[Mux.scala 31:69:@11200.4]
  assign _T_31050 = valid_34_11 ? 6'hb : _T_31049; // @[Mux.scala 31:69:@11201.4]
  assign _T_31051 = valid_34_10 ? 6'ha : _T_31050; // @[Mux.scala 31:69:@11202.4]
  assign _T_31052 = valid_34_9 ? 6'h9 : _T_31051; // @[Mux.scala 31:69:@11203.4]
  assign _T_31053 = valid_34_8 ? 6'h8 : _T_31052; // @[Mux.scala 31:69:@11204.4]
  assign _T_31054 = valid_34_7 ? 6'h7 : _T_31053; // @[Mux.scala 31:69:@11205.4]
  assign _T_31055 = valid_34_6 ? 6'h6 : _T_31054; // @[Mux.scala 31:69:@11206.4]
  assign _T_31056 = valid_34_5 ? 6'h5 : _T_31055; // @[Mux.scala 31:69:@11207.4]
  assign _T_31057 = valid_34_4 ? 6'h4 : _T_31056; // @[Mux.scala 31:69:@11208.4]
  assign _T_31058 = valid_34_3 ? 6'h3 : _T_31057; // @[Mux.scala 31:69:@11209.4]
  assign _T_31059 = valid_34_2 ? 6'h2 : _T_31058; // @[Mux.scala 31:69:@11210.4]
  assign _T_31060 = valid_34_1 ? 6'h1 : _T_31059; // @[Mux.scala 31:69:@11211.4]
  assign select_34 = valid_34_0 ? 6'h0 : _T_31060; // @[Mux.scala 31:69:@11212.4]
  assign _GEN_2177 = 6'h1 == select_34 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2178 = 6'h2 == select_34 ? io_inData_2 : _GEN_2177; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2179 = 6'h3 == select_34 ? io_inData_3 : _GEN_2178; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2180 = 6'h4 == select_34 ? io_inData_4 : _GEN_2179; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2181 = 6'h5 == select_34 ? io_inData_5 : _GEN_2180; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2182 = 6'h6 == select_34 ? io_inData_6 : _GEN_2181; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2183 = 6'h7 == select_34 ? io_inData_7 : _GEN_2182; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2184 = 6'h8 == select_34 ? io_inData_8 : _GEN_2183; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2185 = 6'h9 == select_34 ? io_inData_9 : _GEN_2184; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2186 = 6'ha == select_34 ? io_inData_10 : _GEN_2185; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2187 = 6'hb == select_34 ? io_inData_11 : _GEN_2186; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2188 = 6'hc == select_34 ? io_inData_12 : _GEN_2187; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2189 = 6'hd == select_34 ? io_inData_13 : _GEN_2188; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2190 = 6'he == select_34 ? io_inData_14 : _GEN_2189; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2191 = 6'hf == select_34 ? io_inData_15 : _GEN_2190; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2192 = 6'h10 == select_34 ? io_inData_16 : _GEN_2191; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2193 = 6'h11 == select_34 ? io_inData_17 : _GEN_2192; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2194 = 6'h12 == select_34 ? io_inData_18 : _GEN_2193; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2195 = 6'h13 == select_34 ? io_inData_19 : _GEN_2194; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2196 = 6'h14 == select_34 ? io_inData_20 : _GEN_2195; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2197 = 6'h15 == select_34 ? io_inData_21 : _GEN_2196; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2198 = 6'h16 == select_34 ? io_inData_22 : _GEN_2197; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2199 = 6'h17 == select_34 ? io_inData_23 : _GEN_2198; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2200 = 6'h18 == select_34 ? io_inData_24 : _GEN_2199; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2201 = 6'h19 == select_34 ? io_inData_25 : _GEN_2200; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2202 = 6'h1a == select_34 ? io_inData_26 : _GEN_2201; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2203 = 6'h1b == select_34 ? io_inData_27 : _GEN_2202; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2204 = 6'h1c == select_34 ? io_inData_28 : _GEN_2203; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2205 = 6'h1d == select_34 ? io_inData_29 : _GEN_2204; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2206 = 6'h1e == select_34 ? io_inData_30 : _GEN_2205; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2207 = 6'h1f == select_34 ? io_inData_31 : _GEN_2206; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2208 = 6'h20 == select_34 ? io_inData_32 : _GEN_2207; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2209 = 6'h21 == select_34 ? io_inData_33 : _GEN_2208; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2210 = 6'h22 == select_34 ? io_inData_34 : _GEN_2209; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2211 = 6'h23 == select_34 ? io_inData_35 : _GEN_2210; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2212 = 6'h24 == select_34 ? io_inData_36 : _GEN_2211; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2213 = 6'h25 == select_34 ? io_inData_37 : _GEN_2212; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2214 = 6'h26 == select_34 ? io_inData_38 : _GEN_2213; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2215 = 6'h27 == select_34 ? io_inData_39 : _GEN_2214; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2216 = 6'h28 == select_34 ? io_inData_40 : _GEN_2215; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2217 = 6'h29 == select_34 ? io_inData_41 : _GEN_2216; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2218 = 6'h2a == select_34 ? io_inData_42 : _GEN_2217; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2219 = 6'h2b == select_34 ? io_inData_43 : _GEN_2218; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2220 = 6'h2c == select_34 ? io_inData_44 : _GEN_2219; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2221 = 6'h2d == select_34 ? io_inData_45 : _GEN_2220; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2222 = 6'h2e == select_34 ? io_inData_46 : _GEN_2221; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2223 = 6'h2f == select_34 ? io_inData_47 : _GEN_2222; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2224 = 6'h30 == select_34 ? io_inData_48 : _GEN_2223; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2225 = 6'h31 == select_34 ? io_inData_49 : _GEN_2224; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2226 = 6'h32 == select_34 ? io_inData_50 : _GEN_2225; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2227 = 6'h33 == select_34 ? io_inData_51 : _GEN_2226; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2228 = 6'h34 == select_34 ? io_inData_52 : _GEN_2227; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2229 = 6'h35 == select_34 ? io_inData_53 : _GEN_2228; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2230 = 6'h36 == select_34 ? io_inData_54 : _GEN_2229; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2231 = 6'h37 == select_34 ? io_inData_55 : _GEN_2230; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2232 = 6'h38 == select_34 ? io_inData_56 : _GEN_2231; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2233 = 6'h39 == select_34 ? io_inData_57 : _GEN_2232; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2234 = 6'h3a == select_34 ? io_inData_58 : _GEN_2233; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2235 = 6'h3b == select_34 ? io_inData_59 : _GEN_2234; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2236 = 6'h3c == select_34 ? io_inData_60 : _GEN_2235; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2237 = 6'h3d == select_34 ? io_inData_61 : _GEN_2236; // @[Switch.scala 33:19:@11214.4]
  assign _GEN_2238 = 6'h3e == select_34 ? io_inData_62 : _GEN_2237; // @[Switch.scala 33:19:@11214.4]
  assign _T_31069 = {valid_34_7,valid_34_6,valid_34_5,valid_34_4,valid_34_3,valid_34_2,valid_34_1,valid_34_0}; // @[Switch.scala 34:32:@11221.4]
  assign _T_31077 = {valid_34_15,valid_34_14,valid_34_13,valid_34_12,valid_34_11,valid_34_10,valid_34_9,valid_34_8,_T_31069}; // @[Switch.scala 34:32:@11229.4]
  assign _T_31084 = {valid_34_23,valid_34_22,valid_34_21,valid_34_20,valid_34_19,valid_34_18,valid_34_17,valid_34_16}; // @[Switch.scala 34:32:@11236.4]
  assign _T_31093 = {valid_34_31,valid_34_30,valid_34_29,valid_34_28,valid_34_27,valid_34_26,valid_34_25,valid_34_24,_T_31084,_T_31077}; // @[Switch.scala 34:32:@11245.4]
  assign _T_31100 = {valid_34_39,valid_34_38,valid_34_37,valid_34_36,valid_34_35,valid_34_34,valid_34_33,valid_34_32}; // @[Switch.scala 34:32:@11252.4]
  assign _T_31108 = {valid_34_47,valid_34_46,valid_34_45,valid_34_44,valid_34_43,valid_34_42,valid_34_41,valid_34_40,_T_31100}; // @[Switch.scala 34:32:@11260.4]
  assign _T_31115 = {valid_34_55,valid_34_54,valid_34_53,valid_34_52,valid_34_51,valid_34_50,valid_34_49,valid_34_48}; // @[Switch.scala 34:32:@11267.4]
  assign _T_31124 = {valid_34_63,valid_34_62,valid_34_61,valid_34_60,valid_34_59,valid_34_58,valid_34_57,valid_34_56,_T_31115,_T_31108}; // @[Switch.scala 34:32:@11276.4]
  assign _T_31125 = {_T_31124,_T_31093}; // @[Switch.scala 34:32:@11277.4]
  assign _T_31129 = io_inAddr_0 == 6'h23; // @[Switch.scala 30:53:@11280.4]
  assign valid_35_0 = io_inValid_0 & _T_31129; // @[Switch.scala 30:36:@11281.4]
  assign _T_31132 = io_inAddr_1 == 6'h23; // @[Switch.scala 30:53:@11283.4]
  assign valid_35_1 = io_inValid_1 & _T_31132; // @[Switch.scala 30:36:@11284.4]
  assign _T_31135 = io_inAddr_2 == 6'h23; // @[Switch.scala 30:53:@11286.4]
  assign valid_35_2 = io_inValid_2 & _T_31135; // @[Switch.scala 30:36:@11287.4]
  assign _T_31138 = io_inAddr_3 == 6'h23; // @[Switch.scala 30:53:@11289.4]
  assign valid_35_3 = io_inValid_3 & _T_31138; // @[Switch.scala 30:36:@11290.4]
  assign _T_31141 = io_inAddr_4 == 6'h23; // @[Switch.scala 30:53:@11292.4]
  assign valid_35_4 = io_inValid_4 & _T_31141; // @[Switch.scala 30:36:@11293.4]
  assign _T_31144 = io_inAddr_5 == 6'h23; // @[Switch.scala 30:53:@11295.4]
  assign valid_35_5 = io_inValid_5 & _T_31144; // @[Switch.scala 30:36:@11296.4]
  assign _T_31147 = io_inAddr_6 == 6'h23; // @[Switch.scala 30:53:@11298.4]
  assign valid_35_6 = io_inValid_6 & _T_31147; // @[Switch.scala 30:36:@11299.4]
  assign _T_31150 = io_inAddr_7 == 6'h23; // @[Switch.scala 30:53:@11301.4]
  assign valid_35_7 = io_inValid_7 & _T_31150; // @[Switch.scala 30:36:@11302.4]
  assign _T_31153 = io_inAddr_8 == 6'h23; // @[Switch.scala 30:53:@11304.4]
  assign valid_35_8 = io_inValid_8 & _T_31153; // @[Switch.scala 30:36:@11305.4]
  assign _T_31156 = io_inAddr_9 == 6'h23; // @[Switch.scala 30:53:@11307.4]
  assign valid_35_9 = io_inValid_9 & _T_31156; // @[Switch.scala 30:36:@11308.4]
  assign _T_31159 = io_inAddr_10 == 6'h23; // @[Switch.scala 30:53:@11310.4]
  assign valid_35_10 = io_inValid_10 & _T_31159; // @[Switch.scala 30:36:@11311.4]
  assign _T_31162 = io_inAddr_11 == 6'h23; // @[Switch.scala 30:53:@11313.4]
  assign valid_35_11 = io_inValid_11 & _T_31162; // @[Switch.scala 30:36:@11314.4]
  assign _T_31165 = io_inAddr_12 == 6'h23; // @[Switch.scala 30:53:@11316.4]
  assign valid_35_12 = io_inValid_12 & _T_31165; // @[Switch.scala 30:36:@11317.4]
  assign _T_31168 = io_inAddr_13 == 6'h23; // @[Switch.scala 30:53:@11319.4]
  assign valid_35_13 = io_inValid_13 & _T_31168; // @[Switch.scala 30:36:@11320.4]
  assign _T_31171 = io_inAddr_14 == 6'h23; // @[Switch.scala 30:53:@11322.4]
  assign valid_35_14 = io_inValid_14 & _T_31171; // @[Switch.scala 30:36:@11323.4]
  assign _T_31174 = io_inAddr_15 == 6'h23; // @[Switch.scala 30:53:@11325.4]
  assign valid_35_15 = io_inValid_15 & _T_31174; // @[Switch.scala 30:36:@11326.4]
  assign _T_31177 = io_inAddr_16 == 6'h23; // @[Switch.scala 30:53:@11328.4]
  assign valid_35_16 = io_inValid_16 & _T_31177; // @[Switch.scala 30:36:@11329.4]
  assign _T_31180 = io_inAddr_17 == 6'h23; // @[Switch.scala 30:53:@11331.4]
  assign valid_35_17 = io_inValid_17 & _T_31180; // @[Switch.scala 30:36:@11332.4]
  assign _T_31183 = io_inAddr_18 == 6'h23; // @[Switch.scala 30:53:@11334.4]
  assign valid_35_18 = io_inValid_18 & _T_31183; // @[Switch.scala 30:36:@11335.4]
  assign _T_31186 = io_inAddr_19 == 6'h23; // @[Switch.scala 30:53:@11337.4]
  assign valid_35_19 = io_inValid_19 & _T_31186; // @[Switch.scala 30:36:@11338.4]
  assign _T_31189 = io_inAddr_20 == 6'h23; // @[Switch.scala 30:53:@11340.4]
  assign valid_35_20 = io_inValid_20 & _T_31189; // @[Switch.scala 30:36:@11341.4]
  assign _T_31192 = io_inAddr_21 == 6'h23; // @[Switch.scala 30:53:@11343.4]
  assign valid_35_21 = io_inValid_21 & _T_31192; // @[Switch.scala 30:36:@11344.4]
  assign _T_31195 = io_inAddr_22 == 6'h23; // @[Switch.scala 30:53:@11346.4]
  assign valid_35_22 = io_inValid_22 & _T_31195; // @[Switch.scala 30:36:@11347.4]
  assign _T_31198 = io_inAddr_23 == 6'h23; // @[Switch.scala 30:53:@11349.4]
  assign valid_35_23 = io_inValid_23 & _T_31198; // @[Switch.scala 30:36:@11350.4]
  assign _T_31201 = io_inAddr_24 == 6'h23; // @[Switch.scala 30:53:@11352.4]
  assign valid_35_24 = io_inValid_24 & _T_31201; // @[Switch.scala 30:36:@11353.4]
  assign _T_31204 = io_inAddr_25 == 6'h23; // @[Switch.scala 30:53:@11355.4]
  assign valid_35_25 = io_inValid_25 & _T_31204; // @[Switch.scala 30:36:@11356.4]
  assign _T_31207 = io_inAddr_26 == 6'h23; // @[Switch.scala 30:53:@11358.4]
  assign valid_35_26 = io_inValid_26 & _T_31207; // @[Switch.scala 30:36:@11359.4]
  assign _T_31210 = io_inAddr_27 == 6'h23; // @[Switch.scala 30:53:@11361.4]
  assign valid_35_27 = io_inValid_27 & _T_31210; // @[Switch.scala 30:36:@11362.4]
  assign _T_31213 = io_inAddr_28 == 6'h23; // @[Switch.scala 30:53:@11364.4]
  assign valid_35_28 = io_inValid_28 & _T_31213; // @[Switch.scala 30:36:@11365.4]
  assign _T_31216 = io_inAddr_29 == 6'h23; // @[Switch.scala 30:53:@11367.4]
  assign valid_35_29 = io_inValid_29 & _T_31216; // @[Switch.scala 30:36:@11368.4]
  assign _T_31219 = io_inAddr_30 == 6'h23; // @[Switch.scala 30:53:@11370.4]
  assign valid_35_30 = io_inValid_30 & _T_31219; // @[Switch.scala 30:36:@11371.4]
  assign _T_31222 = io_inAddr_31 == 6'h23; // @[Switch.scala 30:53:@11373.4]
  assign valid_35_31 = io_inValid_31 & _T_31222; // @[Switch.scala 30:36:@11374.4]
  assign _T_31225 = io_inAddr_32 == 6'h23; // @[Switch.scala 30:53:@11376.4]
  assign valid_35_32 = io_inValid_32 & _T_31225; // @[Switch.scala 30:36:@11377.4]
  assign _T_31228 = io_inAddr_33 == 6'h23; // @[Switch.scala 30:53:@11379.4]
  assign valid_35_33 = io_inValid_33 & _T_31228; // @[Switch.scala 30:36:@11380.4]
  assign _T_31231 = io_inAddr_34 == 6'h23; // @[Switch.scala 30:53:@11382.4]
  assign valid_35_34 = io_inValid_34 & _T_31231; // @[Switch.scala 30:36:@11383.4]
  assign _T_31234 = io_inAddr_35 == 6'h23; // @[Switch.scala 30:53:@11385.4]
  assign valid_35_35 = io_inValid_35 & _T_31234; // @[Switch.scala 30:36:@11386.4]
  assign _T_31237 = io_inAddr_36 == 6'h23; // @[Switch.scala 30:53:@11388.4]
  assign valid_35_36 = io_inValid_36 & _T_31237; // @[Switch.scala 30:36:@11389.4]
  assign _T_31240 = io_inAddr_37 == 6'h23; // @[Switch.scala 30:53:@11391.4]
  assign valid_35_37 = io_inValid_37 & _T_31240; // @[Switch.scala 30:36:@11392.4]
  assign _T_31243 = io_inAddr_38 == 6'h23; // @[Switch.scala 30:53:@11394.4]
  assign valid_35_38 = io_inValid_38 & _T_31243; // @[Switch.scala 30:36:@11395.4]
  assign _T_31246 = io_inAddr_39 == 6'h23; // @[Switch.scala 30:53:@11397.4]
  assign valid_35_39 = io_inValid_39 & _T_31246; // @[Switch.scala 30:36:@11398.4]
  assign _T_31249 = io_inAddr_40 == 6'h23; // @[Switch.scala 30:53:@11400.4]
  assign valid_35_40 = io_inValid_40 & _T_31249; // @[Switch.scala 30:36:@11401.4]
  assign _T_31252 = io_inAddr_41 == 6'h23; // @[Switch.scala 30:53:@11403.4]
  assign valid_35_41 = io_inValid_41 & _T_31252; // @[Switch.scala 30:36:@11404.4]
  assign _T_31255 = io_inAddr_42 == 6'h23; // @[Switch.scala 30:53:@11406.4]
  assign valid_35_42 = io_inValid_42 & _T_31255; // @[Switch.scala 30:36:@11407.4]
  assign _T_31258 = io_inAddr_43 == 6'h23; // @[Switch.scala 30:53:@11409.4]
  assign valid_35_43 = io_inValid_43 & _T_31258; // @[Switch.scala 30:36:@11410.4]
  assign _T_31261 = io_inAddr_44 == 6'h23; // @[Switch.scala 30:53:@11412.4]
  assign valid_35_44 = io_inValid_44 & _T_31261; // @[Switch.scala 30:36:@11413.4]
  assign _T_31264 = io_inAddr_45 == 6'h23; // @[Switch.scala 30:53:@11415.4]
  assign valid_35_45 = io_inValid_45 & _T_31264; // @[Switch.scala 30:36:@11416.4]
  assign _T_31267 = io_inAddr_46 == 6'h23; // @[Switch.scala 30:53:@11418.4]
  assign valid_35_46 = io_inValid_46 & _T_31267; // @[Switch.scala 30:36:@11419.4]
  assign _T_31270 = io_inAddr_47 == 6'h23; // @[Switch.scala 30:53:@11421.4]
  assign valid_35_47 = io_inValid_47 & _T_31270; // @[Switch.scala 30:36:@11422.4]
  assign _T_31273 = io_inAddr_48 == 6'h23; // @[Switch.scala 30:53:@11424.4]
  assign valid_35_48 = io_inValid_48 & _T_31273; // @[Switch.scala 30:36:@11425.4]
  assign _T_31276 = io_inAddr_49 == 6'h23; // @[Switch.scala 30:53:@11427.4]
  assign valid_35_49 = io_inValid_49 & _T_31276; // @[Switch.scala 30:36:@11428.4]
  assign _T_31279 = io_inAddr_50 == 6'h23; // @[Switch.scala 30:53:@11430.4]
  assign valid_35_50 = io_inValid_50 & _T_31279; // @[Switch.scala 30:36:@11431.4]
  assign _T_31282 = io_inAddr_51 == 6'h23; // @[Switch.scala 30:53:@11433.4]
  assign valid_35_51 = io_inValid_51 & _T_31282; // @[Switch.scala 30:36:@11434.4]
  assign _T_31285 = io_inAddr_52 == 6'h23; // @[Switch.scala 30:53:@11436.4]
  assign valid_35_52 = io_inValid_52 & _T_31285; // @[Switch.scala 30:36:@11437.4]
  assign _T_31288 = io_inAddr_53 == 6'h23; // @[Switch.scala 30:53:@11439.4]
  assign valid_35_53 = io_inValid_53 & _T_31288; // @[Switch.scala 30:36:@11440.4]
  assign _T_31291 = io_inAddr_54 == 6'h23; // @[Switch.scala 30:53:@11442.4]
  assign valid_35_54 = io_inValid_54 & _T_31291; // @[Switch.scala 30:36:@11443.4]
  assign _T_31294 = io_inAddr_55 == 6'h23; // @[Switch.scala 30:53:@11445.4]
  assign valid_35_55 = io_inValid_55 & _T_31294; // @[Switch.scala 30:36:@11446.4]
  assign _T_31297 = io_inAddr_56 == 6'h23; // @[Switch.scala 30:53:@11448.4]
  assign valid_35_56 = io_inValid_56 & _T_31297; // @[Switch.scala 30:36:@11449.4]
  assign _T_31300 = io_inAddr_57 == 6'h23; // @[Switch.scala 30:53:@11451.4]
  assign valid_35_57 = io_inValid_57 & _T_31300; // @[Switch.scala 30:36:@11452.4]
  assign _T_31303 = io_inAddr_58 == 6'h23; // @[Switch.scala 30:53:@11454.4]
  assign valid_35_58 = io_inValid_58 & _T_31303; // @[Switch.scala 30:36:@11455.4]
  assign _T_31306 = io_inAddr_59 == 6'h23; // @[Switch.scala 30:53:@11457.4]
  assign valid_35_59 = io_inValid_59 & _T_31306; // @[Switch.scala 30:36:@11458.4]
  assign _T_31309 = io_inAddr_60 == 6'h23; // @[Switch.scala 30:53:@11460.4]
  assign valid_35_60 = io_inValid_60 & _T_31309; // @[Switch.scala 30:36:@11461.4]
  assign _T_31312 = io_inAddr_61 == 6'h23; // @[Switch.scala 30:53:@11463.4]
  assign valid_35_61 = io_inValid_61 & _T_31312; // @[Switch.scala 30:36:@11464.4]
  assign _T_31315 = io_inAddr_62 == 6'h23; // @[Switch.scala 30:53:@11466.4]
  assign valid_35_62 = io_inValid_62 & _T_31315; // @[Switch.scala 30:36:@11467.4]
  assign _T_31318 = io_inAddr_63 == 6'h23; // @[Switch.scala 30:53:@11469.4]
  assign valid_35_63 = io_inValid_63 & _T_31318; // @[Switch.scala 30:36:@11470.4]
  assign _T_31384 = valid_35_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@11472.4]
  assign _T_31385 = valid_35_61 ? 6'h3d : _T_31384; // @[Mux.scala 31:69:@11473.4]
  assign _T_31386 = valid_35_60 ? 6'h3c : _T_31385; // @[Mux.scala 31:69:@11474.4]
  assign _T_31387 = valid_35_59 ? 6'h3b : _T_31386; // @[Mux.scala 31:69:@11475.4]
  assign _T_31388 = valid_35_58 ? 6'h3a : _T_31387; // @[Mux.scala 31:69:@11476.4]
  assign _T_31389 = valid_35_57 ? 6'h39 : _T_31388; // @[Mux.scala 31:69:@11477.4]
  assign _T_31390 = valid_35_56 ? 6'h38 : _T_31389; // @[Mux.scala 31:69:@11478.4]
  assign _T_31391 = valid_35_55 ? 6'h37 : _T_31390; // @[Mux.scala 31:69:@11479.4]
  assign _T_31392 = valid_35_54 ? 6'h36 : _T_31391; // @[Mux.scala 31:69:@11480.4]
  assign _T_31393 = valid_35_53 ? 6'h35 : _T_31392; // @[Mux.scala 31:69:@11481.4]
  assign _T_31394 = valid_35_52 ? 6'h34 : _T_31393; // @[Mux.scala 31:69:@11482.4]
  assign _T_31395 = valid_35_51 ? 6'h33 : _T_31394; // @[Mux.scala 31:69:@11483.4]
  assign _T_31396 = valid_35_50 ? 6'h32 : _T_31395; // @[Mux.scala 31:69:@11484.4]
  assign _T_31397 = valid_35_49 ? 6'h31 : _T_31396; // @[Mux.scala 31:69:@11485.4]
  assign _T_31398 = valid_35_48 ? 6'h30 : _T_31397; // @[Mux.scala 31:69:@11486.4]
  assign _T_31399 = valid_35_47 ? 6'h2f : _T_31398; // @[Mux.scala 31:69:@11487.4]
  assign _T_31400 = valid_35_46 ? 6'h2e : _T_31399; // @[Mux.scala 31:69:@11488.4]
  assign _T_31401 = valid_35_45 ? 6'h2d : _T_31400; // @[Mux.scala 31:69:@11489.4]
  assign _T_31402 = valid_35_44 ? 6'h2c : _T_31401; // @[Mux.scala 31:69:@11490.4]
  assign _T_31403 = valid_35_43 ? 6'h2b : _T_31402; // @[Mux.scala 31:69:@11491.4]
  assign _T_31404 = valid_35_42 ? 6'h2a : _T_31403; // @[Mux.scala 31:69:@11492.4]
  assign _T_31405 = valid_35_41 ? 6'h29 : _T_31404; // @[Mux.scala 31:69:@11493.4]
  assign _T_31406 = valid_35_40 ? 6'h28 : _T_31405; // @[Mux.scala 31:69:@11494.4]
  assign _T_31407 = valid_35_39 ? 6'h27 : _T_31406; // @[Mux.scala 31:69:@11495.4]
  assign _T_31408 = valid_35_38 ? 6'h26 : _T_31407; // @[Mux.scala 31:69:@11496.4]
  assign _T_31409 = valid_35_37 ? 6'h25 : _T_31408; // @[Mux.scala 31:69:@11497.4]
  assign _T_31410 = valid_35_36 ? 6'h24 : _T_31409; // @[Mux.scala 31:69:@11498.4]
  assign _T_31411 = valid_35_35 ? 6'h23 : _T_31410; // @[Mux.scala 31:69:@11499.4]
  assign _T_31412 = valid_35_34 ? 6'h22 : _T_31411; // @[Mux.scala 31:69:@11500.4]
  assign _T_31413 = valid_35_33 ? 6'h21 : _T_31412; // @[Mux.scala 31:69:@11501.4]
  assign _T_31414 = valid_35_32 ? 6'h20 : _T_31413; // @[Mux.scala 31:69:@11502.4]
  assign _T_31415 = valid_35_31 ? 6'h1f : _T_31414; // @[Mux.scala 31:69:@11503.4]
  assign _T_31416 = valid_35_30 ? 6'h1e : _T_31415; // @[Mux.scala 31:69:@11504.4]
  assign _T_31417 = valid_35_29 ? 6'h1d : _T_31416; // @[Mux.scala 31:69:@11505.4]
  assign _T_31418 = valid_35_28 ? 6'h1c : _T_31417; // @[Mux.scala 31:69:@11506.4]
  assign _T_31419 = valid_35_27 ? 6'h1b : _T_31418; // @[Mux.scala 31:69:@11507.4]
  assign _T_31420 = valid_35_26 ? 6'h1a : _T_31419; // @[Mux.scala 31:69:@11508.4]
  assign _T_31421 = valid_35_25 ? 6'h19 : _T_31420; // @[Mux.scala 31:69:@11509.4]
  assign _T_31422 = valid_35_24 ? 6'h18 : _T_31421; // @[Mux.scala 31:69:@11510.4]
  assign _T_31423 = valid_35_23 ? 6'h17 : _T_31422; // @[Mux.scala 31:69:@11511.4]
  assign _T_31424 = valid_35_22 ? 6'h16 : _T_31423; // @[Mux.scala 31:69:@11512.4]
  assign _T_31425 = valid_35_21 ? 6'h15 : _T_31424; // @[Mux.scala 31:69:@11513.4]
  assign _T_31426 = valid_35_20 ? 6'h14 : _T_31425; // @[Mux.scala 31:69:@11514.4]
  assign _T_31427 = valid_35_19 ? 6'h13 : _T_31426; // @[Mux.scala 31:69:@11515.4]
  assign _T_31428 = valid_35_18 ? 6'h12 : _T_31427; // @[Mux.scala 31:69:@11516.4]
  assign _T_31429 = valid_35_17 ? 6'h11 : _T_31428; // @[Mux.scala 31:69:@11517.4]
  assign _T_31430 = valid_35_16 ? 6'h10 : _T_31429; // @[Mux.scala 31:69:@11518.4]
  assign _T_31431 = valid_35_15 ? 6'hf : _T_31430; // @[Mux.scala 31:69:@11519.4]
  assign _T_31432 = valid_35_14 ? 6'he : _T_31431; // @[Mux.scala 31:69:@11520.4]
  assign _T_31433 = valid_35_13 ? 6'hd : _T_31432; // @[Mux.scala 31:69:@11521.4]
  assign _T_31434 = valid_35_12 ? 6'hc : _T_31433; // @[Mux.scala 31:69:@11522.4]
  assign _T_31435 = valid_35_11 ? 6'hb : _T_31434; // @[Mux.scala 31:69:@11523.4]
  assign _T_31436 = valid_35_10 ? 6'ha : _T_31435; // @[Mux.scala 31:69:@11524.4]
  assign _T_31437 = valid_35_9 ? 6'h9 : _T_31436; // @[Mux.scala 31:69:@11525.4]
  assign _T_31438 = valid_35_8 ? 6'h8 : _T_31437; // @[Mux.scala 31:69:@11526.4]
  assign _T_31439 = valid_35_7 ? 6'h7 : _T_31438; // @[Mux.scala 31:69:@11527.4]
  assign _T_31440 = valid_35_6 ? 6'h6 : _T_31439; // @[Mux.scala 31:69:@11528.4]
  assign _T_31441 = valid_35_5 ? 6'h5 : _T_31440; // @[Mux.scala 31:69:@11529.4]
  assign _T_31442 = valid_35_4 ? 6'h4 : _T_31441; // @[Mux.scala 31:69:@11530.4]
  assign _T_31443 = valid_35_3 ? 6'h3 : _T_31442; // @[Mux.scala 31:69:@11531.4]
  assign _T_31444 = valid_35_2 ? 6'h2 : _T_31443; // @[Mux.scala 31:69:@11532.4]
  assign _T_31445 = valid_35_1 ? 6'h1 : _T_31444; // @[Mux.scala 31:69:@11533.4]
  assign select_35 = valid_35_0 ? 6'h0 : _T_31445; // @[Mux.scala 31:69:@11534.4]
  assign _GEN_2241 = 6'h1 == select_35 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2242 = 6'h2 == select_35 ? io_inData_2 : _GEN_2241; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2243 = 6'h3 == select_35 ? io_inData_3 : _GEN_2242; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2244 = 6'h4 == select_35 ? io_inData_4 : _GEN_2243; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2245 = 6'h5 == select_35 ? io_inData_5 : _GEN_2244; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2246 = 6'h6 == select_35 ? io_inData_6 : _GEN_2245; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2247 = 6'h7 == select_35 ? io_inData_7 : _GEN_2246; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2248 = 6'h8 == select_35 ? io_inData_8 : _GEN_2247; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2249 = 6'h9 == select_35 ? io_inData_9 : _GEN_2248; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2250 = 6'ha == select_35 ? io_inData_10 : _GEN_2249; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2251 = 6'hb == select_35 ? io_inData_11 : _GEN_2250; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2252 = 6'hc == select_35 ? io_inData_12 : _GEN_2251; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2253 = 6'hd == select_35 ? io_inData_13 : _GEN_2252; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2254 = 6'he == select_35 ? io_inData_14 : _GEN_2253; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2255 = 6'hf == select_35 ? io_inData_15 : _GEN_2254; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2256 = 6'h10 == select_35 ? io_inData_16 : _GEN_2255; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2257 = 6'h11 == select_35 ? io_inData_17 : _GEN_2256; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2258 = 6'h12 == select_35 ? io_inData_18 : _GEN_2257; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2259 = 6'h13 == select_35 ? io_inData_19 : _GEN_2258; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2260 = 6'h14 == select_35 ? io_inData_20 : _GEN_2259; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2261 = 6'h15 == select_35 ? io_inData_21 : _GEN_2260; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2262 = 6'h16 == select_35 ? io_inData_22 : _GEN_2261; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2263 = 6'h17 == select_35 ? io_inData_23 : _GEN_2262; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2264 = 6'h18 == select_35 ? io_inData_24 : _GEN_2263; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2265 = 6'h19 == select_35 ? io_inData_25 : _GEN_2264; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2266 = 6'h1a == select_35 ? io_inData_26 : _GEN_2265; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2267 = 6'h1b == select_35 ? io_inData_27 : _GEN_2266; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2268 = 6'h1c == select_35 ? io_inData_28 : _GEN_2267; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2269 = 6'h1d == select_35 ? io_inData_29 : _GEN_2268; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2270 = 6'h1e == select_35 ? io_inData_30 : _GEN_2269; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2271 = 6'h1f == select_35 ? io_inData_31 : _GEN_2270; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2272 = 6'h20 == select_35 ? io_inData_32 : _GEN_2271; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2273 = 6'h21 == select_35 ? io_inData_33 : _GEN_2272; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2274 = 6'h22 == select_35 ? io_inData_34 : _GEN_2273; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2275 = 6'h23 == select_35 ? io_inData_35 : _GEN_2274; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2276 = 6'h24 == select_35 ? io_inData_36 : _GEN_2275; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2277 = 6'h25 == select_35 ? io_inData_37 : _GEN_2276; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2278 = 6'h26 == select_35 ? io_inData_38 : _GEN_2277; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2279 = 6'h27 == select_35 ? io_inData_39 : _GEN_2278; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2280 = 6'h28 == select_35 ? io_inData_40 : _GEN_2279; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2281 = 6'h29 == select_35 ? io_inData_41 : _GEN_2280; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2282 = 6'h2a == select_35 ? io_inData_42 : _GEN_2281; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2283 = 6'h2b == select_35 ? io_inData_43 : _GEN_2282; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2284 = 6'h2c == select_35 ? io_inData_44 : _GEN_2283; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2285 = 6'h2d == select_35 ? io_inData_45 : _GEN_2284; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2286 = 6'h2e == select_35 ? io_inData_46 : _GEN_2285; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2287 = 6'h2f == select_35 ? io_inData_47 : _GEN_2286; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2288 = 6'h30 == select_35 ? io_inData_48 : _GEN_2287; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2289 = 6'h31 == select_35 ? io_inData_49 : _GEN_2288; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2290 = 6'h32 == select_35 ? io_inData_50 : _GEN_2289; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2291 = 6'h33 == select_35 ? io_inData_51 : _GEN_2290; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2292 = 6'h34 == select_35 ? io_inData_52 : _GEN_2291; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2293 = 6'h35 == select_35 ? io_inData_53 : _GEN_2292; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2294 = 6'h36 == select_35 ? io_inData_54 : _GEN_2293; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2295 = 6'h37 == select_35 ? io_inData_55 : _GEN_2294; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2296 = 6'h38 == select_35 ? io_inData_56 : _GEN_2295; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2297 = 6'h39 == select_35 ? io_inData_57 : _GEN_2296; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2298 = 6'h3a == select_35 ? io_inData_58 : _GEN_2297; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2299 = 6'h3b == select_35 ? io_inData_59 : _GEN_2298; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2300 = 6'h3c == select_35 ? io_inData_60 : _GEN_2299; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2301 = 6'h3d == select_35 ? io_inData_61 : _GEN_2300; // @[Switch.scala 33:19:@11536.4]
  assign _GEN_2302 = 6'h3e == select_35 ? io_inData_62 : _GEN_2301; // @[Switch.scala 33:19:@11536.4]
  assign _T_31454 = {valid_35_7,valid_35_6,valid_35_5,valid_35_4,valid_35_3,valid_35_2,valid_35_1,valid_35_0}; // @[Switch.scala 34:32:@11543.4]
  assign _T_31462 = {valid_35_15,valid_35_14,valid_35_13,valid_35_12,valid_35_11,valid_35_10,valid_35_9,valid_35_8,_T_31454}; // @[Switch.scala 34:32:@11551.4]
  assign _T_31469 = {valid_35_23,valid_35_22,valid_35_21,valid_35_20,valid_35_19,valid_35_18,valid_35_17,valid_35_16}; // @[Switch.scala 34:32:@11558.4]
  assign _T_31478 = {valid_35_31,valid_35_30,valid_35_29,valid_35_28,valid_35_27,valid_35_26,valid_35_25,valid_35_24,_T_31469,_T_31462}; // @[Switch.scala 34:32:@11567.4]
  assign _T_31485 = {valid_35_39,valid_35_38,valid_35_37,valid_35_36,valid_35_35,valid_35_34,valid_35_33,valid_35_32}; // @[Switch.scala 34:32:@11574.4]
  assign _T_31493 = {valid_35_47,valid_35_46,valid_35_45,valid_35_44,valid_35_43,valid_35_42,valid_35_41,valid_35_40,_T_31485}; // @[Switch.scala 34:32:@11582.4]
  assign _T_31500 = {valid_35_55,valid_35_54,valid_35_53,valid_35_52,valid_35_51,valid_35_50,valid_35_49,valid_35_48}; // @[Switch.scala 34:32:@11589.4]
  assign _T_31509 = {valid_35_63,valid_35_62,valid_35_61,valid_35_60,valid_35_59,valid_35_58,valid_35_57,valid_35_56,_T_31500,_T_31493}; // @[Switch.scala 34:32:@11598.4]
  assign _T_31510 = {_T_31509,_T_31478}; // @[Switch.scala 34:32:@11599.4]
  assign _T_31514 = io_inAddr_0 == 6'h24; // @[Switch.scala 30:53:@11602.4]
  assign valid_36_0 = io_inValid_0 & _T_31514; // @[Switch.scala 30:36:@11603.4]
  assign _T_31517 = io_inAddr_1 == 6'h24; // @[Switch.scala 30:53:@11605.4]
  assign valid_36_1 = io_inValid_1 & _T_31517; // @[Switch.scala 30:36:@11606.4]
  assign _T_31520 = io_inAddr_2 == 6'h24; // @[Switch.scala 30:53:@11608.4]
  assign valid_36_2 = io_inValid_2 & _T_31520; // @[Switch.scala 30:36:@11609.4]
  assign _T_31523 = io_inAddr_3 == 6'h24; // @[Switch.scala 30:53:@11611.4]
  assign valid_36_3 = io_inValid_3 & _T_31523; // @[Switch.scala 30:36:@11612.4]
  assign _T_31526 = io_inAddr_4 == 6'h24; // @[Switch.scala 30:53:@11614.4]
  assign valid_36_4 = io_inValid_4 & _T_31526; // @[Switch.scala 30:36:@11615.4]
  assign _T_31529 = io_inAddr_5 == 6'h24; // @[Switch.scala 30:53:@11617.4]
  assign valid_36_5 = io_inValid_5 & _T_31529; // @[Switch.scala 30:36:@11618.4]
  assign _T_31532 = io_inAddr_6 == 6'h24; // @[Switch.scala 30:53:@11620.4]
  assign valid_36_6 = io_inValid_6 & _T_31532; // @[Switch.scala 30:36:@11621.4]
  assign _T_31535 = io_inAddr_7 == 6'h24; // @[Switch.scala 30:53:@11623.4]
  assign valid_36_7 = io_inValid_7 & _T_31535; // @[Switch.scala 30:36:@11624.4]
  assign _T_31538 = io_inAddr_8 == 6'h24; // @[Switch.scala 30:53:@11626.4]
  assign valid_36_8 = io_inValid_8 & _T_31538; // @[Switch.scala 30:36:@11627.4]
  assign _T_31541 = io_inAddr_9 == 6'h24; // @[Switch.scala 30:53:@11629.4]
  assign valid_36_9 = io_inValid_9 & _T_31541; // @[Switch.scala 30:36:@11630.4]
  assign _T_31544 = io_inAddr_10 == 6'h24; // @[Switch.scala 30:53:@11632.4]
  assign valid_36_10 = io_inValid_10 & _T_31544; // @[Switch.scala 30:36:@11633.4]
  assign _T_31547 = io_inAddr_11 == 6'h24; // @[Switch.scala 30:53:@11635.4]
  assign valid_36_11 = io_inValid_11 & _T_31547; // @[Switch.scala 30:36:@11636.4]
  assign _T_31550 = io_inAddr_12 == 6'h24; // @[Switch.scala 30:53:@11638.4]
  assign valid_36_12 = io_inValid_12 & _T_31550; // @[Switch.scala 30:36:@11639.4]
  assign _T_31553 = io_inAddr_13 == 6'h24; // @[Switch.scala 30:53:@11641.4]
  assign valid_36_13 = io_inValid_13 & _T_31553; // @[Switch.scala 30:36:@11642.4]
  assign _T_31556 = io_inAddr_14 == 6'h24; // @[Switch.scala 30:53:@11644.4]
  assign valid_36_14 = io_inValid_14 & _T_31556; // @[Switch.scala 30:36:@11645.4]
  assign _T_31559 = io_inAddr_15 == 6'h24; // @[Switch.scala 30:53:@11647.4]
  assign valid_36_15 = io_inValid_15 & _T_31559; // @[Switch.scala 30:36:@11648.4]
  assign _T_31562 = io_inAddr_16 == 6'h24; // @[Switch.scala 30:53:@11650.4]
  assign valid_36_16 = io_inValid_16 & _T_31562; // @[Switch.scala 30:36:@11651.4]
  assign _T_31565 = io_inAddr_17 == 6'h24; // @[Switch.scala 30:53:@11653.4]
  assign valid_36_17 = io_inValid_17 & _T_31565; // @[Switch.scala 30:36:@11654.4]
  assign _T_31568 = io_inAddr_18 == 6'h24; // @[Switch.scala 30:53:@11656.4]
  assign valid_36_18 = io_inValid_18 & _T_31568; // @[Switch.scala 30:36:@11657.4]
  assign _T_31571 = io_inAddr_19 == 6'h24; // @[Switch.scala 30:53:@11659.4]
  assign valid_36_19 = io_inValid_19 & _T_31571; // @[Switch.scala 30:36:@11660.4]
  assign _T_31574 = io_inAddr_20 == 6'h24; // @[Switch.scala 30:53:@11662.4]
  assign valid_36_20 = io_inValid_20 & _T_31574; // @[Switch.scala 30:36:@11663.4]
  assign _T_31577 = io_inAddr_21 == 6'h24; // @[Switch.scala 30:53:@11665.4]
  assign valid_36_21 = io_inValid_21 & _T_31577; // @[Switch.scala 30:36:@11666.4]
  assign _T_31580 = io_inAddr_22 == 6'h24; // @[Switch.scala 30:53:@11668.4]
  assign valid_36_22 = io_inValid_22 & _T_31580; // @[Switch.scala 30:36:@11669.4]
  assign _T_31583 = io_inAddr_23 == 6'h24; // @[Switch.scala 30:53:@11671.4]
  assign valid_36_23 = io_inValid_23 & _T_31583; // @[Switch.scala 30:36:@11672.4]
  assign _T_31586 = io_inAddr_24 == 6'h24; // @[Switch.scala 30:53:@11674.4]
  assign valid_36_24 = io_inValid_24 & _T_31586; // @[Switch.scala 30:36:@11675.4]
  assign _T_31589 = io_inAddr_25 == 6'h24; // @[Switch.scala 30:53:@11677.4]
  assign valid_36_25 = io_inValid_25 & _T_31589; // @[Switch.scala 30:36:@11678.4]
  assign _T_31592 = io_inAddr_26 == 6'h24; // @[Switch.scala 30:53:@11680.4]
  assign valid_36_26 = io_inValid_26 & _T_31592; // @[Switch.scala 30:36:@11681.4]
  assign _T_31595 = io_inAddr_27 == 6'h24; // @[Switch.scala 30:53:@11683.4]
  assign valid_36_27 = io_inValid_27 & _T_31595; // @[Switch.scala 30:36:@11684.4]
  assign _T_31598 = io_inAddr_28 == 6'h24; // @[Switch.scala 30:53:@11686.4]
  assign valid_36_28 = io_inValid_28 & _T_31598; // @[Switch.scala 30:36:@11687.4]
  assign _T_31601 = io_inAddr_29 == 6'h24; // @[Switch.scala 30:53:@11689.4]
  assign valid_36_29 = io_inValid_29 & _T_31601; // @[Switch.scala 30:36:@11690.4]
  assign _T_31604 = io_inAddr_30 == 6'h24; // @[Switch.scala 30:53:@11692.4]
  assign valid_36_30 = io_inValid_30 & _T_31604; // @[Switch.scala 30:36:@11693.4]
  assign _T_31607 = io_inAddr_31 == 6'h24; // @[Switch.scala 30:53:@11695.4]
  assign valid_36_31 = io_inValid_31 & _T_31607; // @[Switch.scala 30:36:@11696.4]
  assign _T_31610 = io_inAddr_32 == 6'h24; // @[Switch.scala 30:53:@11698.4]
  assign valid_36_32 = io_inValid_32 & _T_31610; // @[Switch.scala 30:36:@11699.4]
  assign _T_31613 = io_inAddr_33 == 6'h24; // @[Switch.scala 30:53:@11701.4]
  assign valid_36_33 = io_inValid_33 & _T_31613; // @[Switch.scala 30:36:@11702.4]
  assign _T_31616 = io_inAddr_34 == 6'h24; // @[Switch.scala 30:53:@11704.4]
  assign valid_36_34 = io_inValid_34 & _T_31616; // @[Switch.scala 30:36:@11705.4]
  assign _T_31619 = io_inAddr_35 == 6'h24; // @[Switch.scala 30:53:@11707.4]
  assign valid_36_35 = io_inValid_35 & _T_31619; // @[Switch.scala 30:36:@11708.4]
  assign _T_31622 = io_inAddr_36 == 6'h24; // @[Switch.scala 30:53:@11710.4]
  assign valid_36_36 = io_inValid_36 & _T_31622; // @[Switch.scala 30:36:@11711.4]
  assign _T_31625 = io_inAddr_37 == 6'h24; // @[Switch.scala 30:53:@11713.4]
  assign valid_36_37 = io_inValid_37 & _T_31625; // @[Switch.scala 30:36:@11714.4]
  assign _T_31628 = io_inAddr_38 == 6'h24; // @[Switch.scala 30:53:@11716.4]
  assign valid_36_38 = io_inValid_38 & _T_31628; // @[Switch.scala 30:36:@11717.4]
  assign _T_31631 = io_inAddr_39 == 6'h24; // @[Switch.scala 30:53:@11719.4]
  assign valid_36_39 = io_inValid_39 & _T_31631; // @[Switch.scala 30:36:@11720.4]
  assign _T_31634 = io_inAddr_40 == 6'h24; // @[Switch.scala 30:53:@11722.4]
  assign valid_36_40 = io_inValid_40 & _T_31634; // @[Switch.scala 30:36:@11723.4]
  assign _T_31637 = io_inAddr_41 == 6'h24; // @[Switch.scala 30:53:@11725.4]
  assign valid_36_41 = io_inValid_41 & _T_31637; // @[Switch.scala 30:36:@11726.4]
  assign _T_31640 = io_inAddr_42 == 6'h24; // @[Switch.scala 30:53:@11728.4]
  assign valid_36_42 = io_inValid_42 & _T_31640; // @[Switch.scala 30:36:@11729.4]
  assign _T_31643 = io_inAddr_43 == 6'h24; // @[Switch.scala 30:53:@11731.4]
  assign valid_36_43 = io_inValid_43 & _T_31643; // @[Switch.scala 30:36:@11732.4]
  assign _T_31646 = io_inAddr_44 == 6'h24; // @[Switch.scala 30:53:@11734.4]
  assign valid_36_44 = io_inValid_44 & _T_31646; // @[Switch.scala 30:36:@11735.4]
  assign _T_31649 = io_inAddr_45 == 6'h24; // @[Switch.scala 30:53:@11737.4]
  assign valid_36_45 = io_inValid_45 & _T_31649; // @[Switch.scala 30:36:@11738.4]
  assign _T_31652 = io_inAddr_46 == 6'h24; // @[Switch.scala 30:53:@11740.4]
  assign valid_36_46 = io_inValid_46 & _T_31652; // @[Switch.scala 30:36:@11741.4]
  assign _T_31655 = io_inAddr_47 == 6'h24; // @[Switch.scala 30:53:@11743.4]
  assign valid_36_47 = io_inValid_47 & _T_31655; // @[Switch.scala 30:36:@11744.4]
  assign _T_31658 = io_inAddr_48 == 6'h24; // @[Switch.scala 30:53:@11746.4]
  assign valid_36_48 = io_inValid_48 & _T_31658; // @[Switch.scala 30:36:@11747.4]
  assign _T_31661 = io_inAddr_49 == 6'h24; // @[Switch.scala 30:53:@11749.4]
  assign valid_36_49 = io_inValid_49 & _T_31661; // @[Switch.scala 30:36:@11750.4]
  assign _T_31664 = io_inAddr_50 == 6'h24; // @[Switch.scala 30:53:@11752.4]
  assign valid_36_50 = io_inValid_50 & _T_31664; // @[Switch.scala 30:36:@11753.4]
  assign _T_31667 = io_inAddr_51 == 6'h24; // @[Switch.scala 30:53:@11755.4]
  assign valid_36_51 = io_inValid_51 & _T_31667; // @[Switch.scala 30:36:@11756.4]
  assign _T_31670 = io_inAddr_52 == 6'h24; // @[Switch.scala 30:53:@11758.4]
  assign valid_36_52 = io_inValid_52 & _T_31670; // @[Switch.scala 30:36:@11759.4]
  assign _T_31673 = io_inAddr_53 == 6'h24; // @[Switch.scala 30:53:@11761.4]
  assign valid_36_53 = io_inValid_53 & _T_31673; // @[Switch.scala 30:36:@11762.4]
  assign _T_31676 = io_inAddr_54 == 6'h24; // @[Switch.scala 30:53:@11764.4]
  assign valid_36_54 = io_inValid_54 & _T_31676; // @[Switch.scala 30:36:@11765.4]
  assign _T_31679 = io_inAddr_55 == 6'h24; // @[Switch.scala 30:53:@11767.4]
  assign valid_36_55 = io_inValid_55 & _T_31679; // @[Switch.scala 30:36:@11768.4]
  assign _T_31682 = io_inAddr_56 == 6'h24; // @[Switch.scala 30:53:@11770.4]
  assign valid_36_56 = io_inValid_56 & _T_31682; // @[Switch.scala 30:36:@11771.4]
  assign _T_31685 = io_inAddr_57 == 6'h24; // @[Switch.scala 30:53:@11773.4]
  assign valid_36_57 = io_inValid_57 & _T_31685; // @[Switch.scala 30:36:@11774.4]
  assign _T_31688 = io_inAddr_58 == 6'h24; // @[Switch.scala 30:53:@11776.4]
  assign valid_36_58 = io_inValid_58 & _T_31688; // @[Switch.scala 30:36:@11777.4]
  assign _T_31691 = io_inAddr_59 == 6'h24; // @[Switch.scala 30:53:@11779.4]
  assign valid_36_59 = io_inValid_59 & _T_31691; // @[Switch.scala 30:36:@11780.4]
  assign _T_31694 = io_inAddr_60 == 6'h24; // @[Switch.scala 30:53:@11782.4]
  assign valid_36_60 = io_inValid_60 & _T_31694; // @[Switch.scala 30:36:@11783.4]
  assign _T_31697 = io_inAddr_61 == 6'h24; // @[Switch.scala 30:53:@11785.4]
  assign valid_36_61 = io_inValid_61 & _T_31697; // @[Switch.scala 30:36:@11786.4]
  assign _T_31700 = io_inAddr_62 == 6'h24; // @[Switch.scala 30:53:@11788.4]
  assign valid_36_62 = io_inValid_62 & _T_31700; // @[Switch.scala 30:36:@11789.4]
  assign _T_31703 = io_inAddr_63 == 6'h24; // @[Switch.scala 30:53:@11791.4]
  assign valid_36_63 = io_inValid_63 & _T_31703; // @[Switch.scala 30:36:@11792.4]
  assign _T_31769 = valid_36_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@11794.4]
  assign _T_31770 = valid_36_61 ? 6'h3d : _T_31769; // @[Mux.scala 31:69:@11795.4]
  assign _T_31771 = valid_36_60 ? 6'h3c : _T_31770; // @[Mux.scala 31:69:@11796.4]
  assign _T_31772 = valid_36_59 ? 6'h3b : _T_31771; // @[Mux.scala 31:69:@11797.4]
  assign _T_31773 = valid_36_58 ? 6'h3a : _T_31772; // @[Mux.scala 31:69:@11798.4]
  assign _T_31774 = valid_36_57 ? 6'h39 : _T_31773; // @[Mux.scala 31:69:@11799.4]
  assign _T_31775 = valid_36_56 ? 6'h38 : _T_31774; // @[Mux.scala 31:69:@11800.4]
  assign _T_31776 = valid_36_55 ? 6'h37 : _T_31775; // @[Mux.scala 31:69:@11801.4]
  assign _T_31777 = valid_36_54 ? 6'h36 : _T_31776; // @[Mux.scala 31:69:@11802.4]
  assign _T_31778 = valid_36_53 ? 6'h35 : _T_31777; // @[Mux.scala 31:69:@11803.4]
  assign _T_31779 = valid_36_52 ? 6'h34 : _T_31778; // @[Mux.scala 31:69:@11804.4]
  assign _T_31780 = valid_36_51 ? 6'h33 : _T_31779; // @[Mux.scala 31:69:@11805.4]
  assign _T_31781 = valid_36_50 ? 6'h32 : _T_31780; // @[Mux.scala 31:69:@11806.4]
  assign _T_31782 = valid_36_49 ? 6'h31 : _T_31781; // @[Mux.scala 31:69:@11807.4]
  assign _T_31783 = valid_36_48 ? 6'h30 : _T_31782; // @[Mux.scala 31:69:@11808.4]
  assign _T_31784 = valid_36_47 ? 6'h2f : _T_31783; // @[Mux.scala 31:69:@11809.4]
  assign _T_31785 = valid_36_46 ? 6'h2e : _T_31784; // @[Mux.scala 31:69:@11810.4]
  assign _T_31786 = valid_36_45 ? 6'h2d : _T_31785; // @[Mux.scala 31:69:@11811.4]
  assign _T_31787 = valid_36_44 ? 6'h2c : _T_31786; // @[Mux.scala 31:69:@11812.4]
  assign _T_31788 = valid_36_43 ? 6'h2b : _T_31787; // @[Mux.scala 31:69:@11813.4]
  assign _T_31789 = valid_36_42 ? 6'h2a : _T_31788; // @[Mux.scala 31:69:@11814.4]
  assign _T_31790 = valid_36_41 ? 6'h29 : _T_31789; // @[Mux.scala 31:69:@11815.4]
  assign _T_31791 = valid_36_40 ? 6'h28 : _T_31790; // @[Mux.scala 31:69:@11816.4]
  assign _T_31792 = valid_36_39 ? 6'h27 : _T_31791; // @[Mux.scala 31:69:@11817.4]
  assign _T_31793 = valid_36_38 ? 6'h26 : _T_31792; // @[Mux.scala 31:69:@11818.4]
  assign _T_31794 = valid_36_37 ? 6'h25 : _T_31793; // @[Mux.scala 31:69:@11819.4]
  assign _T_31795 = valid_36_36 ? 6'h24 : _T_31794; // @[Mux.scala 31:69:@11820.4]
  assign _T_31796 = valid_36_35 ? 6'h23 : _T_31795; // @[Mux.scala 31:69:@11821.4]
  assign _T_31797 = valid_36_34 ? 6'h22 : _T_31796; // @[Mux.scala 31:69:@11822.4]
  assign _T_31798 = valid_36_33 ? 6'h21 : _T_31797; // @[Mux.scala 31:69:@11823.4]
  assign _T_31799 = valid_36_32 ? 6'h20 : _T_31798; // @[Mux.scala 31:69:@11824.4]
  assign _T_31800 = valid_36_31 ? 6'h1f : _T_31799; // @[Mux.scala 31:69:@11825.4]
  assign _T_31801 = valid_36_30 ? 6'h1e : _T_31800; // @[Mux.scala 31:69:@11826.4]
  assign _T_31802 = valid_36_29 ? 6'h1d : _T_31801; // @[Mux.scala 31:69:@11827.4]
  assign _T_31803 = valid_36_28 ? 6'h1c : _T_31802; // @[Mux.scala 31:69:@11828.4]
  assign _T_31804 = valid_36_27 ? 6'h1b : _T_31803; // @[Mux.scala 31:69:@11829.4]
  assign _T_31805 = valid_36_26 ? 6'h1a : _T_31804; // @[Mux.scala 31:69:@11830.4]
  assign _T_31806 = valid_36_25 ? 6'h19 : _T_31805; // @[Mux.scala 31:69:@11831.4]
  assign _T_31807 = valid_36_24 ? 6'h18 : _T_31806; // @[Mux.scala 31:69:@11832.4]
  assign _T_31808 = valid_36_23 ? 6'h17 : _T_31807; // @[Mux.scala 31:69:@11833.4]
  assign _T_31809 = valid_36_22 ? 6'h16 : _T_31808; // @[Mux.scala 31:69:@11834.4]
  assign _T_31810 = valid_36_21 ? 6'h15 : _T_31809; // @[Mux.scala 31:69:@11835.4]
  assign _T_31811 = valid_36_20 ? 6'h14 : _T_31810; // @[Mux.scala 31:69:@11836.4]
  assign _T_31812 = valid_36_19 ? 6'h13 : _T_31811; // @[Mux.scala 31:69:@11837.4]
  assign _T_31813 = valid_36_18 ? 6'h12 : _T_31812; // @[Mux.scala 31:69:@11838.4]
  assign _T_31814 = valid_36_17 ? 6'h11 : _T_31813; // @[Mux.scala 31:69:@11839.4]
  assign _T_31815 = valid_36_16 ? 6'h10 : _T_31814; // @[Mux.scala 31:69:@11840.4]
  assign _T_31816 = valid_36_15 ? 6'hf : _T_31815; // @[Mux.scala 31:69:@11841.4]
  assign _T_31817 = valid_36_14 ? 6'he : _T_31816; // @[Mux.scala 31:69:@11842.4]
  assign _T_31818 = valid_36_13 ? 6'hd : _T_31817; // @[Mux.scala 31:69:@11843.4]
  assign _T_31819 = valid_36_12 ? 6'hc : _T_31818; // @[Mux.scala 31:69:@11844.4]
  assign _T_31820 = valid_36_11 ? 6'hb : _T_31819; // @[Mux.scala 31:69:@11845.4]
  assign _T_31821 = valid_36_10 ? 6'ha : _T_31820; // @[Mux.scala 31:69:@11846.4]
  assign _T_31822 = valid_36_9 ? 6'h9 : _T_31821; // @[Mux.scala 31:69:@11847.4]
  assign _T_31823 = valid_36_8 ? 6'h8 : _T_31822; // @[Mux.scala 31:69:@11848.4]
  assign _T_31824 = valid_36_7 ? 6'h7 : _T_31823; // @[Mux.scala 31:69:@11849.4]
  assign _T_31825 = valid_36_6 ? 6'h6 : _T_31824; // @[Mux.scala 31:69:@11850.4]
  assign _T_31826 = valid_36_5 ? 6'h5 : _T_31825; // @[Mux.scala 31:69:@11851.4]
  assign _T_31827 = valid_36_4 ? 6'h4 : _T_31826; // @[Mux.scala 31:69:@11852.4]
  assign _T_31828 = valid_36_3 ? 6'h3 : _T_31827; // @[Mux.scala 31:69:@11853.4]
  assign _T_31829 = valid_36_2 ? 6'h2 : _T_31828; // @[Mux.scala 31:69:@11854.4]
  assign _T_31830 = valid_36_1 ? 6'h1 : _T_31829; // @[Mux.scala 31:69:@11855.4]
  assign select_36 = valid_36_0 ? 6'h0 : _T_31830; // @[Mux.scala 31:69:@11856.4]
  assign _GEN_2305 = 6'h1 == select_36 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2306 = 6'h2 == select_36 ? io_inData_2 : _GEN_2305; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2307 = 6'h3 == select_36 ? io_inData_3 : _GEN_2306; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2308 = 6'h4 == select_36 ? io_inData_4 : _GEN_2307; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2309 = 6'h5 == select_36 ? io_inData_5 : _GEN_2308; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2310 = 6'h6 == select_36 ? io_inData_6 : _GEN_2309; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2311 = 6'h7 == select_36 ? io_inData_7 : _GEN_2310; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2312 = 6'h8 == select_36 ? io_inData_8 : _GEN_2311; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2313 = 6'h9 == select_36 ? io_inData_9 : _GEN_2312; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2314 = 6'ha == select_36 ? io_inData_10 : _GEN_2313; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2315 = 6'hb == select_36 ? io_inData_11 : _GEN_2314; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2316 = 6'hc == select_36 ? io_inData_12 : _GEN_2315; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2317 = 6'hd == select_36 ? io_inData_13 : _GEN_2316; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2318 = 6'he == select_36 ? io_inData_14 : _GEN_2317; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2319 = 6'hf == select_36 ? io_inData_15 : _GEN_2318; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2320 = 6'h10 == select_36 ? io_inData_16 : _GEN_2319; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2321 = 6'h11 == select_36 ? io_inData_17 : _GEN_2320; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2322 = 6'h12 == select_36 ? io_inData_18 : _GEN_2321; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2323 = 6'h13 == select_36 ? io_inData_19 : _GEN_2322; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2324 = 6'h14 == select_36 ? io_inData_20 : _GEN_2323; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2325 = 6'h15 == select_36 ? io_inData_21 : _GEN_2324; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2326 = 6'h16 == select_36 ? io_inData_22 : _GEN_2325; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2327 = 6'h17 == select_36 ? io_inData_23 : _GEN_2326; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2328 = 6'h18 == select_36 ? io_inData_24 : _GEN_2327; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2329 = 6'h19 == select_36 ? io_inData_25 : _GEN_2328; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2330 = 6'h1a == select_36 ? io_inData_26 : _GEN_2329; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2331 = 6'h1b == select_36 ? io_inData_27 : _GEN_2330; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2332 = 6'h1c == select_36 ? io_inData_28 : _GEN_2331; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2333 = 6'h1d == select_36 ? io_inData_29 : _GEN_2332; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2334 = 6'h1e == select_36 ? io_inData_30 : _GEN_2333; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2335 = 6'h1f == select_36 ? io_inData_31 : _GEN_2334; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2336 = 6'h20 == select_36 ? io_inData_32 : _GEN_2335; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2337 = 6'h21 == select_36 ? io_inData_33 : _GEN_2336; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2338 = 6'h22 == select_36 ? io_inData_34 : _GEN_2337; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2339 = 6'h23 == select_36 ? io_inData_35 : _GEN_2338; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2340 = 6'h24 == select_36 ? io_inData_36 : _GEN_2339; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2341 = 6'h25 == select_36 ? io_inData_37 : _GEN_2340; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2342 = 6'h26 == select_36 ? io_inData_38 : _GEN_2341; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2343 = 6'h27 == select_36 ? io_inData_39 : _GEN_2342; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2344 = 6'h28 == select_36 ? io_inData_40 : _GEN_2343; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2345 = 6'h29 == select_36 ? io_inData_41 : _GEN_2344; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2346 = 6'h2a == select_36 ? io_inData_42 : _GEN_2345; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2347 = 6'h2b == select_36 ? io_inData_43 : _GEN_2346; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2348 = 6'h2c == select_36 ? io_inData_44 : _GEN_2347; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2349 = 6'h2d == select_36 ? io_inData_45 : _GEN_2348; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2350 = 6'h2e == select_36 ? io_inData_46 : _GEN_2349; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2351 = 6'h2f == select_36 ? io_inData_47 : _GEN_2350; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2352 = 6'h30 == select_36 ? io_inData_48 : _GEN_2351; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2353 = 6'h31 == select_36 ? io_inData_49 : _GEN_2352; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2354 = 6'h32 == select_36 ? io_inData_50 : _GEN_2353; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2355 = 6'h33 == select_36 ? io_inData_51 : _GEN_2354; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2356 = 6'h34 == select_36 ? io_inData_52 : _GEN_2355; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2357 = 6'h35 == select_36 ? io_inData_53 : _GEN_2356; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2358 = 6'h36 == select_36 ? io_inData_54 : _GEN_2357; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2359 = 6'h37 == select_36 ? io_inData_55 : _GEN_2358; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2360 = 6'h38 == select_36 ? io_inData_56 : _GEN_2359; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2361 = 6'h39 == select_36 ? io_inData_57 : _GEN_2360; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2362 = 6'h3a == select_36 ? io_inData_58 : _GEN_2361; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2363 = 6'h3b == select_36 ? io_inData_59 : _GEN_2362; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2364 = 6'h3c == select_36 ? io_inData_60 : _GEN_2363; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2365 = 6'h3d == select_36 ? io_inData_61 : _GEN_2364; // @[Switch.scala 33:19:@11858.4]
  assign _GEN_2366 = 6'h3e == select_36 ? io_inData_62 : _GEN_2365; // @[Switch.scala 33:19:@11858.4]
  assign _T_31839 = {valid_36_7,valid_36_6,valid_36_5,valid_36_4,valid_36_3,valid_36_2,valid_36_1,valid_36_0}; // @[Switch.scala 34:32:@11865.4]
  assign _T_31847 = {valid_36_15,valid_36_14,valid_36_13,valid_36_12,valid_36_11,valid_36_10,valid_36_9,valid_36_8,_T_31839}; // @[Switch.scala 34:32:@11873.4]
  assign _T_31854 = {valid_36_23,valid_36_22,valid_36_21,valid_36_20,valid_36_19,valid_36_18,valid_36_17,valid_36_16}; // @[Switch.scala 34:32:@11880.4]
  assign _T_31863 = {valid_36_31,valid_36_30,valid_36_29,valid_36_28,valid_36_27,valid_36_26,valid_36_25,valid_36_24,_T_31854,_T_31847}; // @[Switch.scala 34:32:@11889.4]
  assign _T_31870 = {valid_36_39,valid_36_38,valid_36_37,valid_36_36,valid_36_35,valid_36_34,valid_36_33,valid_36_32}; // @[Switch.scala 34:32:@11896.4]
  assign _T_31878 = {valid_36_47,valid_36_46,valid_36_45,valid_36_44,valid_36_43,valid_36_42,valid_36_41,valid_36_40,_T_31870}; // @[Switch.scala 34:32:@11904.4]
  assign _T_31885 = {valid_36_55,valid_36_54,valid_36_53,valid_36_52,valid_36_51,valid_36_50,valid_36_49,valid_36_48}; // @[Switch.scala 34:32:@11911.4]
  assign _T_31894 = {valid_36_63,valid_36_62,valid_36_61,valid_36_60,valid_36_59,valid_36_58,valid_36_57,valid_36_56,_T_31885,_T_31878}; // @[Switch.scala 34:32:@11920.4]
  assign _T_31895 = {_T_31894,_T_31863}; // @[Switch.scala 34:32:@11921.4]
  assign _T_31899 = io_inAddr_0 == 6'h25; // @[Switch.scala 30:53:@11924.4]
  assign valid_37_0 = io_inValid_0 & _T_31899; // @[Switch.scala 30:36:@11925.4]
  assign _T_31902 = io_inAddr_1 == 6'h25; // @[Switch.scala 30:53:@11927.4]
  assign valid_37_1 = io_inValid_1 & _T_31902; // @[Switch.scala 30:36:@11928.4]
  assign _T_31905 = io_inAddr_2 == 6'h25; // @[Switch.scala 30:53:@11930.4]
  assign valid_37_2 = io_inValid_2 & _T_31905; // @[Switch.scala 30:36:@11931.4]
  assign _T_31908 = io_inAddr_3 == 6'h25; // @[Switch.scala 30:53:@11933.4]
  assign valid_37_3 = io_inValid_3 & _T_31908; // @[Switch.scala 30:36:@11934.4]
  assign _T_31911 = io_inAddr_4 == 6'h25; // @[Switch.scala 30:53:@11936.4]
  assign valid_37_4 = io_inValid_4 & _T_31911; // @[Switch.scala 30:36:@11937.4]
  assign _T_31914 = io_inAddr_5 == 6'h25; // @[Switch.scala 30:53:@11939.4]
  assign valid_37_5 = io_inValid_5 & _T_31914; // @[Switch.scala 30:36:@11940.4]
  assign _T_31917 = io_inAddr_6 == 6'h25; // @[Switch.scala 30:53:@11942.4]
  assign valid_37_6 = io_inValid_6 & _T_31917; // @[Switch.scala 30:36:@11943.4]
  assign _T_31920 = io_inAddr_7 == 6'h25; // @[Switch.scala 30:53:@11945.4]
  assign valid_37_7 = io_inValid_7 & _T_31920; // @[Switch.scala 30:36:@11946.4]
  assign _T_31923 = io_inAddr_8 == 6'h25; // @[Switch.scala 30:53:@11948.4]
  assign valid_37_8 = io_inValid_8 & _T_31923; // @[Switch.scala 30:36:@11949.4]
  assign _T_31926 = io_inAddr_9 == 6'h25; // @[Switch.scala 30:53:@11951.4]
  assign valid_37_9 = io_inValid_9 & _T_31926; // @[Switch.scala 30:36:@11952.4]
  assign _T_31929 = io_inAddr_10 == 6'h25; // @[Switch.scala 30:53:@11954.4]
  assign valid_37_10 = io_inValid_10 & _T_31929; // @[Switch.scala 30:36:@11955.4]
  assign _T_31932 = io_inAddr_11 == 6'h25; // @[Switch.scala 30:53:@11957.4]
  assign valid_37_11 = io_inValid_11 & _T_31932; // @[Switch.scala 30:36:@11958.4]
  assign _T_31935 = io_inAddr_12 == 6'h25; // @[Switch.scala 30:53:@11960.4]
  assign valid_37_12 = io_inValid_12 & _T_31935; // @[Switch.scala 30:36:@11961.4]
  assign _T_31938 = io_inAddr_13 == 6'h25; // @[Switch.scala 30:53:@11963.4]
  assign valid_37_13 = io_inValid_13 & _T_31938; // @[Switch.scala 30:36:@11964.4]
  assign _T_31941 = io_inAddr_14 == 6'h25; // @[Switch.scala 30:53:@11966.4]
  assign valid_37_14 = io_inValid_14 & _T_31941; // @[Switch.scala 30:36:@11967.4]
  assign _T_31944 = io_inAddr_15 == 6'h25; // @[Switch.scala 30:53:@11969.4]
  assign valid_37_15 = io_inValid_15 & _T_31944; // @[Switch.scala 30:36:@11970.4]
  assign _T_31947 = io_inAddr_16 == 6'h25; // @[Switch.scala 30:53:@11972.4]
  assign valid_37_16 = io_inValid_16 & _T_31947; // @[Switch.scala 30:36:@11973.4]
  assign _T_31950 = io_inAddr_17 == 6'h25; // @[Switch.scala 30:53:@11975.4]
  assign valid_37_17 = io_inValid_17 & _T_31950; // @[Switch.scala 30:36:@11976.4]
  assign _T_31953 = io_inAddr_18 == 6'h25; // @[Switch.scala 30:53:@11978.4]
  assign valid_37_18 = io_inValid_18 & _T_31953; // @[Switch.scala 30:36:@11979.4]
  assign _T_31956 = io_inAddr_19 == 6'h25; // @[Switch.scala 30:53:@11981.4]
  assign valid_37_19 = io_inValid_19 & _T_31956; // @[Switch.scala 30:36:@11982.4]
  assign _T_31959 = io_inAddr_20 == 6'h25; // @[Switch.scala 30:53:@11984.4]
  assign valid_37_20 = io_inValid_20 & _T_31959; // @[Switch.scala 30:36:@11985.4]
  assign _T_31962 = io_inAddr_21 == 6'h25; // @[Switch.scala 30:53:@11987.4]
  assign valid_37_21 = io_inValid_21 & _T_31962; // @[Switch.scala 30:36:@11988.4]
  assign _T_31965 = io_inAddr_22 == 6'h25; // @[Switch.scala 30:53:@11990.4]
  assign valid_37_22 = io_inValid_22 & _T_31965; // @[Switch.scala 30:36:@11991.4]
  assign _T_31968 = io_inAddr_23 == 6'h25; // @[Switch.scala 30:53:@11993.4]
  assign valid_37_23 = io_inValid_23 & _T_31968; // @[Switch.scala 30:36:@11994.4]
  assign _T_31971 = io_inAddr_24 == 6'h25; // @[Switch.scala 30:53:@11996.4]
  assign valid_37_24 = io_inValid_24 & _T_31971; // @[Switch.scala 30:36:@11997.4]
  assign _T_31974 = io_inAddr_25 == 6'h25; // @[Switch.scala 30:53:@11999.4]
  assign valid_37_25 = io_inValid_25 & _T_31974; // @[Switch.scala 30:36:@12000.4]
  assign _T_31977 = io_inAddr_26 == 6'h25; // @[Switch.scala 30:53:@12002.4]
  assign valid_37_26 = io_inValid_26 & _T_31977; // @[Switch.scala 30:36:@12003.4]
  assign _T_31980 = io_inAddr_27 == 6'h25; // @[Switch.scala 30:53:@12005.4]
  assign valid_37_27 = io_inValid_27 & _T_31980; // @[Switch.scala 30:36:@12006.4]
  assign _T_31983 = io_inAddr_28 == 6'h25; // @[Switch.scala 30:53:@12008.4]
  assign valid_37_28 = io_inValid_28 & _T_31983; // @[Switch.scala 30:36:@12009.4]
  assign _T_31986 = io_inAddr_29 == 6'h25; // @[Switch.scala 30:53:@12011.4]
  assign valid_37_29 = io_inValid_29 & _T_31986; // @[Switch.scala 30:36:@12012.4]
  assign _T_31989 = io_inAddr_30 == 6'h25; // @[Switch.scala 30:53:@12014.4]
  assign valid_37_30 = io_inValid_30 & _T_31989; // @[Switch.scala 30:36:@12015.4]
  assign _T_31992 = io_inAddr_31 == 6'h25; // @[Switch.scala 30:53:@12017.4]
  assign valid_37_31 = io_inValid_31 & _T_31992; // @[Switch.scala 30:36:@12018.4]
  assign _T_31995 = io_inAddr_32 == 6'h25; // @[Switch.scala 30:53:@12020.4]
  assign valid_37_32 = io_inValid_32 & _T_31995; // @[Switch.scala 30:36:@12021.4]
  assign _T_31998 = io_inAddr_33 == 6'h25; // @[Switch.scala 30:53:@12023.4]
  assign valid_37_33 = io_inValid_33 & _T_31998; // @[Switch.scala 30:36:@12024.4]
  assign _T_32001 = io_inAddr_34 == 6'h25; // @[Switch.scala 30:53:@12026.4]
  assign valid_37_34 = io_inValid_34 & _T_32001; // @[Switch.scala 30:36:@12027.4]
  assign _T_32004 = io_inAddr_35 == 6'h25; // @[Switch.scala 30:53:@12029.4]
  assign valid_37_35 = io_inValid_35 & _T_32004; // @[Switch.scala 30:36:@12030.4]
  assign _T_32007 = io_inAddr_36 == 6'h25; // @[Switch.scala 30:53:@12032.4]
  assign valid_37_36 = io_inValid_36 & _T_32007; // @[Switch.scala 30:36:@12033.4]
  assign _T_32010 = io_inAddr_37 == 6'h25; // @[Switch.scala 30:53:@12035.4]
  assign valid_37_37 = io_inValid_37 & _T_32010; // @[Switch.scala 30:36:@12036.4]
  assign _T_32013 = io_inAddr_38 == 6'h25; // @[Switch.scala 30:53:@12038.4]
  assign valid_37_38 = io_inValid_38 & _T_32013; // @[Switch.scala 30:36:@12039.4]
  assign _T_32016 = io_inAddr_39 == 6'h25; // @[Switch.scala 30:53:@12041.4]
  assign valid_37_39 = io_inValid_39 & _T_32016; // @[Switch.scala 30:36:@12042.4]
  assign _T_32019 = io_inAddr_40 == 6'h25; // @[Switch.scala 30:53:@12044.4]
  assign valid_37_40 = io_inValid_40 & _T_32019; // @[Switch.scala 30:36:@12045.4]
  assign _T_32022 = io_inAddr_41 == 6'h25; // @[Switch.scala 30:53:@12047.4]
  assign valid_37_41 = io_inValid_41 & _T_32022; // @[Switch.scala 30:36:@12048.4]
  assign _T_32025 = io_inAddr_42 == 6'h25; // @[Switch.scala 30:53:@12050.4]
  assign valid_37_42 = io_inValid_42 & _T_32025; // @[Switch.scala 30:36:@12051.4]
  assign _T_32028 = io_inAddr_43 == 6'h25; // @[Switch.scala 30:53:@12053.4]
  assign valid_37_43 = io_inValid_43 & _T_32028; // @[Switch.scala 30:36:@12054.4]
  assign _T_32031 = io_inAddr_44 == 6'h25; // @[Switch.scala 30:53:@12056.4]
  assign valid_37_44 = io_inValid_44 & _T_32031; // @[Switch.scala 30:36:@12057.4]
  assign _T_32034 = io_inAddr_45 == 6'h25; // @[Switch.scala 30:53:@12059.4]
  assign valid_37_45 = io_inValid_45 & _T_32034; // @[Switch.scala 30:36:@12060.4]
  assign _T_32037 = io_inAddr_46 == 6'h25; // @[Switch.scala 30:53:@12062.4]
  assign valid_37_46 = io_inValid_46 & _T_32037; // @[Switch.scala 30:36:@12063.4]
  assign _T_32040 = io_inAddr_47 == 6'h25; // @[Switch.scala 30:53:@12065.4]
  assign valid_37_47 = io_inValid_47 & _T_32040; // @[Switch.scala 30:36:@12066.4]
  assign _T_32043 = io_inAddr_48 == 6'h25; // @[Switch.scala 30:53:@12068.4]
  assign valid_37_48 = io_inValid_48 & _T_32043; // @[Switch.scala 30:36:@12069.4]
  assign _T_32046 = io_inAddr_49 == 6'h25; // @[Switch.scala 30:53:@12071.4]
  assign valid_37_49 = io_inValid_49 & _T_32046; // @[Switch.scala 30:36:@12072.4]
  assign _T_32049 = io_inAddr_50 == 6'h25; // @[Switch.scala 30:53:@12074.4]
  assign valid_37_50 = io_inValid_50 & _T_32049; // @[Switch.scala 30:36:@12075.4]
  assign _T_32052 = io_inAddr_51 == 6'h25; // @[Switch.scala 30:53:@12077.4]
  assign valid_37_51 = io_inValid_51 & _T_32052; // @[Switch.scala 30:36:@12078.4]
  assign _T_32055 = io_inAddr_52 == 6'h25; // @[Switch.scala 30:53:@12080.4]
  assign valid_37_52 = io_inValid_52 & _T_32055; // @[Switch.scala 30:36:@12081.4]
  assign _T_32058 = io_inAddr_53 == 6'h25; // @[Switch.scala 30:53:@12083.4]
  assign valid_37_53 = io_inValid_53 & _T_32058; // @[Switch.scala 30:36:@12084.4]
  assign _T_32061 = io_inAddr_54 == 6'h25; // @[Switch.scala 30:53:@12086.4]
  assign valid_37_54 = io_inValid_54 & _T_32061; // @[Switch.scala 30:36:@12087.4]
  assign _T_32064 = io_inAddr_55 == 6'h25; // @[Switch.scala 30:53:@12089.4]
  assign valid_37_55 = io_inValid_55 & _T_32064; // @[Switch.scala 30:36:@12090.4]
  assign _T_32067 = io_inAddr_56 == 6'h25; // @[Switch.scala 30:53:@12092.4]
  assign valid_37_56 = io_inValid_56 & _T_32067; // @[Switch.scala 30:36:@12093.4]
  assign _T_32070 = io_inAddr_57 == 6'h25; // @[Switch.scala 30:53:@12095.4]
  assign valid_37_57 = io_inValid_57 & _T_32070; // @[Switch.scala 30:36:@12096.4]
  assign _T_32073 = io_inAddr_58 == 6'h25; // @[Switch.scala 30:53:@12098.4]
  assign valid_37_58 = io_inValid_58 & _T_32073; // @[Switch.scala 30:36:@12099.4]
  assign _T_32076 = io_inAddr_59 == 6'h25; // @[Switch.scala 30:53:@12101.4]
  assign valid_37_59 = io_inValid_59 & _T_32076; // @[Switch.scala 30:36:@12102.4]
  assign _T_32079 = io_inAddr_60 == 6'h25; // @[Switch.scala 30:53:@12104.4]
  assign valid_37_60 = io_inValid_60 & _T_32079; // @[Switch.scala 30:36:@12105.4]
  assign _T_32082 = io_inAddr_61 == 6'h25; // @[Switch.scala 30:53:@12107.4]
  assign valid_37_61 = io_inValid_61 & _T_32082; // @[Switch.scala 30:36:@12108.4]
  assign _T_32085 = io_inAddr_62 == 6'h25; // @[Switch.scala 30:53:@12110.4]
  assign valid_37_62 = io_inValid_62 & _T_32085; // @[Switch.scala 30:36:@12111.4]
  assign _T_32088 = io_inAddr_63 == 6'h25; // @[Switch.scala 30:53:@12113.4]
  assign valid_37_63 = io_inValid_63 & _T_32088; // @[Switch.scala 30:36:@12114.4]
  assign _T_32154 = valid_37_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@12116.4]
  assign _T_32155 = valid_37_61 ? 6'h3d : _T_32154; // @[Mux.scala 31:69:@12117.4]
  assign _T_32156 = valid_37_60 ? 6'h3c : _T_32155; // @[Mux.scala 31:69:@12118.4]
  assign _T_32157 = valid_37_59 ? 6'h3b : _T_32156; // @[Mux.scala 31:69:@12119.4]
  assign _T_32158 = valid_37_58 ? 6'h3a : _T_32157; // @[Mux.scala 31:69:@12120.4]
  assign _T_32159 = valid_37_57 ? 6'h39 : _T_32158; // @[Mux.scala 31:69:@12121.4]
  assign _T_32160 = valid_37_56 ? 6'h38 : _T_32159; // @[Mux.scala 31:69:@12122.4]
  assign _T_32161 = valid_37_55 ? 6'h37 : _T_32160; // @[Mux.scala 31:69:@12123.4]
  assign _T_32162 = valid_37_54 ? 6'h36 : _T_32161; // @[Mux.scala 31:69:@12124.4]
  assign _T_32163 = valid_37_53 ? 6'h35 : _T_32162; // @[Mux.scala 31:69:@12125.4]
  assign _T_32164 = valid_37_52 ? 6'h34 : _T_32163; // @[Mux.scala 31:69:@12126.4]
  assign _T_32165 = valid_37_51 ? 6'h33 : _T_32164; // @[Mux.scala 31:69:@12127.4]
  assign _T_32166 = valid_37_50 ? 6'h32 : _T_32165; // @[Mux.scala 31:69:@12128.4]
  assign _T_32167 = valid_37_49 ? 6'h31 : _T_32166; // @[Mux.scala 31:69:@12129.4]
  assign _T_32168 = valid_37_48 ? 6'h30 : _T_32167; // @[Mux.scala 31:69:@12130.4]
  assign _T_32169 = valid_37_47 ? 6'h2f : _T_32168; // @[Mux.scala 31:69:@12131.4]
  assign _T_32170 = valid_37_46 ? 6'h2e : _T_32169; // @[Mux.scala 31:69:@12132.4]
  assign _T_32171 = valid_37_45 ? 6'h2d : _T_32170; // @[Mux.scala 31:69:@12133.4]
  assign _T_32172 = valid_37_44 ? 6'h2c : _T_32171; // @[Mux.scala 31:69:@12134.4]
  assign _T_32173 = valid_37_43 ? 6'h2b : _T_32172; // @[Mux.scala 31:69:@12135.4]
  assign _T_32174 = valid_37_42 ? 6'h2a : _T_32173; // @[Mux.scala 31:69:@12136.4]
  assign _T_32175 = valid_37_41 ? 6'h29 : _T_32174; // @[Mux.scala 31:69:@12137.4]
  assign _T_32176 = valid_37_40 ? 6'h28 : _T_32175; // @[Mux.scala 31:69:@12138.4]
  assign _T_32177 = valid_37_39 ? 6'h27 : _T_32176; // @[Mux.scala 31:69:@12139.4]
  assign _T_32178 = valid_37_38 ? 6'h26 : _T_32177; // @[Mux.scala 31:69:@12140.4]
  assign _T_32179 = valid_37_37 ? 6'h25 : _T_32178; // @[Mux.scala 31:69:@12141.4]
  assign _T_32180 = valid_37_36 ? 6'h24 : _T_32179; // @[Mux.scala 31:69:@12142.4]
  assign _T_32181 = valid_37_35 ? 6'h23 : _T_32180; // @[Mux.scala 31:69:@12143.4]
  assign _T_32182 = valid_37_34 ? 6'h22 : _T_32181; // @[Mux.scala 31:69:@12144.4]
  assign _T_32183 = valid_37_33 ? 6'h21 : _T_32182; // @[Mux.scala 31:69:@12145.4]
  assign _T_32184 = valid_37_32 ? 6'h20 : _T_32183; // @[Mux.scala 31:69:@12146.4]
  assign _T_32185 = valid_37_31 ? 6'h1f : _T_32184; // @[Mux.scala 31:69:@12147.4]
  assign _T_32186 = valid_37_30 ? 6'h1e : _T_32185; // @[Mux.scala 31:69:@12148.4]
  assign _T_32187 = valid_37_29 ? 6'h1d : _T_32186; // @[Mux.scala 31:69:@12149.4]
  assign _T_32188 = valid_37_28 ? 6'h1c : _T_32187; // @[Mux.scala 31:69:@12150.4]
  assign _T_32189 = valid_37_27 ? 6'h1b : _T_32188; // @[Mux.scala 31:69:@12151.4]
  assign _T_32190 = valid_37_26 ? 6'h1a : _T_32189; // @[Mux.scala 31:69:@12152.4]
  assign _T_32191 = valid_37_25 ? 6'h19 : _T_32190; // @[Mux.scala 31:69:@12153.4]
  assign _T_32192 = valid_37_24 ? 6'h18 : _T_32191; // @[Mux.scala 31:69:@12154.4]
  assign _T_32193 = valid_37_23 ? 6'h17 : _T_32192; // @[Mux.scala 31:69:@12155.4]
  assign _T_32194 = valid_37_22 ? 6'h16 : _T_32193; // @[Mux.scala 31:69:@12156.4]
  assign _T_32195 = valid_37_21 ? 6'h15 : _T_32194; // @[Mux.scala 31:69:@12157.4]
  assign _T_32196 = valid_37_20 ? 6'h14 : _T_32195; // @[Mux.scala 31:69:@12158.4]
  assign _T_32197 = valid_37_19 ? 6'h13 : _T_32196; // @[Mux.scala 31:69:@12159.4]
  assign _T_32198 = valid_37_18 ? 6'h12 : _T_32197; // @[Mux.scala 31:69:@12160.4]
  assign _T_32199 = valid_37_17 ? 6'h11 : _T_32198; // @[Mux.scala 31:69:@12161.4]
  assign _T_32200 = valid_37_16 ? 6'h10 : _T_32199; // @[Mux.scala 31:69:@12162.4]
  assign _T_32201 = valid_37_15 ? 6'hf : _T_32200; // @[Mux.scala 31:69:@12163.4]
  assign _T_32202 = valid_37_14 ? 6'he : _T_32201; // @[Mux.scala 31:69:@12164.4]
  assign _T_32203 = valid_37_13 ? 6'hd : _T_32202; // @[Mux.scala 31:69:@12165.4]
  assign _T_32204 = valid_37_12 ? 6'hc : _T_32203; // @[Mux.scala 31:69:@12166.4]
  assign _T_32205 = valid_37_11 ? 6'hb : _T_32204; // @[Mux.scala 31:69:@12167.4]
  assign _T_32206 = valid_37_10 ? 6'ha : _T_32205; // @[Mux.scala 31:69:@12168.4]
  assign _T_32207 = valid_37_9 ? 6'h9 : _T_32206; // @[Mux.scala 31:69:@12169.4]
  assign _T_32208 = valid_37_8 ? 6'h8 : _T_32207; // @[Mux.scala 31:69:@12170.4]
  assign _T_32209 = valid_37_7 ? 6'h7 : _T_32208; // @[Mux.scala 31:69:@12171.4]
  assign _T_32210 = valid_37_6 ? 6'h6 : _T_32209; // @[Mux.scala 31:69:@12172.4]
  assign _T_32211 = valid_37_5 ? 6'h5 : _T_32210; // @[Mux.scala 31:69:@12173.4]
  assign _T_32212 = valid_37_4 ? 6'h4 : _T_32211; // @[Mux.scala 31:69:@12174.4]
  assign _T_32213 = valid_37_3 ? 6'h3 : _T_32212; // @[Mux.scala 31:69:@12175.4]
  assign _T_32214 = valid_37_2 ? 6'h2 : _T_32213; // @[Mux.scala 31:69:@12176.4]
  assign _T_32215 = valid_37_1 ? 6'h1 : _T_32214; // @[Mux.scala 31:69:@12177.4]
  assign select_37 = valid_37_0 ? 6'h0 : _T_32215; // @[Mux.scala 31:69:@12178.4]
  assign _GEN_2369 = 6'h1 == select_37 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2370 = 6'h2 == select_37 ? io_inData_2 : _GEN_2369; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2371 = 6'h3 == select_37 ? io_inData_3 : _GEN_2370; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2372 = 6'h4 == select_37 ? io_inData_4 : _GEN_2371; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2373 = 6'h5 == select_37 ? io_inData_5 : _GEN_2372; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2374 = 6'h6 == select_37 ? io_inData_6 : _GEN_2373; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2375 = 6'h7 == select_37 ? io_inData_7 : _GEN_2374; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2376 = 6'h8 == select_37 ? io_inData_8 : _GEN_2375; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2377 = 6'h9 == select_37 ? io_inData_9 : _GEN_2376; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2378 = 6'ha == select_37 ? io_inData_10 : _GEN_2377; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2379 = 6'hb == select_37 ? io_inData_11 : _GEN_2378; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2380 = 6'hc == select_37 ? io_inData_12 : _GEN_2379; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2381 = 6'hd == select_37 ? io_inData_13 : _GEN_2380; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2382 = 6'he == select_37 ? io_inData_14 : _GEN_2381; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2383 = 6'hf == select_37 ? io_inData_15 : _GEN_2382; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2384 = 6'h10 == select_37 ? io_inData_16 : _GEN_2383; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2385 = 6'h11 == select_37 ? io_inData_17 : _GEN_2384; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2386 = 6'h12 == select_37 ? io_inData_18 : _GEN_2385; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2387 = 6'h13 == select_37 ? io_inData_19 : _GEN_2386; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2388 = 6'h14 == select_37 ? io_inData_20 : _GEN_2387; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2389 = 6'h15 == select_37 ? io_inData_21 : _GEN_2388; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2390 = 6'h16 == select_37 ? io_inData_22 : _GEN_2389; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2391 = 6'h17 == select_37 ? io_inData_23 : _GEN_2390; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2392 = 6'h18 == select_37 ? io_inData_24 : _GEN_2391; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2393 = 6'h19 == select_37 ? io_inData_25 : _GEN_2392; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2394 = 6'h1a == select_37 ? io_inData_26 : _GEN_2393; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2395 = 6'h1b == select_37 ? io_inData_27 : _GEN_2394; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2396 = 6'h1c == select_37 ? io_inData_28 : _GEN_2395; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2397 = 6'h1d == select_37 ? io_inData_29 : _GEN_2396; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2398 = 6'h1e == select_37 ? io_inData_30 : _GEN_2397; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2399 = 6'h1f == select_37 ? io_inData_31 : _GEN_2398; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2400 = 6'h20 == select_37 ? io_inData_32 : _GEN_2399; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2401 = 6'h21 == select_37 ? io_inData_33 : _GEN_2400; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2402 = 6'h22 == select_37 ? io_inData_34 : _GEN_2401; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2403 = 6'h23 == select_37 ? io_inData_35 : _GEN_2402; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2404 = 6'h24 == select_37 ? io_inData_36 : _GEN_2403; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2405 = 6'h25 == select_37 ? io_inData_37 : _GEN_2404; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2406 = 6'h26 == select_37 ? io_inData_38 : _GEN_2405; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2407 = 6'h27 == select_37 ? io_inData_39 : _GEN_2406; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2408 = 6'h28 == select_37 ? io_inData_40 : _GEN_2407; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2409 = 6'h29 == select_37 ? io_inData_41 : _GEN_2408; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2410 = 6'h2a == select_37 ? io_inData_42 : _GEN_2409; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2411 = 6'h2b == select_37 ? io_inData_43 : _GEN_2410; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2412 = 6'h2c == select_37 ? io_inData_44 : _GEN_2411; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2413 = 6'h2d == select_37 ? io_inData_45 : _GEN_2412; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2414 = 6'h2e == select_37 ? io_inData_46 : _GEN_2413; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2415 = 6'h2f == select_37 ? io_inData_47 : _GEN_2414; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2416 = 6'h30 == select_37 ? io_inData_48 : _GEN_2415; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2417 = 6'h31 == select_37 ? io_inData_49 : _GEN_2416; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2418 = 6'h32 == select_37 ? io_inData_50 : _GEN_2417; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2419 = 6'h33 == select_37 ? io_inData_51 : _GEN_2418; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2420 = 6'h34 == select_37 ? io_inData_52 : _GEN_2419; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2421 = 6'h35 == select_37 ? io_inData_53 : _GEN_2420; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2422 = 6'h36 == select_37 ? io_inData_54 : _GEN_2421; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2423 = 6'h37 == select_37 ? io_inData_55 : _GEN_2422; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2424 = 6'h38 == select_37 ? io_inData_56 : _GEN_2423; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2425 = 6'h39 == select_37 ? io_inData_57 : _GEN_2424; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2426 = 6'h3a == select_37 ? io_inData_58 : _GEN_2425; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2427 = 6'h3b == select_37 ? io_inData_59 : _GEN_2426; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2428 = 6'h3c == select_37 ? io_inData_60 : _GEN_2427; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2429 = 6'h3d == select_37 ? io_inData_61 : _GEN_2428; // @[Switch.scala 33:19:@12180.4]
  assign _GEN_2430 = 6'h3e == select_37 ? io_inData_62 : _GEN_2429; // @[Switch.scala 33:19:@12180.4]
  assign _T_32224 = {valid_37_7,valid_37_6,valid_37_5,valid_37_4,valid_37_3,valid_37_2,valid_37_1,valid_37_0}; // @[Switch.scala 34:32:@12187.4]
  assign _T_32232 = {valid_37_15,valid_37_14,valid_37_13,valid_37_12,valid_37_11,valid_37_10,valid_37_9,valid_37_8,_T_32224}; // @[Switch.scala 34:32:@12195.4]
  assign _T_32239 = {valid_37_23,valid_37_22,valid_37_21,valid_37_20,valid_37_19,valid_37_18,valid_37_17,valid_37_16}; // @[Switch.scala 34:32:@12202.4]
  assign _T_32248 = {valid_37_31,valid_37_30,valid_37_29,valid_37_28,valid_37_27,valid_37_26,valid_37_25,valid_37_24,_T_32239,_T_32232}; // @[Switch.scala 34:32:@12211.4]
  assign _T_32255 = {valid_37_39,valid_37_38,valid_37_37,valid_37_36,valid_37_35,valid_37_34,valid_37_33,valid_37_32}; // @[Switch.scala 34:32:@12218.4]
  assign _T_32263 = {valid_37_47,valid_37_46,valid_37_45,valid_37_44,valid_37_43,valid_37_42,valid_37_41,valid_37_40,_T_32255}; // @[Switch.scala 34:32:@12226.4]
  assign _T_32270 = {valid_37_55,valid_37_54,valid_37_53,valid_37_52,valid_37_51,valid_37_50,valid_37_49,valid_37_48}; // @[Switch.scala 34:32:@12233.4]
  assign _T_32279 = {valid_37_63,valid_37_62,valid_37_61,valid_37_60,valid_37_59,valid_37_58,valid_37_57,valid_37_56,_T_32270,_T_32263}; // @[Switch.scala 34:32:@12242.4]
  assign _T_32280 = {_T_32279,_T_32248}; // @[Switch.scala 34:32:@12243.4]
  assign _T_32284 = io_inAddr_0 == 6'h26; // @[Switch.scala 30:53:@12246.4]
  assign valid_38_0 = io_inValid_0 & _T_32284; // @[Switch.scala 30:36:@12247.4]
  assign _T_32287 = io_inAddr_1 == 6'h26; // @[Switch.scala 30:53:@12249.4]
  assign valid_38_1 = io_inValid_1 & _T_32287; // @[Switch.scala 30:36:@12250.4]
  assign _T_32290 = io_inAddr_2 == 6'h26; // @[Switch.scala 30:53:@12252.4]
  assign valid_38_2 = io_inValid_2 & _T_32290; // @[Switch.scala 30:36:@12253.4]
  assign _T_32293 = io_inAddr_3 == 6'h26; // @[Switch.scala 30:53:@12255.4]
  assign valid_38_3 = io_inValid_3 & _T_32293; // @[Switch.scala 30:36:@12256.4]
  assign _T_32296 = io_inAddr_4 == 6'h26; // @[Switch.scala 30:53:@12258.4]
  assign valid_38_4 = io_inValid_4 & _T_32296; // @[Switch.scala 30:36:@12259.4]
  assign _T_32299 = io_inAddr_5 == 6'h26; // @[Switch.scala 30:53:@12261.4]
  assign valid_38_5 = io_inValid_5 & _T_32299; // @[Switch.scala 30:36:@12262.4]
  assign _T_32302 = io_inAddr_6 == 6'h26; // @[Switch.scala 30:53:@12264.4]
  assign valid_38_6 = io_inValid_6 & _T_32302; // @[Switch.scala 30:36:@12265.4]
  assign _T_32305 = io_inAddr_7 == 6'h26; // @[Switch.scala 30:53:@12267.4]
  assign valid_38_7 = io_inValid_7 & _T_32305; // @[Switch.scala 30:36:@12268.4]
  assign _T_32308 = io_inAddr_8 == 6'h26; // @[Switch.scala 30:53:@12270.4]
  assign valid_38_8 = io_inValid_8 & _T_32308; // @[Switch.scala 30:36:@12271.4]
  assign _T_32311 = io_inAddr_9 == 6'h26; // @[Switch.scala 30:53:@12273.4]
  assign valid_38_9 = io_inValid_9 & _T_32311; // @[Switch.scala 30:36:@12274.4]
  assign _T_32314 = io_inAddr_10 == 6'h26; // @[Switch.scala 30:53:@12276.4]
  assign valid_38_10 = io_inValid_10 & _T_32314; // @[Switch.scala 30:36:@12277.4]
  assign _T_32317 = io_inAddr_11 == 6'h26; // @[Switch.scala 30:53:@12279.4]
  assign valid_38_11 = io_inValid_11 & _T_32317; // @[Switch.scala 30:36:@12280.4]
  assign _T_32320 = io_inAddr_12 == 6'h26; // @[Switch.scala 30:53:@12282.4]
  assign valid_38_12 = io_inValid_12 & _T_32320; // @[Switch.scala 30:36:@12283.4]
  assign _T_32323 = io_inAddr_13 == 6'h26; // @[Switch.scala 30:53:@12285.4]
  assign valid_38_13 = io_inValid_13 & _T_32323; // @[Switch.scala 30:36:@12286.4]
  assign _T_32326 = io_inAddr_14 == 6'h26; // @[Switch.scala 30:53:@12288.4]
  assign valid_38_14 = io_inValid_14 & _T_32326; // @[Switch.scala 30:36:@12289.4]
  assign _T_32329 = io_inAddr_15 == 6'h26; // @[Switch.scala 30:53:@12291.4]
  assign valid_38_15 = io_inValid_15 & _T_32329; // @[Switch.scala 30:36:@12292.4]
  assign _T_32332 = io_inAddr_16 == 6'h26; // @[Switch.scala 30:53:@12294.4]
  assign valid_38_16 = io_inValid_16 & _T_32332; // @[Switch.scala 30:36:@12295.4]
  assign _T_32335 = io_inAddr_17 == 6'h26; // @[Switch.scala 30:53:@12297.4]
  assign valid_38_17 = io_inValid_17 & _T_32335; // @[Switch.scala 30:36:@12298.4]
  assign _T_32338 = io_inAddr_18 == 6'h26; // @[Switch.scala 30:53:@12300.4]
  assign valid_38_18 = io_inValid_18 & _T_32338; // @[Switch.scala 30:36:@12301.4]
  assign _T_32341 = io_inAddr_19 == 6'h26; // @[Switch.scala 30:53:@12303.4]
  assign valid_38_19 = io_inValid_19 & _T_32341; // @[Switch.scala 30:36:@12304.4]
  assign _T_32344 = io_inAddr_20 == 6'h26; // @[Switch.scala 30:53:@12306.4]
  assign valid_38_20 = io_inValid_20 & _T_32344; // @[Switch.scala 30:36:@12307.4]
  assign _T_32347 = io_inAddr_21 == 6'h26; // @[Switch.scala 30:53:@12309.4]
  assign valid_38_21 = io_inValid_21 & _T_32347; // @[Switch.scala 30:36:@12310.4]
  assign _T_32350 = io_inAddr_22 == 6'h26; // @[Switch.scala 30:53:@12312.4]
  assign valid_38_22 = io_inValid_22 & _T_32350; // @[Switch.scala 30:36:@12313.4]
  assign _T_32353 = io_inAddr_23 == 6'h26; // @[Switch.scala 30:53:@12315.4]
  assign valid_38_23 = io_inValid_23 & _T_32353; // @[Switch.scala 30:36:@12316.4]
  assign _T_32356 = io_inAddr_24 == 6'h26; // @[Switch.scala 30:53:@12318.4]
  assign valid_38_24 = io_inValid_24 & _T_32356; // @[Switch.scala 30:36:@12319.4]
  assign _T_32359 = io_inAddr_25 == 6'h26; // @[Switch.scala 30:53:@12321.4]
  assign valid_38_25 = io_inValid_25 & _T_32359; // @[Switch.scala 30:36:@12322.4]
  assign _T_32362 = io_inAddr_26 == 6'h26; // @[Switch.scala 30:53:@12324.4]
  assign valid_38_26 = io_inValid_26 & _T_32362; // @[Switch.scala 30:36:@12325.4]
  assign _T_32365 = io_inAddr_27 == 6'h26; // @[Switch.scala 30:53:@12327.4]
  assign valid_38_27 = io_inValid_27 & _T_32365; // @[Switch.scala 30:36:@12328.4]
  assign _T_32368 = io_inAddr_28 == 6'h26; // @[Switch.scala 30:53:@12330.4]
  assign valid_38_28 = io_inValid_28 & _T_32368; // @[Switch.scala 30:36:@12331.4]
  assign _T_32371 = io_inAddr_29 == 6'h26; // @[Switch.scala 30:53:@12333.4]
  assign valid_38_29 = io_inValid_29 & _T_32371; // @[Switch.scala 30:36:@12334.4]
  assign _T_32374 = io_inAddr_30 == 6'h26; // @[Switch.scala 30:53:@12336.4]
  assign valid_38_30 = io_inValid_30 & _T_32374; // @[Switch.scala 30:36:@12337.4]
  assign _T_32377 = io_inAddr_31 == 6'h26; // @[Switch.scala 30:53:@12339.4]
  assign valid_38_31 = io_inValid_31 & _T_32377; // @[Switch.scala 30:36:@12340.4]
  assign _T_32380 = io_inAddr_32 == 6'h26; // @[Switch.scala 30:53:@12342.4]
  assign valid_38_32 = io_inValid_32 & _T_32380; // @[Switch.scala 30:36:@12343.4]
  assign _T_32383 = io_inAddr_33 == 6'h26; // @[Switch.scala 30:53:@12345.4]
  assign valid_38_33 = io_inValid_33 & _T_32383; // @[Switch.scala 30:36:@12346.4]
  assign _T_32386 = io_inAddr_34 == 6'h26; // @[Switch.scala 30:53:@12348.4]
  assign valid_38_34 = io_inValid_34 & _T_32386; // @[Switch.scala 30:36:@12349.4]
  assign _T_32389 = io_inAddr_35 == 6'h26; // @[Switch.scala 30:53:@12351.4]
  assign valid_38_35 = io_inValid_35 & _T_32389; // @[Switch.scala 30:36:@12352.4]
  assign _T_32392 = io_inAddr_36 == 6'h26; // @[Switch.scala 30:53:@12354.4]
  assign valid_38_36 = io_inValid_36 & _T_32392; // @[Switch.scala 30:36:@12355.4]
  assign _T_32395 = io_inAddr_37 == 6'h26; // @[Switch.scala 30:53:@12357.4]
  assign valid_38_37 = io_inValid_37 & _T_32395; // @[Switch.scala 30:36:@12358.4]
  assign _T_32398 = io_inAddr_38 == 6'h26; // @[Switch.scala 30:53:@12360.4]
  assign valid_38_38 = io_inValid_38 & _T_32398; // @[Switch.scala 30:36:@12361.4]
  assign _T_32401 = io_inAddr_39 == 6'h26; // @[Switch.scala 30:53:@12363.4]
  assign valid_38_39 = io_inValid_39 & _T_32401; // @[Switch.scala 30:36:@12364.4]
  assign _T_32404 = io_inAddr_40 == 6'h26; // @[Switch.scala 30:53:@12366.4]
  assign valid_38_40 = io_inValid_40 & _T_32404; // @[Switch.scala 30:36:@12367.4]
  assign _T_32407 = io_inAddr_41 == 6'h26; // @[Switch.scala 30:53:@12369.4]
  assign valid_38_41 = io_inValid_41 & _T_32407; // @[Switch.scala 30:36:@12370.4]
  assign _T_32410 = io_inAddr_42 == 6'h26; // @[Switch.scala 30:53:@12372.4]
  assign valid_38_42 = io_inValid_42 & _T_32410; // @[Switch.scala 30:36:@12373.4]
  assign _T_32413 = io_inAddr_43 == 6'h26; // @[Switch.scala 30:53:@12375.4]
  assign valid_38_43 = io_inValid_43 & _T_32413; // @[Switch.scala 30:36:@12376.4]
  assign _T_32416 = io_inAddr_44 == 6'h26; // @[Switch.scala 30:53:@12378.4]
  assign valid_38_44 = io_inValid_44 & _T_32416; // @[Switch.scala 30:36:@12379.4]
  assign _T_32419 = io_inAddr_45 == 6'h26; // @[Switch.scala 30:53:@12381.4]
  assign valid_38_45 = io_inValid_45 & _T_32419; // @[Switch.scala 30:36:@12382.4]
  assign _T_32422 = io_inAddr_46 == 6'h26; // @[Switch.scala 30:53:@12384.4]
  assign valid_38_46 = io_inValid_46 & _T_32422; // @[Switch.scala 30:36:@12385.4]
  assign _T_32425 = io_inAddr_47 == 6'h26; // @[Switch.scala 30:53:@12387.4]
  assign valid_38_47 = io_inValid_47 & _T_32425; // @[Switch.scala 30:36:@12388.4]
  assign _T_32428 = io_inAddr_48 == 6'h26; // @[Switch.scala 30:53:@12390.4]
  assign valid_38_48 = io_inValid_48 & _T_32428; // @[Switch.scala 30:36:@12391.4]
  assign _T_32431 = io_inAddr_49 == 6'h26; // @[Switch.scala 30:53:@12393.4]
  assign valid_38_49 = io_inValid_49 & _T_32431; // @[Switch.scala 30:36:@12394.4]
  assign _T_32434 = io_inAddr_50 == 6'h26; // @[Switch.scala 30:53:@12396.4]
  assign valid_38_50 = io_inValid_50 & _T_32434; // @[Switch.scala 30:36:@12397.4]
  assign _T_32437 = io_inAddr_51 == 6'h26; // @[Switch.scala 30:53:@12399.4]
  assign valid_38_51 = io_inValid_51 & _T_32437; // @[Switch.scala 30:36:@12400.4]
  assign _T_32440 = io_inAddr_52 == 6'h26; // @[Switch.scala 30:53:@12402.4]
  assign valid_38_52 = io_inValid_52 & _T_32440; // @[Switch.scala 30:36:@12403.4]
  assign _T_32443 = io_inAddr_53 == 6'h26; // @[Switch.scala 30:53:@12405.4]
  assign valid_38_53 = io_inValid_53 & _T_32443; // @[Switch.scala 30:36:@12406.4]
  assign _T_32446 = io_inAddr_54 == 6'h26; // @[Switch.scala 30:53:@12408.4]
  assign valid_38_54 = io_inValid_54 & _T_32446; // @[Switch.scala 30:36:@12409.4]
  assign _T_32449 = io_inAddr_55 == 6'h26; // @[Switch.scala 30:53:@12411.4]
  assign valid_38_55 = io_inValid_55 & _T_32449; // @[Switch.scala 30:36:@12412.4]
  assign _T_32452 = io_inAddr_56 == 6'h26; // @[Switch.scala 30:53:@12414.4]
  assign valid_38_56 = io_inValid_56 & _T_32452; // @[Switch.scala 30:36:@12415.4]
  assign _T_32455 = io_inAddr_57 == 6'h26; // @[Switch.scala 30:53:@12417.4]
  assign valid_38_57 = io_inValid_57 & _T_32455; // @[Switch.scala 30:36:@12418.4]
  assign _T_32458 = io_inAddr_58 == 6'h26; // @[Switch.scala 30:53:@12420.4]
  assign valid_38_58 = io_inValid_58 & _T_32458; // @[Switch.scala 30:36:@12421.4]
  assign _T_32461 = io_inAddr_59 == 6'h26; // @[Switch.scala 30:53:@12423.4]
  assign valid_38_59 = io_inValid_59 & _T_32461; // @[Switch.scala 30:36:@12424.4]
  assign _T_32464 = io_inAddr_60 == 6'h26; // @[Switch.scala 30:53:@12426.4]
  assign valid_38_60 = io_inValid_60 & _T_32464; // @[Switch.scala 30:36:@12427.4]
  assign _T_32467 = io_inAddr_61 == 6'h26; // @[Switch.scala 30:53:@12429.4]
  assign valid_38_61 = io_inValid_61 & _T_32467; // @[Switch.scala 30:36:@12430.4]
  assign _T_32470 = io_inAddr_62 == 6'h26; // @[Switch.scala 30:53:@12432.4]
  assign valid_38_62 = io_inValid_62 & _T_32470; // @[Switch.scala 30:36:@12433.4]
  assign _T_32473 = io_inAddr_63 == 6'h26; // @[Switch.scala 30:53:@12435.4]
  assign valid_38_63 = io_inValid_63 & _T_32473; // @[Switch.scala 30:36:@12436.4]
  assign _T_32539 = valid_38_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@12438.4]
  assign _T_32540 = valid_38_61 ? 6'h3d : _T_32539; // @[Mux.scala 31:69:@12439.4]
  assign _T_32541 = valid_38_60 ? 6'h3c : _T_32540; // @[Mux.scala 31:69:@12440.4]
  assign _T_32542 = valid_38_59 ? 6'h3b : _T_32541; // @[Mux.scala 31:69:@12441.4]
  assign _T_32543 = valid_38_58 ? 6'h3a : _T_32542; // @[Mux.scala 31:69:@12442.4]
  assign _T_32544 = valid_38_57 ? 6'h39 : _T_32543; // @[Mux.scala 31:69:@12443.4]
  assign _T_32545 = valid_38_56 ? 6'h38 : _T_32544; // @[Mux.scala 31:69:@12444.4]
  assign _T_32546 = valid_38_55 ? 6'h37 : _T_32545; // @[Mux.scala 31:69:@12445.4]
  assign _T_32547 = valid_38_54 ? 6'h36 : _T_32546; // @[Mux.scala 31:69:@12446.4]
  assign _T_32548 = valid_38_53 ? 6'h35 : _T_32547; // @[Mux.scala 31:69:@12447.4]
  assign _T_32549 = valid_38_52 ? 6'h34 : _T_32548; // @[Mux.scala 31:69:@12448.4]
  assign _T_32550 = valid_38_51 ? 6'h33 : _T_32549; // @[Mux.scala 31:69:@12449.4]
  assign _T_32551 = valid_38_50 ? 6'h32 : _T_32550; // @[Mux.scala 31:69:@12450.4]
  assign _T_32552 = valid_38_49 ? 6'h31 : _T_32551; // @[Mux.scala 31:69:@12451.4]
  assign _T_32553 = valid_38_48 ? 6'h30 : _T_32552; // @[Mux.scala 31:69:@12452.4]
  assign _T_32554 = valid_38_47 ? 6'h2f : _T_32553; // @[Mux.scala 31:69:@12453.4]
  assign _T_32555 = valid_38_46 ? 6'h2e : _T_32554; // @[Mux.scala 31:69:@12454.4]
  assign _T_32556 = valid_38_45 ? 6'h2d : _T_32555; // @[Mux.scala 31:69:@12455.4]
  assign _T_32557 = valid_38_44 ? 6'h2c : _T_32556; // @[Mux.scala 31:69:@12456.4]
  assign _T_32558 = valid_38_43 ? 6'h2b : _T_32557; // @[Mux.scala 31:69:@12457.4]
  assign _T_32559 = valid_38_42 ? 6'h2a : _T_32558; // @[Mux.scala 31:69:@12458.4]
  assign _T_32560 = valid_38_41 ? 6'h29 : _T_32559; // @[Mux.scala 31:69:@12459.4]
  assign _T_32561 = valid_38_40 ? 6'h28 : _T_32560; // @[Mux.scala 31:69:@12460.4]
  assign _T_32562 = valid_38_39 ? 6'h27 : _T_32561; // @[Mux.scala 31:69:@12461.4]
  assign _T_32563 = valid_38_38 ? 6'h26 : _T_32562; // @[Mux.scala 31:69:@12462.4]
  assign _T_32564 = valid_38_37 ? 6'h25 : _T_32563; // @[Mux.scala 31:69:@12463.4]
  assign _T_32565 = valid_38_36 ? 6'h24 : _T_32564; // @[Mux.scala 31:69:@12464.4]
  assign _T_32566 = valid_38_35 ? 6'h23 : _T_32565; // @[Mux.scala 31:69:@12465.4]
  assign _T_32567 = valid_38_34 ? 6'h22 : _T_32566; // @[Mux.scala 31:69:@12466.4]
  assign _T_32568 = valid_38_33 ? 6'h21 : _T_32567; // @[Mux.scala 31:69:@12467.4]
  assign _T_32569 = valid_38_32 ? 6'h20 : _T_32568; // @[Mux.scala 31:69:@12468.4]
  assign _T_32570 = valid_38_31 ? 6'h1f : _T_32569; // @[Mux.scala 31:69:@12469.4]
  assign _T_32571 = valid_38_30 ? 6'h1e : _T_32570; // @[Mux.scala 31:69:@12470.4]
  assign _T_32572 = valid_38_29 ? 6'h1d : _T_32571; // @[Mux.scala 31:69:@12471.4]
  assign _T_32573 = valid_38_28 ? 6'h1c : _T_32572; // @[Mux.scala 31:69:@12472.4]
  assign _T_32574 = valid_38_27 ? 6'h1b : _T_32573; // @[Mux.scala 31:69:@12473.4]
  assign _T_32575 = valid_38_26 ? 6'h1a : _T_32574; // @[Mux.scala 31:69:@12474.4]
  assign _T_32576 = valid_38_25 ? 6'h19 : _T_32575; // @[Mux.scala 31:69:@12475.4]
  assign _T_32577 = valid_38_24 ? 6'h18 : _T_32576; // @[Mux.scala 31:69:@12476.4]
  assign _T_32578 = valid_38_23 ? 6'h17 : _T_32577; // @[Mux.scala 31:69:@12477.4]
  assign _T_32579 = valid_38_22 ? 6'h16 : _T_32578; // @[Mux.scala 31:69:@12478.4]
  assign _T_32580 = valid_38_21 ? 6'h15 : _T_32579; // @[Mux.scala 31:69:@12479.4]
  assign _T_32581 = valid_38_20 ? 6'h14 : _T_32580; // @[Mux.scala 31:69:@12480.4]
  assign _T_32582 = valid_38_19 ? 6'h13 : _T_32581; // @[Mux.scala 31:69:@12481.4]
  assign _T_32583 = valid_38_18 ? 6'h12 : _T_32582; // @[Mux.scala 31:69:@12482.4]
  assign _T_32584 = valid_38_17 ? 6'h11 : _T_32583; // @[Mux.scala 31:69:@12483.4]
  assign _T_32585 = valid_38_16 ? 6'h10 : _T_32584; // @[Mux.scala 31:69:@12484.4]
  assign _T_32586 = valid_38_15 ? 6'hf : _T_32585; // @[Mux.scala 31:69:@12485.4]
  assign _T_32587 = valid_38_14 ? 6'he : _T_32586; // @[Mux.scala 31:69:@12486.4]
  assign _T_32588 = valid_38_13 ? 6'hd : _T_32587; // @[Mux.scala 31:69:@12487.4]
  assign _T_32589 = valid_38_12 ? 6'hc : _T_32588; // @[Mux.scala 31:69:@12488.4]
  assign _T_32590 = valid_38_11 ? 6'hb : _T_32589; // @[Mux.scala 31:69:@12489.4]
  assign _T_32591 = valid_38_10 ? 6'ha : _T_32590; // @[Mux.scala 31:69:@12490.4]
  assign _T_32592 = valid_38_9 ? 6'h9 : _T_32591; // @[Mux.scala 31:69:@12491.4]
  assign _T_32593 = valid_38_8 ? 6'h8 : _T_32592; // @[Mux.scala 31:69:@12492.4]
  assign _T_32594 = valid_38_7 ? 6'h7 : _T_32593; // @[Mux.scala 31:69:@12493.4]
  assign _T_32595 = valid_38_6 ? 6'h6 : _T_32594; // @[Mux.scala 31:69:@12494.4]
  assign _T_32596 = valid_38_5 ? 6'h5 : _T_32595; // @[Mux.scala 31:69:@12495.4]
  assign _T_32597 = valid_38_4 ? 6'h4 : _T_32596; // @[Mux.scala 31:69:@12496.4]
  assign _T_32598 = valid_38_3 ? 6'h3 : _T_32597; // @[Mux.scala 31:69:@12497.4]
  assign _T_32599 = valid_38_2 ? 6'h2 : _T_32598; // @[Mux.scala 31:69:@12498.4]
  assign _T_32600 = valid_38_1 ? 6'h1 : _T_32599; // @[Mux.scala 31:69:@12499.4]
  assign select_38 = valid_38_0 ? 6'h0 : _T_32600; // @[Mux.scala 31:69:@12500.4]
  assign _GEN_2433 = 6'h1 == select_38 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2434 = 6'h2 == select_38 ? io_inData_2 : _GEN_2433; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2435 = 6'h3 == select_38 ? io_inData_3 : _GEN_2434; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2436 = 6'h4 == select_38 ? io_inData_4 : _GEN_2435; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2437 = 6'h5 == select_38 ? io_inData_5 : _GEN_2436; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2438 = 6'h6 == select_38 ? io_inData_6 : _GEN_2437; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2439 = 6'h7 == select_38 ? io_inData_7 : _GEN_2438; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2440 = 6'h8 == select_38 ? io_inData_8 : _GEN_2439; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2441 = 6'h9 == select_38 ? io_inData_9 : _GEN_2440; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2442 = 6'ha == select_38 ? io_inData_10 : _GEN_2441; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2443 = 6'hb == select_38 ? io_inData_11 : _GEN_2442; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2444 = 6'hc == select_38 ? io_inData_12 : _GEN_2443; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2445 = 6'hd == select_38 ? io_inData_13 : _GEN_2444; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2446 = 6'he == select_38 ? io_inData_14 : _GEN_2445; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2447 = 6'hf == select_38 ? io_inData_15 : _GEN_2446; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2448 = 6'h10 == select_38 ? io_inData_16 : _GEN_2447; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2449 = 6'h11 == select_38 ? io_inData_17 : _GEN_2448; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2450 = 6'h12 == select_38 ? io_inData_18 : _GEN_2449; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2451 = 6'h13 == select_38 ? io_inData_19 : _GEN_2450; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2452 = 6'h14 == select_38 ? io_inData_20 : _GEN_2451; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2453 = 6'h15 == select_38 ? io_inData_21 : _GEN_2452; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2454 = 6'h16 == select_38 ? io_inData_22 : _GEN_2453; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2455 = 6'h17 == select_38 ? io_inData_23 : _GEN_2454; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2456 = 6'h18 == select_38 ? io_inData_24 : _GEN_2455; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2457 = 6'h19 == select_38 ? io_inData_25 : _GEN_2456; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2458 = 6'h1a == select_38 ? io_inData_26 : _GEN_2457; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2459 = 6'h1b == select_38 ? io_inData_27 : _GEN_2458; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2460 = 6'h1c == select_38 ? io_inData_28 : _GEN_2459; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2461 = 6'h1d == select_38 ? io_inData_29 : _GEN_2460; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2462 = 6'h1e == select_38 ? io_inData_30 : _GEN_2461; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2463 = 6'h1f == select_38 ? io_inData_31 : _GEN_2462; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2464 = 6'h20 == select_38 ? io_inData_32 : _GEN_2463; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2465 = 6'h21 == select_38 ? io_inData_33 : _GEN_2464; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2466 = 6'h22 == select_38 ? io_inData_34 : _GEN_2465; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2467 = 6'h23 == select_38 ? io_inData_35 : _GEN_2466; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2468 = 6'h24 == select_38 ? io_inData_36 : _GEN_2467; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2469 = 6'h25 == select_38 ? io_inData_37 : _GEN_2468; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2470 = 6'h26 == select_38 ? io_inData_38 : _GEN_2469; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2471 = 6'h27 == select_38 ? io_inData_39 : _GEN_2470; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2472 = 6'h28 == select_38 ? io_inData_40 : _GEN_2471; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2473 = 6'h29 == select_38 ? io_inData_41 : _GEN_2472; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2474 = 6'h2a == select_38 ? io_inData_42 : _GEN_2473; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2475 = 6'h2b == select_38 ? io_inData_43 : _GEN_2474; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2476 = 6'h2c == select_38 ? io_inData_44 : _GEN_2475; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2477 = 6'h2d == select_38 ? io_inData_45 : _GEN_2476; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2478 = 6'h2e == select_38 ? io_inData_46 : _GEN_2477; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2479 = 6'h2f == select_38 ? io_inData_47 : _GEN_2478; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2480 = 6'h30 == select_38 ? io_inData_48 : _GEN_2479; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2481 = 6'h31 == select_38 ? io_inData_49 : _GEN_2480; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2482 = 6'h32 == select_38 ? io_inData_50 : _GEN_2481; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2483 = 6'h33 == select_38 ? io_inData_51 : _GEN_2482; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2484 = 6'h34 == select_38 ? io_inData_52 : _GEN_2483; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2485 = 6'h35 == select_38 ? io_inData_53 : _GEN_2484; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2486 = 6'h36 == select_38 ? io_inData_54 : _GEN_2485; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2487 = 6'h37 == select_38 ? io_inData_55 : _GEN_2486; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2488 = 6'h38 == select_38 ? io_inData_56 : _GEN_2487; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2489 = 6'h39 == select_38 ? io_inData_57 : _GEN_2488; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2490 = 6'h3a == select_38 ? io_inData_58 : _GEN_2489; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2491 = 6'h3b == select_38 ? io_inData_59 : _GEN_2490; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2492 = 6'h3c == select_38 ? io_inData_60 : _GEN_2491; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2493 = 6'h3d == select_38 ? io_inData_61 : _GEN_2492; // @[Switch.scala 33:19:@12502.4]
  assign _GEN_2494 = 6'h3e == select_38 ? io_inData_62 : _GEN_2493; // @[Switch.scala 33:19:@12502.4]
  assign _T_32609 = {valid_38_7,valid_38_6,valid_38_5,valid_38_4,valid_38_3,valid_38_2,valid_38_1,valid_38_0}; // @[Switch.scala 34:32:@12509.4]
  assign _T_32617 = {valid_38_15,valid_38_14,valid_38_13,valid_38_12,valid_38_11,valid_38_10,valid_38_9,valid_38_8,_T_32609}; // @[Switch.scala 34:32:@12517.4]
  assign _T_32624 = {valid_38_23,valid_38_22,valid_38_21,valid_38_20,valid_38_19,valid_38_18,valid_38_17,valid_38_16}; // @[Switch.scala 34:32:@12524.4]
  assign _T_32633 = {valid_38_31,valid_38_30,valid_38_29,valid_38_28,valid_38_27,valid_38_26,valid_38_25,valid_38_24,_T_32624,_T_32617}; // @[Switch.scala 34:32:@12533.4]
  assign _T_32640 = {valid_38_39,valid_38_38,valid_38_37,valid_38_36,valid_38_35,valid_38_34,valid_38_33,valid_38_32}; // @[Switch.scala 34:32:@12540.4]
  assign _T_32648 = {valid_38_47,valid_38_46,valid_38_45,valid_38_44,valid_38_43,valid_38_42,valid_38_41,valid_38_40,_T_32640}; // @[Switch.scala 34:32:@12548.4]
  assign _T_32655 = {valid_38_55,valid_38_54,valid_38_53,valid_38_52,valid_38_51,valid_38_50,valid_38_49,valid_38_48}; // @[Switch.scala 34:32:@12555.4]
  assign _T_32664 = {valid_38_63,valid_38_62,valid_38_61,valid_38_60,valid_38_59,valid_38_58,valid_38_57,valid_38_56,_T_32655,_T_32648}; // @[Switch.scala 34:32:@12564.4]
  assign _T_32665 = {_T_32664,_T_32633}; // @[Switch.scala 34:32:@12565.4]
  assign _T_32669 = io_inAddr_0 == 6'h27; // @[Switch.scala 30:53:@12568.4]
  assign valid_39_0 = io_inValid_0 & _T_32669; // @[Switch.scala 30:36:@12569.4]
  assign _T_32672 = io_inAddr_1 == 6'h27; // @[Switch.scala 30:53:@12571.4]
  assign valid_39_1 = io_inValid_1 & _T_32672; // @[Switch.scala 30:36:@12572.4]
  assign _T_32675 = io_inAddr_2 == 6'h27; // @[Switch.scala 30:53:@12574.4]
  assign valid_39_2 = io_inValid_2 & _T_32675; // @[Switch.scala 30:36:@12575.4]
  assign _T_32678 = io_inAddr_3 == 6'h27; // @[Switch.scala 30:53:@12577.4]
  assign valid_39_3 = io_inValid_3 & _T_32678; // @[Switch.scala 30:36:@12578.4]
  assign _T_32681 = io_inAddr_4 == 6'h27; // @[Switch.scala 30:53:@12580.4]
  assign valid_39_4 = io_inValid_4 & _T_32681; // @[Switch.scala 30:36:@12581.4]
  assign _T_32684 = io_inAddr_5 == 6'h27; // @[Switch.scala 30:53:@12583.4]
  assign valid_39_5 = io_inValid_5 & _T_32684; // @[Switch.scala 30:36:@12584.4]
  assign _T_32687 = io_inAddr_6 == 6'h27; // @[Switch.scala 30:53:@12586.4]
  assign valid_39_6 = io_inValid_6 & _T_32687; // @[Switch.scala 30:36:@12587.4]
  assign _T_32690 = io_inAddr_7 == 6'h27; // @[Switch.scala 30:53:@12589.4]
  assign valid_39_7 = io_inValid_7 & _T_32690; // @[Switch.scala 30:36:@12590.4]
  assign _T_32693 = io_inAddr_8 == 6'h27; // @[Switch.scala 30:53:@12592.4]
  assign valid_39_8 = io_inValid_8 & _T_32693; // @[Switch.scala 30:36:@12593.4]
  assign _T_32696 = io_inAddr_9 == 6'h27; // @[Switch.scala 30:53:@12595.4]
  assign valid_39_9 = io_inValid_9 & _T_32696; // @[Switch.scala 30:36:@12596.4]
  assign _T_32699 = io_inAddr_10 == 6'h27; // @[Switch.scala 30:53:@12598.4]
  assign valid_39_10 = io_inValid_10 & _T_32699; // @[Switch.scala 30:36:@12599.4]
  assign _T_32702 = io_inAddr_11 == 6'h27; // @[Switch.scala 30:53:@12601.4]
  assign valid_39_11 = io_inValid_11 & _T_32702; // @[Switch.scala 30:36:@12602.4]
  assign _T_32705 = io_inAddr_12 == 6'h27; // @[Switch.scala 30:53:@12604.4]
  assign valid_39_12 = io_inValid_12 & _T_32705; // @[Switch.scala 30:36:@12605.4]
  assign _T_32708 = io_inAddr_13 == 6'h27; // @[Switch.scala 30:53:@12607.4]
  assign valid_39_13 = io_inValid_13 & _T_32708; // @[Switch.scala 30:36:@12608.4]
  assign _T_32711 = io_inAddr_14 == 6'h27; // @[Switch.scala 30:53:@12610.4]
  assign valid_39_14 = io_inValid_14 & _T_32711; // @[Switch.scala 30:36:@12611.4]
  assign _T_32714 = io_inAddr_15 == 6'h27; // @[Switch.scala 30:53:@12613.4]
  assign valid_39_15 = io_inValid_15 & _T_32714; // @[Switch.scala 30:36:@12614.4]
  assign _T_32717 = io_inAddr_16 == 6'h27; // @[Switch.scala 30:53:@12616.4]
  assign valid_39_16 = io_inValid_16 & _T_32717; // @[Switch.scala 30:36:@12617.4]
  assign _T_32720 = io_inAddr_17 == 6'h27; // @[Switch.scala 30:53:@12619.4]
  assign valid_39_17 = io_inValid_17 & _T_32720; // @[Switch.scala 30:36:@12620.4]
  assign _T_32723 = io_inAddr_18 == 6'h27; // @[Switch.scala 30:53:@12622.4]
  assign valid_39_18 = io_inValid_18 & _T_32723; // @[Switch.scala 30:36:@12623.4]
  assign _T_32726 = io_inAddr_19 == 6'h27; // @[Switch.scala 30:53:@12625.4]
  assign valid_39_19 = io_inValid_19 & _T_32726; // @[Switch.scala 30:36:@12626.4]
  assign _T_32729 = io_inAddr_20 == 6'h27; // @[Switch.scala 30:53:@12628.4]
  assign valid_39_20 = io_inValid_20 & _T_32729; // @[Switch.scala 30:36:@12629.4]
  assign _T_32732 = io_inAddr_21 == 6'h27; // @[Switch.scala 30:53:@12631.4]
  assign valid_39_21 = io_inValid_21 & _T_32732; // @[Switch.scala 30:36:@12632.4]
  assign _T_32735 = io_inAddr_22 == 6'h27; // @[Switch.scala 30:53:@12634.4]
  assign valid_39_22 = io_inValid_22 & _T_32735; // @[Switch.scala 30:36:@12635.4]
  assign _T_32738 = io_inAddr_23 == 6'h27; // @[Switch.scala 30:53:@12637.4]
  assign valid_39_23 = io_inValid_23 & _T_32738; // @[Switch.scala 30:36:@12638.4]
  assign _T_32741 = io_inAddr_24 == 6'h27; // @[Switch.scala 30:53:@12640.4]
  assign valid_39_24 = io_inValid_24 & _T_32741; // @[Switch.scala 30:36:@12641.4]
  assign _T_32744 = io_inAddr_25 == 6'h27; // @[Switch.scala 30:53:@12643.4]
  assign valid_39_25 = io_inValid_25 & _T_32744; // @[Switch.scala 30:36:@12644.4]
  assign _T_32747 = io_inAddr_26 == 6'h27; // @[Switch.scala 30:53:@12646.4]
  assign valid_39_26 = io_inValid_26 & _T_32747; // @[Switch.scala 30:36:@12647.4]
  assign _T_32750 = io_inAddr_27 == 6'h27; // @[Switch.scala 30:53:@12649.4]
  assign valid_39_27 = io_inValid_27 & _T_32750; // @[Switch.scala 30:36:@12650.4]
  assign _T_32753 = io_inAddr_28 == 6'h27; // @[Switch.scala 30:53:@12652.4]
  assign valid_39_28 = io_inValid_28 & _T_32753; // @[Switch.scala 30:36:@12653.4]
  assign _T_32756 = io_inAddr_29 == 6'h27; // @[Switch.scala 30:53:@12655.4]
  assign valid_39_29 = io_inValid_29 & _T_32756; // @[Switch.scala 30:36:@12656.4]
  assign _T_32759 = io_inAddr_30 == 6'h27; // @[Switch.scala 30:53:@12658.4]
  assign valid_39_30 = io_inValid_30 & _T_32759; // @[Switch.scala 30:36:@12659.4]
  assign _T_32762 = io_inAddr_31 == 6'h27; // @[Switch.scala 30:53:@12661.4]
  assign valid_39_31 = io_inValid_31 & _T_32762; // @[Switch.scala 30:36:@12662.4]
  assign _T_32765 = io_inAddr_32 == 6'h27; // @[Switch.scala 30:53:@12664.4]
  assign valid_39_32 = io_inValid_32 & _T_32765; // @[Switch.scala 30:36:@12665.4]
  assign _T_32768 = io_inAddr_33 == 6'h27; // @[Switch.scala 30:53:@12667.4]
  assign valid_39_33 = io_inValid_33 & _T_32768; // @[Switch.scala 30:36:@12668.4]
  assign _T_32771 = io_inAddr_34 == 6'h27; // @[Switch.scala 30:53:@12670.4]
  assign valid_39_34 = io_inValid_34 & _T_32771; // @[Switch.scala 30:36:@12671.4]
  assign _T_32774 = io_inAddr_35 == 6'h27; // @[Switch.scala 30:53:@12673.4]
  assign valid_39_35 = io_inValid_35 & _T_32774; // @[Switch.scala 30:36:@12674.4]
  assign _T_32777 = io_inAddr_36 == 6'h27; // @[Switch.scala 30:53:@12676.4]
  assign valid_39_36 = io_inValid_36 & _T_32777; // @[Switch.scala 30:36:@12677.4]
  assign _T_32780 = io_inAddr_37 == 6'h27; // @[Switch.scala 30:53:@12679.4]
  assign valid_39_37 = io_inValid_37 & _T_32780; // @[Switch.scala 30:36:@12680.4]
  assign _T_32783 = io_inAddr_38 == 6'h27; // @[Switch.scala 30:53:@12682.4]
  assign valid_39_38 = io_inValid_38 & _T_32783; // @[Switch.scala 30:36:@12683.4]
  assign _T_32786 = io_inAddr_39 == 6'h27; // @[Switch.scala 30:53:@12685.4]
  assign valid_39_39 = io_inValid_39 & _T_32786; // @[Switch.scala 30:36:@12686.4]
  assign _T_32789 = io_inAddr_40 == 6'h27; // @[Switch.scala 30:53:@12688.4]
  assign valid_39_40 = io_inValid_40 & _T_32789; // @[Switch.scala 30:36:@12689.4]
  assign _T_32792 = io_inAddr_41 == 6'h27; // @[Switch.scala 30:53:@12691.4]
  assign valid_39_41 = io_inValid_41 & _T_32792; // @[Switch.scala 30:36:@12692.4]
  assign _T_32795 = io_inAddr_42 == 6'h27; // @[Switch.scala 30:53:@12694.4]
  assign valid_39_42 = io_inValid_42 & _T_32795; // @[Switch.scala 30:36:@12695.4]
  assign _T_32798 = io_inAddr_43 == 6'h27; // @[Switch.scala 30:53:@12697.4]
  assign valid_39_43 = io_inValid_43 & _T_32798; // @[Switch.scala 30:36:@12698.4]
  assign _T_32801 = io_inAddr_44 == 6'h27; // @[Switch.scala 30:53:@12700.4]
  assign valid_39_44 = io_inValid_44 & _T_32801; // @[Switch.scala 30:36:@12701.4]
  assign _T_32804 = io_inAddr_45 == 6'h27; // @[Switch.scala 30:53:@12703.4]
  assign valid_39_45 = io_inValid_45 & _T_32804; // @[Switch.scala 30:36:@12704.4]
  assign _T_32807 = io_inAddr_46 == 6'h27; // @[Switch.scala 30:53:@12706.4]
  assign valid_39_46 = io_inValid_46 & _T_32807; // @[Switch.scala 30:36:@12707.4]
  assign _T_32810 = io_inAddr_47 == 6'h27; // @[Switch.scala 30:53:@12709.4]
  assign valid_39_47 = io_inValid_47 & _T_32810; // @[Switch.scala 30:36:@12710.4]
  assign _T_32813 = io_inAddr_48 == 6'h27; // @[Switch.scala 30:53:@12712.4]
  assign valid_39_48 = io_inValid_48 & _T_32813; // @[Switch.scala 30:36:@12713.4]
  assign _T_32816 = io_inAddr_49 == 6'h27; // @[Switch.scala 30:53:@12715.4]
  assign valid_39_49 = io_inValid_49 & _T_32816; // @[Switch.scala 30:36:@12716.4]
  assign _T_32819 = io_inAddr_50 == 6'h27; // @[Switch.scala 30:53:@12718.4]
  assign valid_39_50 = io_inValid_50 & _T_32819; // @[Switch.scala 30:36:@12719.4]
  assign _T_32822 = io_inAddr_51 == 6'h27; // @[Switch.scala 30:53:@12721.4]
  assign valid_39_51 = io_inValid_51 & _T_32822; // @[Switch.scala 30:36:@12722.4]
  assign _T_32825 = io_inAddr_52 == 6'h27; // @[Switch.scala 30:53:@12724.4]
  assign valid_39_52 = io_inValid_52 & _T_32825; // @[Switch.scala 30:36:@12725.4]
  assign _T_32828 = io_inAddr_53 == 6'h27; // @[Switch.scala 30:53:@12727.4]
  assign valid_39_53 = io_inValid_53 & _T_32828; // @[Switch.scala 30:36:@12728.4]
  assign _T_32831 = io_inAddr_54 == 6'h27; // @[Switch.scala 30:53:@12730.4]
  assign valid_39_54 = io_inValid_54 & _T_32831; // @[Switch.scala 30:36:@12731.4]
  assign _T_32834 = io_inAddr_55 == 6'h27; // @[Switch.scala 30:53:@12733.4]
  assign valid_39_55 = io_inValid_55 & _T_32834; // @[Switch.scala 30:36:@12734.4]
  assign _T_32837 = io_inAddr_56 == 6'h27; // @[Switch.scala 30:53:@12736.4]
  assign valid_39_56 = io_inValid_56 & _T_32837; // @[Switch.scala 30:36:@12737.4]
  assign _T_32840 = io_inAddr_57 == 6'h27; // @[Switch.scala 30:53:@12739.4]
  assign valid_39_57 = io_inValid_57 & _T_32840; // @[Switch.scala 30:36:@12740.4]
  assign _T_32843 = io_inAddr_58 == 6'h27; // @[Switch.scala 30:53:@12742.4]
  assign valid_39_58 = io_inValid_58 & _T_32843; // @[Switch.scala 30:36:@12743.4]
  assign _T_32846 = io_inAddr_59 == 6'h27; // @[Switch.scala 30:53:@12745.4]
  assign valid_39_59 = io_inValid_59 & _T_32846; // @[Switch.scala 30:36:@12746.4]
  assign _T_32849 = io_inAddr_60 == 6'h27; // @[Switch.scala 30:53:@12748.4]
  assign valid_39_60 = io_inValid_60 & _T_32849; // @[Switch.scala 30:36:@12749.4]
  assign _T_32852 = io_inAddr_61 == 6'h27; // @[Switch.scala 30:53:@12751.4]
  assign valid_39_61 = io_inValid_61 & _T_32852; // @[Switch.scala 30:36:@12752.4]
  assign _T_32855 = io_inAddr_62 == 6'h27; // @[Switch.scala 30:53:@12754.4]
  assign valid_39_62 = io_inValid_62 & _T_32855; // @[Switch.scala 30:36:@12755.4]
  assign _T_32858 = io_inAddr_63 == 6'h27; // @[Switch.scala 30:53:@12757.4]
  assign valid_39_63 = io_inValid_63 & _T_32858; // @[Switch.scala 30:36:@12758.4]
  assign _T_32924 = valid_39_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@12760.4]
  assign _T_32925 = valid_39_61 ? 6'h3d : _T_32924; // @[Mux.scala 31:69:@12761.4]
  assign _T_32926 = valid_39_60 ? 6'h3c : _T_32925; // @[Mux.scala 31:69:@12762.4]
  assign _T_32927 = valid_39_59 ? 6'h3b : _T_32926; // @[Mux.scala 31:69:@12763.4]
  assign _T_32928 = valid_39_58 ? 6'h3a : _T_32927; // @[Mux.scala 31:69:@12764.4]
  assign _T_32929 = valid_39_57 ? 6'h39 : _T_32928; // @[Mux.scala 31:69:@12765.4]
  assign _T_32930 = valid_39_56 ? 6'h38 : _T_32929; // @[Mux.scala 31:69:@12766.4]
  assign _T_32931 = valid_39_55 ? 6'h37 : _T_32930; // @[Mux.scala 31:69:@12767.4]
  assign _T_32932 = valid_39_54 ? 6'h36 : _T_32931; // @[Mux.scala 31:69:@12768.4]
  assign _T_32933 = valid_39_53 ? 6'h35 : _T_32932; // @[Mux.scala 31:69:@12769.4]
  assign _T_32934 = valid_39_52 ? 6'h34 : _T_32933; // @[Mux.scala 31:69:@12770.4]
  assign _T_32935 = valid_39_51 ? 6'h33 : _T_32934; // @[Mux.scala 31:69:@12771.4]
  assign _T_32936 = valid_39_50 ? 6'h32 : _T_32935; // @[Mux.scala 31:69:@12772.4]
  assign _T_32937 = valid_39_49 ? 6'h31 : _T_32936; // @[Mux.scala 31:69:@12773.4]
  assign _T_32938 = valid_39_48 ? 6'h30 : _T_32937; // @[Mux.scala 31:69:@12774.4]
  assign _T_32939 = valid_39_47 ? 6'h2f : _T_32938; // @[Mux.scala 31:69:@12775.4]
  assign _T_32940 = valid_39_46 ? 6'h2e : _T_32939; // @[Mux.scala 31:69:@12776.4]
  assign _T_32941 = valid_39_45 ? 6'h2d : _T_32940; // @[Mux.scala 31:69:@12777.4]
  assign _T_32942 = valid_39_44 ? 6'h2c : _T_32941; // @[Mux.scala 31:69:@12778.4]
  assign _T_32943 = valid_39_43 ? 6'h2b : _T_32942; // @[Mux.scala 31:69:@12779.4]
  assign _T_32944 = valid_39_42 ? 6'h2a : _T_32943; // @[Mux.scala 31:69:@12780.4]
  assign _T_32945 = valid_39_41 ? 6'h29 : _T_32944; // @[Mux.scala 31:69:@12781.4]
  assign _T_32946 = valid_39_40 ? 6'h28 : _T_32945; // @[Mux.scala 31:69:@12782.4]
  assign _T_32947 = valid_39_39 ? 6'h27 : _T_32946; // @[Mux.scala 31:69:@12783.4]
  assign _T_32948 = valid_39_38 ? 6'h26 : _T_32947; // @[Mux.scala 31:69:@12784.4]
  assign _T_32949 = valid_39_37 ? 6'h25 : _T_32948; // @[Mux.scala 31:69:@12785.4]
  assign _T_32950 = valid_39_36 ? 6'h24 : _T_32949; // @[Mux.scala 31:69:@12786.4]
  assign _T_32951 = valid_39_35 ? 6'h23 : _T_32950; // @[Mux.scala 31:69:@12787.4]
  assign _T_32952 = valid_39_34 ? 6'h22 : _T_32951; // @[Mux.scala 31:69:@12788.4]
  assign _T_32953 = valid_39_33 ? 6'h21 : _T_32952; // @[Mux.scala 31:69:@12789.4]
  assign _T_32954 = valid_39_32 ? 6'h20 : _T_32953; // @[Mux.scala 31:69:@12790.4]
  assign _T_32955 = valid_39_31 ? 6'h1f : _T_32954; // @[Mux.scala 31:69:@12791.4]
  assign _T_32956 = valid_39_30 ? 6'h1e : _T_32955; // @[Mux.scala 31:69:@12792.4]
  assign _T_32957 = valid_39_29 ? 6'h1d : _T_32956; // @[Mux.scala 31:69:@12793.4]
  assign _T_32958 = valid_39_28 ? 6'h1c : _T_32957; // @[Mux.scala 31:69:@12794.4]
  assign _T_32959 = valid_39_27 ? 6'h1b : _T_32958; // @[Mux.scala 31:69:@12795.4]
  assign _T_32960 = valid_39_26 ? 6'h1a : _T_32959; // @[Mux.scala 31:69:@12796.4]
  assign _T_32961 = valid_39_25 ? 6'h19 : _T_32960; // @[Mux.scala 31:69:@12797.4]
  assign _T_32962 = valid_39_24 ? 6'h18 : _T_32961; // @[Mux.scala 31:69:@12798.4]
  assign _T_32963 = valid_39_23 ? 6'h17 : _T_32962; // @[Mux.scala 31:69:@12799.4]
  assign _T_32964 = valid_39_22 ? 6'h16 : _T_32963; // @[Mux.scala 31:69:@12800.4]
  assign _T_32965 = valid_39_21 ? 6'h15 : _T_32964; // @[Mux.scala 31:69:@12801.4]
  assign _T_32966 = valid_39_20 ? 6'h14 : _T_32965; // @[Mux.scala 31:69:@12802.4]
  assign _T_32967 = valid_39_19 ? 6'h13 : _T_32966; // @[Mux.scala 31:69:@12803.4]
  assign _T_32968 = valid_39_18 ? 6'h12 : _T_32967; // @[Mux.scala 31:69:@12804.4]
  assign _T_32969 = valid_39_17 ? 6'h11 : _T_32968; // @[Mux.scala 31:69:@12805.4]
  assign _T_32970 = valid_39_16 ? 6'h10 : _T_32969; // @[Mux.scala 31:69:@12806.4]
  assign _T_32971 = valid_39_15 ? 6'hf : _T_32970; // @[Mux.scala 31:69:@12807.4]
  assign _T_32972 = valid_39_14 ? 6'he : _T_32971; // @[Mux.scala 31:69:@12808.4]
  assign _T_32973 = valid_39_13 ? 6'hd : _T_32972; // @[Mux.scala 31:69:@12809.4]
  assign _T_32974 = valid_39_12 ? 6'hc : _T_32973; // @[Mux.scala 31:69:@12810.4]
  assign _T_32975 = valid_39_11 ? 6'hb : _T_32974; // @[Mux.scala 31:69:@12811.4]
  assign _T_32976 = valid_39_10 ? 6'ha : _T_32975; // @[Mux.scala 31:69:@12812.4]
  assign _T_32977 = valid_39_9 ? 6'h9 : _T_32976; // @[Mux.scala 31:69:@12813.4]
  assign _T_32978 = valid_39_8 ? 6'h8 : _T_32977; // @[Mux.scala 31:69:@12814.4]
  assign _T_32979 = valid_39_7 ? 6'h7 : _T_32978; // @[Mux.scala 31:69:@12815.4]
  assign _T_32980 = valid_39_6 ? 6'h6 : _T_32979; // @[Mux.scala 31:69:@12816.4]
  assign _T_32981 = valid_39_5 ? 6'h5 : _T_32980; // @[Mux.scala 31:69:@12817.4]
  assign _T_32982 = valid_39_4 ? 6'h4 : _T_32981; // @[Mux.scala 31:69:@12818.4]
  assign _T_32983 = valid_39_3 ? 6'h3 : _T_32982; // @[Mux.scala 31:69:@12819.4]
  assign _T_32984 = valid_39_2 ? 6'h2 : _T_32983; // @[Mux.scala 31:69:@12820.4]
  assign _T_32985 = valid_39_1 ? 6'h1 : _T_32984; // @[Mux.scala 31:69:@12821.4]
  assign select_39 = valid_39_0 ? 6'h0 : _T_32985; // @[Mux.scala 31:69:@12822.4]
  assign _GEN_2497 = 6'h1 == select_39 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2498 = 6'h2 == select_39 ? io_inData_2 : _GEN_2497; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2499 = 6'h3 == select_39 ? io_inData_3 : _GEN_2498; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2500 = 6'h4 == select_39 ? io_inData_4 : _GEN_2499; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2501 = 6'h5 == select_39 ? io_inData_5 : _GEN_2500; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2502 = 6'h6 == select_39 ? io_inData_6 : _GEN_2501; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2503 = 6'h7 == select_39 ? io_inData_7 : _GEN_2502; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2504 = 6'h8 == select_39 ? io_inData_8 : _GEN_2503; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2505 = 6'h9 == select_39 ? io_inData_9 : _GEN_2504; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2506 = 6'ha == select_39 ? io_inData_10 : _GEN_2505; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2507 = 6'hb == select_39 ? io_inData_11 : _GEN_2506; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2508 = 6'hc == select_39 ? io_inData_12 : _GEN_2507; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2509 = 6'hd == select_39 ? io_inData_13 : _GEN_2508; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2510 = 6'he == select_39 ? io_inData_14 : _GEN_2509; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2511 = 6'hf == select_39 ? io_inData_15 : _GEN_2510; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2512 = 6'h10 == select_39 ? io_inData_16 : _GEN_2511; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2513 = 6'h11 == select_39 ? io_inData_17 : _GEN_2512; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2514 = 6'h12 == select_39 ? io_inData_18 : _GEN_2513; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2515 = 6'h13 == select_39 ? io_inData_19 : _GEN_2514; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2516 = 6'h14 == select_39 ? io_inData_20 : _GEN_2515; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2517 = 6'h15 == select_39 ? io_inData_21 : _GEN_2516; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2518 = 6'h16 == select_39 ? io_inData_22 : _GEN_2517; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2519 = 6'h17 == select_39 ? io_inData_23 : _GEN_2518; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2520 = 6'h18 == select_39 ? io_inData_24 : _GEN_2519; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2521 = 6'h19 == select_39 ? io_inData_25 : _GEN_2520; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2522 = 6'h1a == select_39 ? io_inData_26 : _GEN_2521; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2523 = 6'h1b == select_39 ? io_inData_27 : _GEN_2522; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2524 = 6'h1c == select_39 ? io_inData_28 : _GEN_2523; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2525 = 6'h1d == select_39 ? io_inData_29 : _GEN_2524; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2526 = 6'h1e == select_39 ? io_inData_30 : _GEN_2525; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2527 = 6'h1f == select_39 ? io_inData_31 : _GEN_2526; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2528 = 6'h20 == select_39 ? io_inData_32 : _GEN_2527; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2529 = 6'h21 == select_39 ? io_inData_33 : _GEN_2528; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2530 = 6'h22 == select_39 ? io_inData_34 : _GEN_2529; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2531 = 6'h23 == select_39 ? io_inData_35 : _GEN_2530; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2532 = 6'h24 == select_39 ? io_inData_36 : _GEN_2531; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2533 = 6'h25 == select_39 ? io_inData_37 : _GEN_2532; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2534 = 6'h26 == select_39 ? io_inData_38 : _GEN_2533; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2535 = 6'h27 == select_39 ? io_inData_39 : _GEN_2534; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2536 = 6'h28 == select_39 ? io_inData_40 : _GEN_2535; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2537 = 6'h29 == select_39 ? io_inData_41 : _GEN_2536; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2538 = 6'h2a == select_39 ? io_inData_42 : _GEN_2537; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2539 = 6'h2b == select_39 ? io_inData_43 : _GEN_2538; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2540 = 6'h2c == select_39 ? io_inData_44 : _GEN_2539; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2541 = 6'h2d == select_39 ? io_inData_45 : _GEN_2540; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2542 = 6'h2e == select_39 ? io_inData_46 : _GEN_2541; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2543 = 6'h2f == select_39 ? io_inData_47 : _GEN_2542; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2544 = 6'h30 == select_39 ? io_inData_48 : _GEN_2543; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2545 = 6'h31 == select_39 ? io_inData_49 : _GEN_2544; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2546 = 6'h32 == select_39 ? io_inData_50 : _GEN_2545; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2547 = 6'h33 == select_39 ? io_inData_51 : _GEN_2546; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2548 = 6'h34 == select_39 ? io_inData_52 : _GEN_2547; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2549 = 6'h35 == select_39 ? io_inData_53 : _GEN_2548; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2550 = 6'h36 == select_39 ? io_inData_54 : _GEN_2549; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2551 = 6'h37 == select_39 ? io_inData_55 : _GEN_2550; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2552 = 6'h38 == select_39 ? io_inData_56 : _GEN_2551; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2553 = 6'h39 == select_39 ? io_inData_57 : _GEN_2552; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2554 = 6'h3a == select_39 ? io_inData_58 : _GEN_2553; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2555 = 6'h3b == select_39 ? io_inData_59 : _GEN_2554; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2556 = 6'h3c == select_39 ? io_inData_60 : _GEN_2555; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2557 = 6'h3d == select_39 ? io_inData_61 : _GEN_2556; // @[Switch.scala 33:19:@12824.4]
  assign _GEN_2558 = 6'h3e == select_39 ? io_inData_62 : _GEN_2557; // @[Switch.scala 33:19:@12824.4]
  assign _T_32994 = {valid_39_7,valid_39_6,valid_39_5,valid_39_4,valid_39_3,valid_39_2,valid_39_1,valid_39_0}; // @[Switch.scala 34:32:@12831.4]
  assign _T_33002 = {valid_39_15,valid_39_14,valid_39_13,valid_39_12,valid_39_11,valid_39_10,valid_39_9,valid_39_8,_T_32994}; // @[Switch.scala 34:32:@12839.4]
  assign _T_33009 = {valid_39_23,valid_39_22,valid_39_21,valid_39_20,valid_39_19,valid_39_18,valid_39_17,valid_39_16}; // @[Switch.scala 34:32:@12846.4]
  assign _T_33018 = {valid_39_31,valid_39_30,valid_39_29,valid_39_28,valid_39_27,valid_39_26,valid_39_25,valid_39_24,_T_33009,_T_33002}; // @[Switch.scala 34:32:@12855.4]
  assign _T_33025 = {valid_39_39,valid_39_38,valid_39_37,valid_39_36,valid_39_35,valid_39_34,valid_39_33,valid_39_32}; // @[Switch.scala 34:32:@12862.4]
  assign _T_33033 = {valid_39_47,valid_39_46,valid_39_45,valid_39_44,valid_39_43,valid_39_42,valid_39_41,valid_39_40,_T_33025}; // @[Switch.scala 34:32:@12870.4]
  assign _T_33040 = {valid_39_55,valid_39_54,valid_39_53,valid_39_52,valid_39_51,valid_39_50,valid_39_49,valid_39_48}; // @[Switch.scala 34:32:@12877.4]
  assign _T_33049 = {valid_39_63,valid_39_62,valid_39_61,valid_39_60,valid_39_59,valid_39_58,valid_39_57,valid_39_56,_T_33040,_T_33033}; // @[Switch.scala 34:32:@12886.4]
  assign _T_33050 = {_T_33049,_T_33018}; // @[Switch.scala 34:32:@12887.4]
  assign _T_33054 = io_inAddr_0 == 6'h28; // @[Switch.scala 30:53:@12890.4]
  assign valid_40_0 = io_inValid_0 & _T_33054; // @[Switch.scala 30:36:@12891.4]
  assign _T_33057 = io_inAddr_1 == 6'h28; // @[Switch.scala 30:53:@12893.4]
  assign valid_40_1 = io_inValid_1 & _T_33057; // @[Switch.scala 30:36:@12894.4]
  assign _T_33060 = io_inAddr_2 == 6'h28; // @[Switch.scala 30:53:@12896.4]
  assign valid_40_2 = io_inValid_2 & _T_33060; // @[Switch.scala 30:36:@12897.4]
  assign _T_33063 = io_inAddr_3 == 6'h28; // @[Switch.scala 30:53:@12899.4]
  assign valid_40_3 = io_inValid_3 & _T_33063; // @[Switch.scala 30:36:@12900.4]
  assign _T_33066 = io_inAddr_4 == 6'h28; // @[Switch.scala 30:53:@12902.4]
  assign valid_40_4 = io_inValid_4 & _T_33066; // @[Switch.scala 30:36:@12903.4]
  assign _T_33069 = io_inAddr_5 == 6'h28; // @[Switch.scala 30:53:@12905.4]
  assign valid_40_5 = io_inValid_5 & _T_33069; // @[Switch.scala 30:36:@12906.4]
  assign _T_33072 = io_inAddr_6 == 6'h28; // @[Switch.scala 30:53:@12908.4]
  assign valid_40_6 = io_inValid_6 & _T_33072; // @[Switch.scala 30:36:@12909.4]
  assign _T_33075 = io_inAddr_7 == 6'h28; // @[Switch.scala 30:53:@12911.4]
  assign valid_40_7 = io_inValid_7 & _T_33075; // @[Switch.scala 30:36:@12912.4]
  assign _T_33078 = io_inAddr_8 == 6'h28; // @[Switch.scala 30:53:@12914.4]
  assign valid_40_8 = io_inValid_8 & _T_33078; // @[Switch.scala 30:36:@12915.4]
  assign _T_33081 = io_inAddr_9 == 6'h28; // @[Switch.scala 30:53:@12917.4]
  assign valid_40_9 = io_inValid_9 & _T_33081; // @[Switch.scala 30:36:@12918.4]
  assign _T_33084 = io_inAddr_10 == 6'h28; // @[Switch.scala 30:53:@12920.4]
  assign valid_40_10 = io_inValid_10 & _T_33084; // @[Switch.scala 30:36:@12921.4]
  assign _T_33087 = io_inAddr_11 == 6'h28; // @[Switch.scala 30:53:@12923.4]
  assign valid_40_11 = io_inValid_11 & _T_33087; // @[Switch.scala 30:36:@12924.4]
  assign _T_33090 = io_inAddr_12 == 6'h28; // @[Switch.scala 30:53:@12926.4]
  assign valid_40_12 = io_inValid_12 & _T_33090; // @[Switch.scala 30:36:@12927.4]
  assign _T_33093 = io_inAddr_13 == 6'h28; // @[Switch.scala 30:53:@12929.4]
  assign valid_40_13 = io_inValid_13 & _T_33093; // @[Switch.scala 30:36:@12930.4]
  assign _T_33096 = io_inAddr_14 == 6'h28; // @[Switch.scala 30:53:@12932.4]
  assign valid_40_14 = io_inValid_14 & _T_33096; // @[Switch.scala 30:36:@12933.4]
  assign _T_33099 = io_inAddr_15 == 6'h28; // @[Switch.scala 30:53:@12935.4]
  assign valid_40_15 = io_inValid_15 & _T_33099; // @[Switch.scala 30:36:@12936.4]
  assign _T_33102 = io_inAddr_16 == 6'h28; // @[Switch.scala 30:53:@12938.4]
  assign valid_40_16 = io_inValid_16 & _T_33102; // @[Switch.scala 30:36:@12939.4]
  assign _T_33105 = io_inAddr_17 == 6'h28; // @[Switch.scala 30:53:@12941.4]
  assign valid_40_17 = io_inValid_17 & _T_33105; // @[Switch.scala 30:36:@12942.4]
  assign _T_33108 = io_inAddr_18 == 6'h28; // @[Switch.scala 30:53:@12944.4]
  assign valid_40_18 = io_inValid_18 & _T_33108; // @[Switch.scala 30:36:@12945.4]
  assign _T_33111 = io_inAddr_19 == 6'h28; // @[Switch.scala 30:53:@12947.4]
  assign valid_40_19 = io_inValid_19 & _T_33111; // @[Switch.scala 30:36:@12948.4]
  assign _T_33114 = io_inAddr_20 == 6'h28; // @[Switch.scala 30:53:@12950.4]
  assign valid_40_20 = io_inValid_20 & _T_33114; // @[Switch.scala 30:36:@12951.4]
  assign _T_33117 = io_inAddr_21 == 6'h28; // @[Switch.scala 30:53:@12953.4]
  assign valid_40_21 = io_inValid_21 & _T_33117; // @[Switch.scala 30:36:@12954.4]
  assign _T_33120 = io_inAddr_22 == 6'h28; // @[Switch.scala 30:53:@12956.4]
  assign valid_40_22 = io_inValid_22 & _T_33120; // @[Switch.scala 30:36:@12957.4]
  assign _T_33123 = io_inAddr_23 == 6'h28; // @[Switch.scala 30:53:@12959.4]
  assign valid_40_23 = io_inValid_23 & _T_33123; // @[Switch.scala 30:36:@12960.4]
  assign _T_33126 = io_inAddr_24 == 6'h28; // @[Switch.scala 30:53:@12962.4]
  assign valid_40_24 = io_inValid_24 & _T_33126; // @[Switch.scala 30:36:@12963.4]
  assign _T_33129 = io_inAddr_25 == 6'h28; // @[Switch.scala 30:53:@12965.4]
  assign valid_40_25 = io_inValid_25 & _T_33129; // @[Switch.scala 30:36:@12966.4]
  assign _T_33132 = io_inAddr_26 == 6'h28; // @[Switch.scala 30:53:@12968.4]
  assign valid_40_26 = io_inValid_26 & _T_33132; // @[Switch.scala 30:36:@12969.4]
  assign _T_33135 = io_inAddr_27 == 6'h28; // @[Switch.scala 30:53:@12971.4]
  assign valid_40_27 = io_inValid_27 & _T_33135; // @[Switch.scala 30:36:@12972.4]
  assign _T_33138 = io_inAddr_28 == 6'h28; // @[Switch.scala 30:53:@12974.4]
  assign valid_40_28 = io_inValid_28 & _T_33138; // @[Switch.scala 30:36:@12975.4]
  assign _T_33141 = io_inAddr_29 == 6'h28; // @[Switch.scala 30:53:@12977.4]
  assign valid_40_29 = io_inValid_29 & _T_33141; // @[Switch.scala 30:36:@12978.4]
  assign _T_33144 = io_inAddr_30 == 6'h28; // @[Switch.scala 30:53:@12980.4]
  assign valid_40_30 = io_inValid_30 & _T_33144; // @[Switch.scala 30:36:@12981.4]
  assign _T_33147 = io_inAddr_31 == 6'h28; // @[Switch.scala 30:53:@12983.4]
  assign valid_40_31 = io_inValid_31 & _T_33147; // @[Switch.scala 30:36:@12984.4]
  assign _T_33150 = io_inAddr_32 == 6'h28; // @[Switch.scala 30:53:@12986.4]
  assign valid_40_32 = io_inValid_32 & _T_33150; // @[Switch.scala 30:36:@12987.4]
  assign _T_33153 = io_inAddr_33 == 6'h28; // @[Switch.scala 30:53:@12989.4]
  assign valid_40_33 = io_inValid_33 & _T_33153; // @[Switch.scala 30:36:@12990.4]
  assign _T_33156 = io_inAddr_34 == 6'h28; // @[Switch.scala 30:53:@12992.4]
  assign valid_40_34 = io_inValid_34 & _T_33156; // @[Switch.scala 30:36:@12993.4]
  assign _T_33159 = io_inAddr_35 == 6'h28; // @[Switch.scala 30:53:@12995.4]
  assign valid_40_35 = io_inValid_35 & _T_33159; // @[Switch.scala 30:36:@12996.4]
  assign _T_33162 = io_inAddr_36 == 6'h28; // @[Switch.scala 30:53:@12998.4]
  assign valid_40_36 = io_inValid_36 & _T_33162; // @[Switch.scala 30:36:@12999.4]
  assign _T_33165 = io_inAddr_37 == 6'h28; // @[Switch.scala 30:53:@13001.4]
  assign valid_40_37 = io_inValid_37 & _T_33165; // @[Switch.scala 30:36:@13002.4]
  assign _T_33168 = io_inAddr_38 == 6'h28; // @[Switch.scala 30:53:@13004.4]
  assign valid_40_38 = io_inValid_38 & _T_33168; // @[Switch.scala 30:36:@13005.4]
  assign _T_33171 = io_inAddr_39 == 6'h28; // @[Switch.scala 30:53:@13007.4]
  assign valid_40_39 = io_inValid_39 & _T_33171; // @[Switch.scala 30:36:@13008.4]
  assign _T_33174 = io_inAddr_40 == 6'h28; // @[Switch.scala 30:53:@13010.4]
  assign valid_40_40 = io_inValid_40 & _T_33174; // @[Switch.scala 30:36:@13011.4]
  assign _T_33177 = io_inAddr_41 == 6'h28; // @[Switch.scala 30:53:@13013.4]
  assign valid_40_41 = io_inValid_41 & _T_33177; // @[Switch.scala 30:36:@13014.4]
  assign _T_33180 = io_inAddr_42 == 6'h28; // @[Switch.scala 30:53:@13016.4]
  assign valid_40_42 = io_inValid_42 & _T_33180; // @[Switch.scala 30:36:@13017.4]
  assign _T_33183 = io_inAddr_43 == 6'h28; // @[Switch.scala 30:53:@13019.4]
  assign valid_40_43 = io_inValid_43 & _T_33183; // @[Switch.scala 30:36:@13020.4]
  assign _T_33186 = io_inAddr_44 == 6'h28; // @[Switch.scala 30:53:@13022.4]
  assign valid_40_44 = io_inValid_44 & _T_33186; // @[Switch.scala 30:36:@13023.4]
  assign _T_33189 = io_inAddr_45 == 6'h28; // @[Switch.scala 30:53:@13025.4]
  assign valid_40_45 = io_inValid_45 & _T_33189; // @[Switch.scala 30:36:@13026.4]
  assign _T_33192 = io_inAddr_46 == 6'h28; // @[Switch.scala 30:53:@13028.4]
  assign valid_40_46 = io_inValid_46 & _T_33192; // @[Switch.scala 30:36:@13029.4]
  assign _T_33195 = io_inAddr_47 == 6'h28; // @[Switch.scala 30:53:@13031.4]
  assign valid_40_47 = io_inValid_47 & _T_33195; // @[Switch.scala 30:36:@13032.4]
  assign _T_33198 = io_inAddr_48 == 6'h28; // @[Switch.scala 30:53:@13034.4]
  assign valid_40_48 = io_inValid_48 & _T_33198; // @[Switch.scala 30:36:@13035.4]
  assign _T_33201 = io_inAddr_49 == 6'h28; // @[Switch.scala 30:53:@13037.4]
  assign valid_40_49 = io_inValid_49 & _T_33201; // @[Switch.scala 30:36:@13038.4]
  assign _T_33204 = io_inAddr_50 == 6'h28; // @[Switch.scala 30:53:@13040.4]
  assign valid_40_50 = io_inValid_50 & _T_33204; // @[Switch.scala 30:36:@13041.4]
  assign _T_33207 = io_inAddr_51 == 6'h28; // @[Switch.scala 30:53:@13043.4]
  assign valid_40_51 = io_inValid_51 & _T_33207; // @[Switch.scala 30:36:@13044.4]
  assign _T_33210 = io_inAddr_52 == 6'h28; // @[Switch.scala 30:53:@13046.4]
  assign valid_40_52 = io_inValid_52 & _T_33210; // @[Switch.scala 30:36:@13047.4]
  assign _T_33213 = io_inAddr_53 == 6'h28; // @[Switch.scala 30:53:@13049.4]
  assign valid_40_53 = io_inValid_53 & _T_33213; // @[Switch.scala 30:36:@13050.4]
  assign _T_33216 = io_inAddr_54 == 6'h28; // @[Switch.scala 30:53:@13052.4]
  assign valid_40_54 = io_inValid_54 & _T_33216; // @[Switch.scala 30:36:@13053.4]
  assign _T_33219 = io_inAddr_55 == 6'h28; // @[Switch.scala 30:53:@13055.4]
  assign valid_40_55 = io_inValid_55 & _T_33219; // @[Switch.scala 30:36:@13056.4]
  assign _T_33222 = io_inAddr_56 == 6'h28; // @[Switch.scala 30:53:@13058.4]
  assign valid_40_56 = io_inValid_56 & _T_33222; // @[Switch.scala 30:36:@13059.4]
  assign _T_33225 = io_inAddr_57 == 6'h28; // @[Switch.scala 30:53:@13061.4]
  assign valid_40_57 = io_inValid_57 & _T_33225; // @[Switch.scala 30:36:@13062.4]
  assign _T_33228 = io_inAddr_58 == 6'h28; // @[Switch.scala 30:53:@13064.4]
  assign valid_40_58 = io_inValid_58 & _T_33228; // @[Switch.scala 30:36:@13065.4]
  assign _T_33231 = io_inAddr_59 == 6'h28; // @[Switch.scala 30:53:@13067.4]
  assign valid_40_59 = io_inValid_59 & _T_33231; // @[Switch.scala 30:36:@13068.4]
  assign _T_33234 = io_inAddr_60 == 6'h28; // @[Switch.scala 30:53:@13070.4]
  assign valid_40_60 = io_inValid_60 & _T_33234; // @[Switch.scala 30:36:@13071.4]
  assign _T_33237 = io_inAddr_61 == 6'h28; // @[Switch.scala 30:53:@13073.4]
  assign valid_40_61 = io_inValid_61 & _T_33237; // @[Switch.scala 30:36:@13074.4]
  assign _T_33240 = io_inAddr_62 == 6'h28; // @[Switch.scala 30:53:@13076.4]
  assign valid_40_62 = io_inValid_62 & _T_33240; // @[Switch.scala 30:36:@13077.4]
  assign _T_33243 = io_inAddr_63 == 6'h28; // @[Switch.scala 30:53:@13079.4]
  assign valid_40_63 = io_inValid_63 & _T_33243; // @[Switch.scala 30:36:@13080.4]
  assign _T_33309 = valid_40_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@13082.4]
  assign _T_33310 = valid_40_61 ? 6'h3d : _T_33309; // @[Mux.scala 31:69:@13083.4]
  assign _T_33311 = valid_40_60 ? 6'h3c : _T_33310; // @[Mux.scala 31:69:@13084.4]
  assign _T_33312 = valid_40_59 ? 6'h3b : _T_33311; // @[Mux.scala 31:69:@13085.4]
  assign _T_33313 = valid_40_58 ? 6'h3a : _T_33312; // @[Mux.scala 31:69:@13086.4]
  assign _T_33314 = valid_40_57 ? 6'h39 : _T_33313; // @[Mux.scala 31:69:@13087.4]
  assign _T_33315 = valid_40_56 ? 6'h38 : _T_33314; // @[Mux.scala 31:69:@13088.4]
  assign _T_33316 = valid_40_55 ? 6'h37 : _T_33315; // @[Mux.scala 31:69:@13089.4]
  assign _T_33317 = valid_40_54 ? 6'h36 : _T_33316; // @[Mux.scala 31:69:@13090.4]
  assign _T_33318 = valid_40_53 ? 6'h35 : _T_33317; // @[Mux.scala 31:69:@13091.4]
  assign _T_33319 = valid_40_52 ? 6'h34 : _T_33318; // @[Mux.scala 31:69:@13092.4]
  assign _T_33320 = valid_40_51 ? 6'h33 : _T_33319; // @[Mux.scala 31:69:@13093.4]
  assign _T_33321 = valid_40_50 ? 6'h32 : _T_33320; // @[Mux.scala 31:69:@13094.4]
  assign _T_33322 = valid_40_49 ? 6'h31 : _T_33321; // @[Mux.scala 31:69:@13095.4]
  assign _T_33323 = valid_40_48 ? 6'h30 : _T_33322; // @[Mux.scala 31:69:@13096.4]
  assign _T_33324 = valid_40_47 ? 6'h2f : _T_33323; // @[Mux.scala 31:69:@13097.4]
  assign _T_33325 = valid_40_46 ? 6'h2e : _T_33324; // @[Mux.scala 31:69:@13098.4]
  assign _T_33326 = valid_40_45 ? 6'h2d : _T_33325; // @[Mux.scala 31:69:@13099.4]
  assign _T_33327 = valid_40_44 ? 6'h2c : _T_33326; // @[Mux.scala 31:69:@13100.4]
  assign _T_33328 = valid_40_43 ? 6'h2b : _T_33327; // @[Mux.scala 31:69:@13101.4]
  assign _T_33329 = valid_40_42 ? 6'h2a : _T_33328; // @[Mux.scala 31:69:@13102.4]
  assign _T_33330 = valid_40_41 ? 6'h29 : _T_33329; // @[Mux.scala 31:69:@13103.4]
  assign _T_33331 = valid_40_40 ? 6'h28 : _T_33330; // @[Mux.scala 31:69:@13104.4]
  assign _T_33332 = valid_40_39 ? 6'h27 : _T_33331; // @[Mux.scala 31:69:@13105.4]
  assign _T_33333 = valid_40_38 ? 6'h26 : _T_33332; // @[Mux.scala 31:69:@13106.4]
  assign _T_33334 = valid_40_37 ? 6'h25 : _T_33333; // @[Mux.scala 31:69:@13107.4]
  assign _T_33335 = valid_40_36 ? 6'h24 : _T_33334; // @[Mux.scala 31:69:@13108.4]
  assign _T_33336 = valid_40_35 ? 6'h23 : _T_33335; // @[Mux.scala 31:69:@13109.4]
  assign _T_33337 = valid_40_34 ? 6'h22 : _T_33336; // @[Mux.scala 31:69:@13110.4]
  assign _T_33338 = valid_40_33 ? 6'h21 : _T_33337; // @[Mux.scala 31:69:@13111.4]
  assign _T_33339 = valid_40_32 ? 6'h20 : _T_33338; // @[Mux.scala 31:69:@13112.4]
  assign _T_33340 = valid_40_31 ? 6'h1f : _T_33339; // @[Mux.scala 31:69:@13113.4]
  assign _T_33341 = valid_40_30 ? 6'h1e : _T_33340; // @[Mux.scala 31:69:@13114.4]
  assign _T_33342 = valid_40_29 ? 6'h1d : _T_33341; // @[Mux.scala 31:69:@13115.4]
  assign _T_33343 = valid_40_28 ? 6'h1c : _T_33342; // @[Mux.scala 31:69:@13116.4]
  assign _T_33344 = valid_40_27 ? 6'h1b : _T_33343; // @[Mux.scala 31:69:@13117.4]
  assign _T_33345 = valid_40_26 ? 6'h1a : _T_33344; // @[Mux.scala 31:69:@13118.4]
  assign _T_33346 = valid_40_25 ? 6'h19 : _T_33345; // @[Mux.scala 31:69:@13119.4]
  assign _T_33347 = valid_40_24 ? 6'h18 : _T_33346; // @[Mux.scala 31:69:@13120.4]
  assign _T_33348 = valid_40_23 ? 6'h17 : _T_33347; // @[Mux.scala 31:69:@13121.4]
  assign _T_33349 = valid_40_22 ? 6'h16 : _T_33348; // @[Mux.scala 31:69:@13122.4]
  assign _T_33350 = valid_40_21 ? 6'h15 : _T_33349; // @[Mux.scala 31:69:@13123.4]
  assign _T_33351 = valid_40_20 ? 6'h14 : _T_33350; // @[Mux.scala 31:69:@13124.4]
  assign _T_33352 = valid_40_19 ? 6'h13 : _T_33351; // @[Mux.scala 31:69:@13125.4]
  assign _T_33353 = valid_40_18 ? 6'h12 : _T_33352; // @[Mux.scala 31:69:@13126.4]
  assign _T_33354 = valid_40_17 ? 6'h11 : _T_33353; // @[Mux.scala 31:69:@13127.4]
  assign _T_33355 = valid_40_16 ? 6'h10 : _T_33354; // @[Mux.scala 31:69:@13128.4]
  assign _T_33356 = valid_40_15 ? 6'hf : _T_33355; // @[Mux.scala 31:69:@13129.4]
  assign _T_33357 = valid_40_14 ? 6'he : _T_33356; // @[Mux.scala 31:69:@13130.4]
  assign _T_33358 = valid_40_13 ? 6'hd : _T_33357; // @[Mux.scala 31:69:@13131.4]
  assign _T_33359 = valid_40_12 ? 6'hc : _T_33358; // @[Mux.scala 31:69:@13132.4]
  assign _T_33360 = valid_40_11 ? 6'hb : _T_33359; // @[Mux.scala 31:69:@13133.4]
  assign _T_33361 = valid_40_10 ? 6'ha : _T_33360; // @[Mux.scala 31:69:@13134.4]
  assign _T_33362 = valid_40_9 ? 6'h9 : _T_33361; // @[Mux.scala 31:69:@13135.4]
  assign _T_33363 = valid_40_8 ? 6'h8 : _T_33362; // @[Mux.scala 31:69:@13136.4]
  assign _T_33364 = valid_40_7 ? 6'h7 : _T_33363; // @[Mux.scala 31:69:@13137.4]
  assign _T_33365 = valid_40_6 ? 6'h6 : _T_33364; // @[Mux.scala 31:69:@13138.4]
  assign _T_33366 = valid_40_5 ? 6'h5 : _T_33365; // @[Mux.scala 31:69:@13139.4]
  assign _T_33367 = valid_40_4 ? 6'h4 : _T_33366; // @[Mux.scala 31:69:@13140.4]
  assign _T_33368 = valid_40_3 ? 6'h3 : _T_33367; // @[Mux.scala 31:69:@13141.4]
  assign _T_33369 = valid_40_2 ? 6'h2 : _T_33368; // @[Mux.scala 31:69:@13142.4]
  assign _T_33370 = valid_40_1 ? 6'h1 : _T_33369; // @[Mux.scala 31:69:@13143.4]
  assign select_40 = valid_40_0 ? 6'h0 : _T_33370; // @[Mux.scala 31:69:@13144.4]
  assign _GEN_2561 = 6'h1 == select_40 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2562 = 6'h2 == select_40 ? io_inData_2 : _GEN_2561; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2563 = 6'h3 == select_40 ? io_inData_3 : _GEN_2562; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2564 = 6'h4 == select_40 ? io_inData_4 : _GEN_2563; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2565 = 6'h5 == select_40 ? io_inData_5 : _GEN_2564; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2566 = 6'h6 == select_40 ? io_inData_6 : _GEN_2565; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2567 = 6'h7 == select_40 ? io_inData_7 : _GEN_2566; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2568 = 6'h8 == select_40 ? io_inData_8 : _GEN_2567; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2569 = 6'h9 == select_40 ? io_inData_9 : _GEN_2568; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2570 = 6'ha == select_40 ? io_inData_10 : _GEN_2569; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2571 = 6'hb == select_40 ? io_inData_11 : _GEN_2570; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2572 = 6'hc == select_40 ? io_inData_12 : _GEN_2571; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2573 = 6'hd == select_40 ? io_inData_13 : _GEN_2572; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2574 = 6'he == select_40 ? io_inData_14 : _GEN_2573; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2575 = 6'hf == select_40 ? io_inData_15 : _GEN_2574; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2576 = 6'h10 == select_40 ? io_inData_16 : _GEN_2575; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2577 = 6'h11 == select_40 ? io_inData_17 : _GEN_2576; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2578 = 6'h12 == select_40 ? io_inData_18 : _GEN_2577; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2579 = 6'h13 == select_40 ? io_inData_19 : _GEN_2578; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2580 = 6'h14 == select_40 ? io_inData_20 : _GEN_2579; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2581 = 6'h15 == select_40 ? io_inData_21 : _GEN_2580; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2582 = 6'h16 == select_40 ? io_inData_22 : _GEN_2581; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2583 = 6'h17 == select_40 ? io_inData_23 : _GEN_2582; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2584 = 6'h18 == select_40 ? io_inData_24 : _GEN_2583; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2585 = 6'h19 == select_40 ? io_inData_25 : _GEN_2584; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2586 = 6'h1a == select_40 ? io_inData_26 : _GEN_2585; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2587 = 6'h1b == select_40 ? io_inData_27 : _GEN_2586; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2588 = 6'h1c == select_40 ? io_inData_28 : _GEN_2587; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2589 = 6'h1d == select_40 ? io_inData_29 : _GEN_2588; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2590 = 6'h1e == select_40 ? io_inData_30 : _GEN_2589; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2591 = 6'h1f == select_40 ? io_inData_31 : _GEN_2590; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2592 = 6'h20 == select_40 ? io_inData_32 : _GEN_2591; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2593 = 6'h21 == select_40 ? io_inData_33 : _GEN_2592; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2594 = 6'h22 == select_40 ? io_inData_34 : _GEN_2593; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2595 = 6'h23 == select_40 ? io_inData_35 : _GEN_2594; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2596 = 6'h24 == select_40 ? io_inData_36 : _GEN_2595; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2597 = 6'h25 == select_40 ? io_inData_37 : _GEN_2596; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2598 = 6'h26 == select_40 ? io_inData_38 : _GEN_2597; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2599 = 6'h27 == select_40 ? io_inData_39 : _GEN_2598; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2600 = 6'h28 == select_40 ? io_inData_40 : _GEN_2599; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2601 = 6'h29 == select_40 ? io_inData_41 : _GEN_2600; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2602 = 6'h2a == select_40 ? io_inData_42 : _GEN_2601; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2603 = 6'h2b == select_40 ? io_inData_43 : _GEN_2602; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2604 = 6'h2c == select_40 ? io_inData_44 : _GEN_2603; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2605 = 6'h2d == select_40 ? io_inData_45 : _GEN_2604; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2606 = 6'h2e == select_40 ? io_inData_46 : _GEN_2605; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2607 = 6'h2f == select_40 ? io_inData_47 : _GEN_2606; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2608 = 6'h30 == select_40 ? io_inData_48 : _GEN_2607; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2609 = 6'h31 == select_40 ? io_inData_49 : _GEN_2608; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2610 = 6'h32 == select_40 ? io_inData_50 : _GEN_2609; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2611 = 6'h33 == select_40 ? io_inData_51 : _GEN_2610; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2612 = 6'h34 == select_40 ? io_inData_52 : _GEN_2611; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2613 = 6'h35 == select_40 ? io_inData_53 : _GEN_2612; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2614 = 6'h36 == select_40 ? io_inData_54 : _GEN_2613; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2615 = 6'h37 == select_40 ? io_inData_55 : _GEN_2614; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2616 = 6'h38 == select_40 ? io_inData_56 : _GEN_2615; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2617 = 6'h39 == select_40 ? io_inData_57 : _GEN_2616; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2618 = 6'h3a == select_40 ? io_inData_58 : _GEN_2617; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2619 = 6'h3b == select_40 ? io_inData_59 : _GEN_2618; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2620 = 6'h3c == select_40 ? io_inData_60 : _GEN_2619; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2621 = 6'h3d == select_40 ? io_inData_61 : _GEN_2620; // @[Switch.scala 33:19:@13146.4]
  assign _GEN_2622 = 6'h3e == select_40 ? io_inData_62 : _GEN_2621; // @[Switch.scala 33:19:@13146.4]
  assign _T_33379 = {valid_40_7,valid_40_6,valid_40_5,valid_40_4,valid_40_3,valid_40_2,valid_40_1,valid_40_0}; // @[Switch.scala 34:32:@13153.4]
  assign _T_33387 = {valid_40_15,valid_40_14,valid_40_13,valid_40_12,valid_40_11,valid_40_10,valid_40_9,valid_40_8,_T_33379}; // @[Switch.scala 34:32:@13161.4]
  assign _T_33394 = {valid_40_23,valid_40_22,valid_40_21,valid_40_20,valid_40_19,valid_40_18,valid_40_17,valid_40_16}; // @[Switch.scala 34:32:@13168.4]
  assign _T_33403 = {valid_40_31,valid_40_30,valid_40_29,valid_40_28,valid_40_27,valid_40_26,valid_40_25,valid_40_24,_T_33394,_T_33387}; // @[Switch.scala 34:32:@13177.4]
  assign _T_33410 = {valid_40_39,valid_40_38,valid_40_37,valid_40_36,valid_40_35,valid_40_34,valid_40_33,valid_40_32}; // @[Switch.scala 34:32:@13184.4]
  assign _T_33418 = {valid_40_47,valid_40_46,valid_40_45,valid_40_44,valid_40_43,valid_40_42,valid_40_41,valid_40_40,_T_33410}; // @[Switch.scala 34:32:@13192.4]
  assign _T_33425 = {valid_40_55,valid_40_54,valid_40_53,valid_40_52,valid_40_51,valid_40_50,valid_40_49,valid_40_48}; // @[Switch.scala 34:32:@13199.4]
  assign _T_33434 = {valid_40_63,valid_40_62,valid_40_61,valid_40_60,valid_40_59,valid_40_58,valid_40_57,valid_40_56,_T_33425,_T_33418}; // @[Switch.scala 34:32:@13208.4]
  assign _T_33435 = {_T_33434,_T_33403}; // @[Switch.scala 34:32:@13209.4]
  assign _T_33439 = io_inAddr_0 == 6'h29; // @[Switch.scala 30:53:@13212.4]
  assign valid_41_0 = io_inValid_0 & _T_33439; // @[Switch.scala 30:36:@13213.4]
  assign _T_33442 = io_inAddr_1 == 6'h29; // @[Switch.scala 30:53:@13215.4]
  assign valid_41_1 = io_inValid_1 & _T_33442; // @[Switch.scala 30:36:@13216.4]
  assign _T_33445 = io_inAddr_2 == 6'h29; // @[Switch.scala 30:53:@13218.4]
  assign valid_41_2 = io_inValid_2 & _T_33445; // @[Switch.scala 30:36:@13219.4]
  assign _T_33448 = io_inAddr_3 == 6'h29; // @[Switch.scala 30:53:@13221.4]
  assign valid_41_3 = io_inValid_3 & _T_33448; // @[Switch.scala 30:36:@13222.4]
  assign _T_33451 = io_inAddr_4 == 6'h29; // @[Switch.scala 30:53:@13224.4]
  assign valid_41_4 = io_inValid_4 & _T_33451; // @[Switch.scala 30:36:@13225.4]
  assign _T_33454 = io_inAddr_5 == 6'h29; // @[Switch.scala 30:53:@13227.4]
  assign valid_41_5 = io_inValid_5 & _T_33454; // @[Switch.scala 30:36:@13228.4]
  assign _T_33457 = io_inAddr_6 == 6'h29; // @[Switch.scala 30:53:@13230.4]
  assign valid_41_6 = io_inValid_6 & _T_33457; // @[Switch.scala 30:36:@13231.4]
  assign _T_33460 = io_inAddr_7 == 6'h29; // @[Switch.scala 30:53:@13233.4]
  assign valid_41_7 = io_inValid_7 & _T_33460; // @[Switch.scala 30:36:@13234.4]
  assign _T_33463 = io_inAddr_8 == 6'h29; // @[Switch.scala 30:53:@13236.4]
  assign valid_41_8 = io_inValid_8 & _T_33463; // @[Switch.scala 30:36:@13237.4]
  assign _T_33466 = io_inAddr_9 == 6'h29; // @[Switch.scala 30:53:@13239.4]
  assign valid_41_9 = io_inValid_9 & _T_33466; // @[Switch.scala 30:36:@13240.4]
  assign _T_33469 = io_inAddr_10 == 6'h29; // @[Switch.scala 30:53:@13242.4]
  assign valid_41_10 = io_inValid_10 & _T_33469; // @[Switch.scala 30:36:@13243.4]
  assign _T_33472 = io_inAddr_11 == 6'h29; // @[Switch.scala 30:53:@13245.4]
  assign valid_41_11 = io_inValid_11 & _T_33472; // @[Switch.scala 30:36:@13246.4]
  assign _T_33475 = io_inAddr_12 == 6'h29; // @[Switch.scala 30:53:@13248.4]
  assign valid_41_12 = io_inValid_12 & _T_33475; // @[Switch.scala 30:36:@13249.4]
  assign _T_33478 = io_inAddr_13 == 6'h29; // @[Switch.scala 30:53:@13251.4]
  assign valid_41_13 = io_inValid_13 & _T_33478; // @[Switch.scala 30:36:@13252.4]
  assign _T_33481 = io_inAddr_14 == 6'h29; // @[Switch.scala 30:53:@13254.4]
  assign valid_41_14 = io_inValid_14 & _T_33481; // @[Switch.scala 30:36:@13255.4]
  assign _T_33484 = io_inAddr_15 == 6'h29; // @[Switch.scala 30:53:@13257.4]
  assign valid_41_15 = io_inValid_15 & _T_33484; // @[Switch.scala 30:36:@13258.4]
  assign _T_33487 = io_inAddr_16 == 6'h29; // @[Switch.scala 30:53:@13260.4]
  assign valid_41_16 = io_inValid_16 & _T_33487; // @[Switch.scala 30:36:@13261.4]
  assign _T_33490 = io_inAddr_17 == 6'h29; // @[Switch.scala 30:53:@13263.4]
  assign valid_41_17 = io_inValid_17 & _T_33490; // @[Switch.scala 30:36:@13264.4]
  assign _T_33493 = io_inAddr_18 == 6'h29; // @[Switch.scala 30:53:@13266.4]
  assign valid_41_18 = io_inValid_18 & _T_33493; // @[Switch.scala 30:36:@13267.4]
  assign _T_33496 = io_inAddr_19 == 6'h29; // @[Switch.scala 30:53:@13269.4]
  assign valid_41_19 = io_inValid_19 & _T_33496; // @[Switch.scala 30:36:@13270.4]
  assign _T_33499 = io_inAddr_20 == 6'h29; // @[Switch.scala 30:53:@13272.4]
  assign valid_41_20 = io_inValid_20 & _T_33499; // @[Switch.scala 30:36:@13273.4]
  assign _T_33502 = io_inAddr_21 == 6'h29; // @[Switch.scala 30:53:@13275.4]
  assign valid_41_21 = io_inValid_21 & _T_33502; // @[Switch.scala 30:36:@13276.4]
  assign _T_33505 = io_inAddr_22 == 6'h29; // @[Switch.scala 30:53:@13278.4]
  assign valid_41_22 = io_inValid_22 & _T_33505; // @[Switch.scala 30:36:@13279.4]
  assign _T_33508 = io_inAddr_23 == 6'h29; // @[Switch.scala 30:53:@13281.4]
  assign valid_41_23 = io_inValid_23 & _T_33508; // @[Switch.scala 30:36:@13282.4]
  assign _T_33511 = io_inAddr_24 == 6'h29; // @[Switch.scala 30:53:@13284.4]
  assign valid_41_24 = io_inValid_24 & _T_33511; // @[Switch.scala 30:36:@13285.4]
  assign _T_33514 = io_inAddr_25 == 6'h29; // @[Switch.scala 30:53:@13287.4]
  assign valid_41_25 = io_inValid_25 & _T_33514; // @[Switch.scala 30:36:@13288.4]
  assign _T_33517 = io_inAddr_26 == 6'h29; // @[Switch.scala 30:53:@13290.4]
  assign valid_41_26 = io_inValid_26 & _T_33517; // @[Switch.scala 30:36:@13291.4]
  assign _T_33520 = io_inAddr_27 == 6'h29; // @[Switch.scala 30:53:@13293.4]
  assign valid_41_27 = io_inValid_27 & _T_33520; // @[Switch.scala 30:36:@13294.4]
  assign _T_33523 = io_inAddr_28 == 6'h29; // @[Switch.scala 30:53:@13296.4]
  assign valid_41_28 = io_inValid_28 & _T_33523; // @[Switch.scala 30:36:@13297.4]
  assign _T_33526 = io_inAddr_29 == 6'h29; // @[Switch.scala 30:53:@13299.4]
  assign valid_41_29 = io_inValid_29 & _T_33526; // @[Switch.scala 30:36:@13300.4]
  assign _T_33529 = io_inAddr_30 == 6'h29; // @[Switch.scala 30:53:@13302.4]
  assign valid_41_30 = io_inValid_30 & _T_33529; // @[Switch.scala 30:36:@13303.4]
  assign _T_33532 = io_inAddr_31 == 6'h29; // @[Switch.scala 30:53:@13305.4]
  assign valid_41_31 = io_inValid_31 & _T_33532; // @[Switch.scala 30:36:@13306.4]
  assign _T_33535 = io_inAddr_32 == 6'h29; // @[Switch.scala 30:53:@13308.4]
  assign valid_41_32 = io_inValid_32 & _T_33535; // @[Switch.scala 30:36:@13309.4]
  assign _T_33538 = io_inAddr_33 == 6'h29; // @[Switch.scala 30:53:@13311.4]
  assign valid_41_33 = io_inValid_33 & _T_33538; // @[Switch.scala 30:36:@13312.4]
  assign _T_33541 = io_inAddr_34 == 6'h29; // @[Switch.scala 30:53:@13314.4]
  assign valid_41_34 = io_inValid_34 & _T_33541; // @[Switch.scala 30:36:@13315.4]
  assign _T_33544 = io_inAddr_35 == 6'h29; // @[Switch.scala 30:53:@13317.4]
  assign valid_41_35 = io_inValid_35 & _T_33544; // @[Switch.scala 30:36:@13318.4]
  assign _T_33547 = io_inAddr_36 == 6'h29; // @[Switch.scala 30:53:@13320.4]
  assign valid_41_36 = io_inValid_36 & _T_33547; // @[Switch.scala 30:36:@13321.4]
  assign _T_33550 = io_inAddr_37 == 6'h29; // @[Switch.scala 30:53:@13323.4]
  assign valid_41_37 = io_inValid_37 & _T_33550; // @[Switch.scala 30:36:@13324.4]
  assign _T_33553 = io_inAddr_38 == 6'h29; // @[Switch.scala 30:53:@13326.4]
  assign valid_41_38 = io_inValid_38 & _T_33553; // @[Switch.scala 30:36:@13327.4]
  assign _T_33556 = io_inAddr_39 == 6'h29; // @[Switch.scala 30:53:@13329.4]
  assign valid_41_39 = io_inValid_39 & _T_33556; // @[Switch.scala 30:36:@13330.4]
  assign _T_33559 = io_inAddr_40 == 6'h29; // @[Switch.scala 30:53:@13332.4]
  assign valid_41_40 = io_inValid_40 & _T_33559; // @[Switch.scala 30:36:@13333.4]
  assign _T_33562 = io_inAddr_41 == 6'h29; // @[Switch.scala 30:53:@13335.4]
  assign valid_41_41 = io_inValid_41 & _T_33562; // @[Switch.scala 30:36:@13336.4]
  assign _T_33565 = io_inAddr_42 == 6'h29; // @[Switch.scala 30:53:@13338.4]
  assign valid_41_42 = io_inValid_42 & _T_33565; // @[Switch.scala 30:36:@13339.4]
  assign _T_33568 = io_inAddr_43 == 6'h29; // @[Switch.scala 30:53:@13341.4]
  assign valid_41_43 = io_inValid_43 & _T_33568; // @[Switch.scala 30:36:@13342.4]
  assign _T_33571 = io_inAddr_44 == 6'h29; // @[Switch.scala 30:53:@13344.4]
  assign valid_41_44 = io_inValid_44 & _T_33571; // @[Switch.scala 30:36:@13345.4]
  assign _T_33574 = io_inAddr_45 == 6'h29; // @[Switch.scala 30:53:@13347.4]
  assign valid_41_45 = io_inValid_45 & _T_33574; // @[Switch.scala 30:36:@13348.4]
  assign _T_33577 = io_inAddr_46 == 6'h29; // @[Switch.scala 30:53:@13350.4]
  assign valid_41_46 = io_inValid_46 & _T_33577; // @[Switch.scala 30:36:@13351.4]
  assign _T_33580 = io_inAddr_47 == 6'h29; // @[Switch.scala 30:53:@13353.4]
  assign valid_41_47 = io_inValid_47 & _T_33580; // @[Switch.scala 30:36:@13354.4]
  assign _T_33583 = io_inAddr_48 == 6'h29; // @[Switch.scala 30:53:@13356.4]
  assign valid_41_48 = io_inValid_48 & _T_33583; // @[Switch.scala 30:36:@13357.4]
  assign _T_33586 = io_inAddr_49 == 6'h29; // @[Switch.scala 30:53:@13359.4]
  assign valid_41_49 = io_inValid_49 & _T_33586; // @[Switch.scala 30:36:@13360.4]
  assign _T_33589 = io_inAddr_50 == 6'h29; // @[Switch.scala 30:53:@13362.4]
  assign valid_41_50 = io_inValid_50 & _T_33589; // @[Switch.scala 30:36:@13363.4]
  assign _T_33592 = io_inAddr_51 == 6'h29; // @[Switch.scala 30:53:@13365.4]
  assign valid_41_51 = io_inValid_51 & _T_33592; // @[Switch.scala 30:36:@13366.4]
  assign _T_33595 = io_inAddr_52 == 6'h29; // @[Switch.scala 30:53:@13368.4]
  assign valid_41_52 = io_inValid_52 & _T_33595; // @[Switch.scala 30:36:@13369.4]
  assign _T_33598 = io_inAddr_53 == 6'h29; // @[Switch.scala 30:53:@13371.4]
  assign valid_41_53 = io_inValid_53 & _T_33598; // @[Switch.scala 30:36:@13372.4]
  assign _T_33601 = io_inAddr_54 == 6'h29; // @[Switch.scala 30:53:@13374.4]
  assign valid_41_54 = io_inValid_54 & _T_33601; // @[Switch.scala 30:36:@13375.4]
  assign _T_33604 = io_inAddr_55 == 6'h29; // @[Switch.scala 30:53:@13377.4]
  assign valid_41_55 = io_inValid_55 & _T_33604; // @[Switch.scala 30:36:@13378.4]
  assign _T_33607 = io_inAddr_56 == 6'h29; // @[Switch.scala 30:53:@13380.4]
  assign valid_41_56 = io_inValid_56 & _T_33607; // @[Switch.scala 30:36:@13381.4]
  assign _T_33610 = io_inAddr_57 == 6'h29; // @[Switch.scala 30:53:@13383.4]
  assign valid_41_57 = io_inValid_57 & _T_33610; // @[Switch.scala 30:36:@13384.4]
  assign _T_33613 = io_inAddr_58 == 6'h29; // @[Switch.scala 30:53:@13386.4]
  assign valid_41_58 = io_inValid_58 & _T_33613; // @[Switch.scala 30:36:@13387.4]
  assign _T_33616 = io_inAddr_59 == 6'h29; // @[Switch.scala 30:53:@13389.4]
  assign valid_41_59 = io_inValid_59 & _T_33616; // @[Switch.scala 30:36:@13390.4]
  assign _T_33619 = io_inAddr_60 == 6'h29; // @[Switch.scala 30:53:@13392.4]
  assign valid_41_60 = io_inValid_60 & _T_33619; // @[Switch.scala 30:36:@13393.4]
  assign _T_33622 = io_inAddr_61 == 6'h29; // @[Switch.scala 30:53:@13395.4]
  assign valid_41_61 = io_inValid_61 & _T_33622; // @[Switch.scala 30:36:@13396.4]
  assign _T_33625 = io_inAddr_62 == 6'h29; // @[Switch.scala 30:53:@13398.4]
  assign valid_41_62 = io_inValid_62 & _T_33625; // @[Switch.scala 30:36:@13399.4]
  assign _T_33628 = io_inAddr_63 == 6'h29; // @[Switch.scala 30:53:@13401.4]
  assign valid_41_63 = io_inValid_63 & _T_33628; // @[Switch.scala 30:36:@13402.4]
  assign _T_33694 = valid_41_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@13404.4]
  assign _T_33695 = valid_41_61 ? 6'h3d : _T_33694; // @[Mux.scala 31:69:@13405.4]
  assign _T_33696 = valid_41_60 ? 6'h3c : _T_33695; // @[Mux.scala 31:69:@13406.4]
  assign _T_33697 = valid_41_59 ? 6'h3b : _T_33696; // @[Mux.scala 31:69:@13407.4]
  assign _T_33698 = valid_41_58 ? 6'h3a : _T_33697; // @[Mux.scala 31:69:@13408.4]
  assign _T_33699 = valid_41_57 ? 6'h39 : _T_33698; // @[Mux.scala 31:69:@13409.4]
  assign _T_33700 = valid_41_56 ? 6'h38 : _T_33699; // @[Mux.scala 31:69:@13410.4]
  assign _T_33701 = valid_41_55 ? 6'h37 : _T_33700; // @[Mux.scala 31:69:@13411.4]
  assign _T_33702 = valid_41_54 ? 6'h36 : _T_33701; // @[Mux.scala 31:69:@13412.4]
  assign _T_33703 = valid_41_53 ? 6'h35 : _T_33702; // @[Mux.scala 31:69:@13413.4]
  assign _T_33704 = valid_41_52 ? 6'h34 : _T_33703; // @[Mux.scala 31:69:@13414.4]
  assign _T_33705 = valid_41_51 ? 6'h33 : _T_33704; // @[Mux.scala 31:69:@13415.4]
  assign _T_33706 = valid_41_50 ? 6'h32 : _T_33705; // @[Mux.scala 31:69:@13416.4]
  assign _T_33707 = valid_41_49 ? 6'h31 : _T_33706; // @[Mux.scala 31:69:@13417.4]
  assign _T_33708 = valid_41_48 ? 6'h30 : _T_33707; // @[Mux.scala 31:69:@13418.4]
  assign _T_33709 = valid_41_47 ? 6'h2f : _T_33708; // @[Mux.scala 31:69:@13419.4]
  assign _T_33710 = valid_41_46 ? 6'h2e : _T_33709; // @[Mux.scala 31:69:@13420.4]
  assign _T_33711 = valid_41_45 ? 6'h2d : _T_33710; // @[Mux.scala 31:69:@13421.4]
  assign _T_33712 = valid_41_44 ? 6'h2c : _T_33711; // @[Mux.scala 31:69:@13422.4]
  assign _T_33713 = valid_41_43 ? 6'h2b : _T_33712; // @[Mux.scala 31:69:@13423.4]
  assign _T_33714 = valid_41_42 ? 6'h2a : _T_33713; // @[Mux.scala 31:69:@13424.4]
  assign _T_33715 = valid_41_41 ? 6'h29 : _T_33714; // @[Mux.scala 31:69:@13425.4]
  assign _T_33716 = valid_41_40 ? 6'h28 : _T_33715; // @[Mux.scala 31:69:@13426.4]
  assign _T_33717 = valid_41_39 ? 6'h27 : _T_33716; // @[Mux.scala 31:69:@13427.4]
  assign _T_33718 = valid_41_38 ? 6'h26 : _T_33717; // @[Mux.scala 31:69:@13428.4]
  assign _T_33719 = valid_41_37 ? 6'h25 : _T_33718; // @[Mux.scala 31:69:@13429.4]
  assign _T_33720 = valid_41_36 ? 6'h24 : _T_33719; // @[Mux.scala 31:69:@13430.4]
  assign _T_33721 = valid_41_35 ? 6'h23 : _T_33720; // @[Mux.scala 31:69:@13431.4]
  assign _T_33722 = valid_41_34 ? 6'h22 : _T_33721; // @[Mux.scala 31:69:@13432.4]
  assign _T_33723 = valid_41_33 ? 6'h21 : _T_33722; // @[Mux.scala 31:69:@13433.4]
  assign _T_33724 = valid_41_32 ? 6'h20 : _T_33723; // @[Mux.scala 31:69:@13434.4]
  assign _T_33725 = valid_41_31 ? 6'h1f : _T_33724; // @[Mux.scala 31:69:@13435.4]
  assign _T_33726 = valid_41_30 ? 6'h1e : _T_33725; // @[Mux.scala 31:69:@13436.4]
  assign _T_33727 = valid_41_29 ? 6'h1d : _T_33726; // @[Mux.scala 31:69:@13437.4]
  assign _T_33728 = valid_41_28 ? 6'h1c : _T_33727; // @[Mux.scala 31:69:@13438.4]
  assign _T_33729 = valid_41_27 ? 6'h1b : _T_33728; // @[Mux.scala 31:69:@13439.4]
  assign _T_33730 = valid_41_26 ? 6'h1a : _T_33729; // @[Mux.scala 31:69:@13440.4]
  assign _T_33731 = valid_41_25 ? 6'h19 : _T_33730; // @[Mux.scala 31:69:@13441.4]
  assign _T_33732 = valid_41_24 ? 6'h18 : _T_33731; // @[Mux.scala 31:69:@13442.4]
  assign _T_33733 = valid_41_23 ? 6'h17 : _T_33732; // @[Mux.scala 31:69:@13443.4]
  assign _T_33734 = valid_41_22 ? 6'h16 : _T_33733; // @[Mux.scala 31:69:@13444.4]
  assign _T_33735 = valid_41_21 ? 6'h15 : _T_33734; // @[Mux.scala 31:69:@13445.4]
  assign _T_33736 = valid_41_20 ? 6'h14 : _T_33735; // @[Mux.scala 31:69:@13446.4]
  assign _T_33737 = valid_41_19 ? 6'h13 : _T_33736; // @[Mux.scala 31:69:@13447.4]
  assign _T_33738 = valid_41_18 ? 6'h12 : _T_33737; // @[Mux.scala 31:69:@13448.4]
  assign _T_33739 = valid_41_17 ? 6'h11 : _T_33738; // @[Mux.scala 31:69:@13449.4]
  assign _T_33740 = valid_41_16 ? 6'h10 : _T_33739; // @[Mux.scala 31:69:@13450.4]
  assign _T_33741 = valid_41_15 ? 6'hf : _T_33740; // @[Mux.scala 31:69:@13451.4]
  assign _T_33742 = valid_41_14 ? 6'he : _T_33741; // @[Mux.scala 31:69:@13452.4]
  assign _T_33743 = valid_41_13 ? 6'hd : _T_33742; // @[Mux.scala 31:69:@13453.4]
  assign _T_33744 = valid_41_12 ? 6'hc : _T_33743; // @[Mux.scala 31:69:@13454.4]
  assign _T_33745 = valid_41_11 ? 6'hb : _T_33744; // @[Mux.scala 31:69:@13455.4]
  assign _T_33746 = valid_41_10 ? 6'ha : _T_33745; // @[Mux.scala 31:69:@13456.4]
  assign _T_33747 = valid_41_9 ? 6'h9 : _T_33746; // @[Mux.scala 31:69:@13457.4]
  assign _T_33748 = valid_41_8 ? 6'h8 : _T_33747; // @[Mux.scala 31:69:@13458.4]
  assign _T_33749 = valid_41_7 ? 6'h7 : _T_33748; // @[Mux.scala 31:69:@13459.4]
  assign _T_33750 = valid_41_6 ? 6'h6 : _T_33749; // @[Mux.scala 31:69:@13460.4]
  assign _T_33751 = valid_41_5 ? 6'h5 : _T_33750; // @[Mux.scala 31:69:@13461.4]
  assign _T_33752 = valid_41_4 ? 6'h4 : _T_33751; // @[Mux.scala 31:69:@13462.4]
  assign _T_33753 = valid_41_3 ? 6'h3 : _T_33752; // @[Mux.scala 31:69:@13463.4]
  assign _T_33754 = valid_41_2 ? 6'h2 : _T_33753; // @[Mux.scala 31:69:@13464.4]
  assign _T_33755 = valid_41_1 ? 6'h1 : _T_33754; // @[Mux.scala 31:69:@13465.4]
  assign select_41 = valid_41_0 ? 6'h0 : _T_33755; // @[Mux.scala 31:69:@13466.4]
  assign _GEN_2625 = 6'h1 == select_41 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2626 = 6'h2 == select_41 ? io_inData_2 : _GEN_2625; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2627 = 6'h3 == select_41 ? io_inData_3 : _GEN_2626; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2628 = 6'h4 == select_41 ? io_inData_4 : _GEN_2627; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2629 = 6'h5 == select_41 ? io_inData_5 : _GEN_2628; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2630 = 6'h6 == select_41 ? io_inData_6 : _GEN_2629; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2631 = 6'h7 == select_41 ? io_inData_7 : _GEN_2630; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2632 = 6'h8 == select_41 ? io_inData_8 : _GEN_2631; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2633 = 6'h9 == select_41 ? io_inData_9 : _GEN_2632; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2634 = 6'ha == select_41 ? io_inData_10 : _GEN_2633; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2635 = 6'hb == select_41 ? io_inData_11 : _GEN_2634; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2636 = 6'hc == select_41 ? io_inData_12 : _GEN_2635; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2637 = 6'hd == select_41 ? io_inData_13 : _GEN_2636; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2638 = 6'he == select_41 ? io_inData_14 : _GEN_2637; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2639 = 6'hf == select_41 ? io_inData_15 : _GEN_2638; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2640 = 6'h10 == select_41 ? io_inData_16 : _GEN_2639; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2641 = 6'h11 == select_41 ? io_inData_17 : _GEN_2640; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2642 = 6'h12 == select_41 ? io_inData_18 : _GEN_2641; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2643 = 6'h13 == select_41 ? io_inData_19 : _GEN_2642; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2644 = 6'h14 == select_41 ? io_inData_20 : _GEN_2643; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2645 = 6'h15 == select_41 ? io_inData_21 : _GEN_2644; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2646 = 6'h16 == select_41 ? io_inData_22 : _GEN_2645; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2647 = 6'h17 == select_41 ? io_inData_23 : _GEN_2646; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2648 = 6'h18 == select_41 ? io_inData_24 : _GEN_2647; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2649 = 6'h19 == select_41 ? io_inData_25 : _GEN_2648; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2650 = 6'h1a == select_41 ? io_inData_26 : _GEN_2649; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2651 = 6'h1b == select_41 ? io_inData_27 : _GEN_2650; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2652 = 6'h1c == select_41 ? io_inData_28 : _GEN_2651; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2653 = 6'h1d == select_41 ? io_inData_29 : _GEN_2652; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2654 = 6'h1e == select_41 ? io_inData_30 : _GEN_2653; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2655 = 6'h1f == select_41 ? io_inData_31 : _GEN_2654; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2656 = 6'h20 == select_41 ? io_inData_32 : _GEN_2655; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2657 = 6'h21 == select_41 ? io_inData_33 : _GEN_2656; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2658 = 6'h22 == select_41 ? io_inData_34 : _GEN_2657; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2659 = 6'h23 == select_41 ? io_inData_35 : _GEN_2658; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2660 = 6'h24 == select_41 ? io_inData_36 : _GEN_2659; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2661 = 6'h25 == select_41 ? io_inData_37 : _GEN_2660; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2662 = 6'h26 == select_41 ? io_inData_38 : _GEN_2661; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2663 = 6'h27 == select_41 ? io_inData_39 : _GEN_2662; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2664 = 6'h28 == select_41 ? io_inData_40 : _GEN_2663; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2665 = 6'h29 == select_41 ? io_inData_41 : _GEN_2664; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2666 = 6'h2a == select_41 ? io_inData_42 : _GEN_2665; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2667 = 6'h2b == select_41 ? io_inData_43 : _GEN_2666; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2668 = 6'h2c == select_41 ? io_inData_44 : _GEN_2667; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2669 = 6'h2d == select_41 ? io_inData_45 : _GEN_2668; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2670 = 6'h2e == select_41 ? io_inData_46 : _GEN_2669; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2671 = 6'h2f == select_41 ? io_inData_47 : _GEN_2670; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2672 = 6'h30 == select_41 ? io_inData_48 : _GEN_2671; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2673 = 6'h31 == select_41 ? io_inData_49 : _GEN_2672; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2674 = 6'h32 == select_41 ? io_inData_50 : _GEN_2673; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2675 = 6'h33 == select_41 ? io_inData_51 : _GEN_2674; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2676 = 6'h34 == select_41 ? io_inData_52 : _GEN_2675; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2677 = 6'h35 == select_41 ? io_inData_53 : _GEN_2676; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2678 = 6'h36 == select_41 ? io_inData_54 : _GEN_2677; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2679 = 6'h37 == select_41 ? io_inData_55 : _GEN_2678; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2680 = 6'h38 == select_41 ? io_inData_56 : _GEN_2679; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2681 = 6'h39 == select_41 ? io_inData_57 : _GEN_2680; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2682 = 6'h3a == select_41 ? io_inData_58 : _GEN_2681; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2683 = 6'h3b == select_41 ? io_inData_59 : _GEN_2682; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2684 = 6'h3c == select_41 ? io_inData_60 : _GEN_2683; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2685 = 6'h3d == select_41 ? io_inData_61 : _GEN_2684; // @[Switch.scala 33:19:@13468.4]
  assign _GEN_2686 = 6'h3e == select_41 ? io_inData_62 : _GEN_2685; // @[Switch.scala 33:19:@13468.4]
  assign _T_33764 = {valid_41_7,valid_41_6,valid_41_5,valid_41_4,valid_41_3,valid_41_2,valid_41_1,valid_41_0}; // @[Switch.scala 34:32:@13475.4]
  assign _T_33772 = {valid_41_15,valid_41_14,valid_41_13,valid_41_12,valid_41_11,valid_41_10,valid_41_9,valid_41_8,_T_33764}; // @[Switch.scala 34:32:@13483.4]
  assign _T_33779 = {valid_41_23,valid_41_22,valid_41_21,valid_41_20,valid_41_19,valid_41_18,valid_41_17,valid_41_16}; // @[Switch.scala 34:32:@13490.4]
  assign _T_33788 = {valid_41_31,valid_41_30,valid_41_29,valid_41_28,valid_41_27,valid_41_26,valid_41_25,valid_41_24,_T_33779,_T_33772}; // @[Switch.scala 34:32:@13499.4]
  assign _T_33795 = {valid_41_39,valid_41_38,valid_41_37,valid_41_36,valid_41_35,valid_41_34,valid_41_33,valid_41_32}; // @[Switch.scala 34:32:@13506.4]
  assign _T_33803 = {valid_41_47,valid_41_46,valid_41_45,valid_41_44,valid_41_43,valid_41_42,valid_41_41,valid_41_40,_T_33795}; // @[Switch.scala 34:32:@13514.4]
  assign _T_33810 = {valid_41_55,valid_41_54,valid_41_53,valid_41_52,valid_41_51,valid_41_50,valid_41_49,valid_41_48}; // @[Switch.scala 34:32:@13521.4]
  assign _T_33819 = {valid_41_63,valid_41_62,valid_41_61,valid_41_60,valid_41_59,valid_41_58,valid_41_57,valid_41_56,_T_33810,_T_33803}; // @[Switch.scala 34:32:@13530.4]
  assign _T_33820 = {_T_33819,_T_33788}; // @[Switch.scala 34:32:@13531.4]
  assign _T_33824 = io_inAddr_0 == 6'h2a; // @[Switch.scala 30:53:@13534.4]
  assign valid_42_0 = io_inValid_0 & _T_33824; // @[Switch.scala 30:36:@13535.4]
  assign _T_33827 = io_inAddr_1 == 6'h2a; // @[Switch.scala 30:53:@13537.4]
  assign valid_42_1 = io_inValid_1 & _T_33827; // @[Switch.scala 30:36:@13538.4]
  assign _T_33830 = io_inAddr_2 == 6'h2a; // @[Switch.scala 30:53:@13540.4]
  assign valid_42_2 = io_inValid_2 & _T_33830; // @[Switch.scala 30:36:@13541.4]
  assign _T_33833 = io_inAddr_3 == 6'h2a; // @[Switch.scala 30:53:@13543.4]
  assign valid_42_3 = io_inValid_3 & _T_33833; // @[Switch.scala 30:36:@13544.4]
  assign _T_33836 = io_inAddr_4 == 6'h2a; // @[Switch.scala 30:53:@13546.4]
  assign valid_42_4 = io_inValid_4 & _T_33836; // @[Switch.scala 30:36:@13547.4]
  assign _T_33839 = io_inAddr_5 == 6'h2a; // @[Switch.scala 30:53:@13549.4]
  assign valid_42_5 = io_inValid_5 & _T_33839; // @[Switch.scala 30:36:@13550.4]
  assign _T_33842 = io_inAddr_6 == 6'h2a; // @[Switch.scala 30:53:@13552.4]
  assign valid_42_6 = io_inValid_6 & _T_33842; // @[Switch.scala 30:36:@13553.4]
  assign _T_33845 = io_inAddr_7 == 6'h2a; // @[Switch.scala 30:53:@13555.4]
  assign valid_42_7 = io_inValid_7 & _T_33845; // @[Switch.scala 30:36:@13556.4]
  assign _T_33848 = io_inAddr_8 == 6'h2a; // @[Switch.scala 30:53:@13558.4]
  assign valid_42_8 = io_inValid_8 & _T_33848; // @[Switch.scala 30:36:@13559.4]
  assign _T_33851 = io_inAddr_9 == 6'h2a; // @[Switch.scala 30:53:@13561.4]
  assign valid_42_9 = io_inValid_9 & _T_33851; // @[Switch.scala 30:36:@13562.4]
  assign _T_33854 = io_inAddr_10 == 6'h2a; // @[Switch.scala 30:53:@13564.4]
  assign valid_42_10 = io_inValid_10 & _T_33854; // @[Switch.scala 30:36:@13565.4]
  assign _T_33857 = io_inAddr_11 == 6'h2a; // @[Switch.scala 30:53:@13567.4]
  assign valid_42_11 = io_inValid_11 & _T_33857; // @[Switch.scala 30:36:@13568.4]
  assign _T_33860 = io_inAddr_12 == 6'h2a; // @[Switch.scala 30:53:@13570.4]
  assign valid_42_12 = io_inValid_12 & _T_33860; // @[Switch.scala 30:36:@13571.4]
  assign _T_33863 = io_inAddr_13 == 6'h2a; // @[Switch.scala 30:53:@13573.4]
  assign valid_42_13 = io_inValid_13 & _T_33863; // @[Switch.scala 30:36:@13574.4]
  assign _T_33866 = io_inAddr_14 == 6'h2a; // @[Switch.scala 30:53:@13576.4]
  assign valid_42_14 = io_inValid_14 & _T_33866; // @[Switch.scala 30:36:@13577.4]
  assign _T_33869 = io_inAddr_15 == 6'h2a; // @[Switch.scala 30:53:@13579.4]
  assign valid_42_15 = io_inValid_15 & _T_33869; // @[Switch.scala 30:36:@13580.4]
  assign _T_33872 = io_inAddr_16 == 6'h2a; // @[Switch.scala 30:53:@13582.4]
  assign valid_42_16 = io_inValid_16 & _T_33872; // @[Switch.scala 30:36:@13583.4]
  assign _T_33875 = io_inAddr_17 == 6'h2a; // @[Switch.scala 30:53:@13585.4]
  assign valid_42_17 = io_inValid_17 & _T_33875; // @[Switch.scala 30:36:@13586.4]
  assign _T_33878 = io_inAddr_18 == 6'h2a; // @[Switch.scala 30:53:@13588.4]
  assign valid_42_18 = io_inValid_18 & _T_33878; // @[Switch.scala 30:36:@13589.4]
  assign _T_33881 = io_inAddr_19 == 6'h2a; // @[Switch.scala 30:53:@13591.4]
  assign valid_42_19 = io_inValid_19 & _T_33881; // @[Switch.scala 30:36:@13592.4]
  assign _T_33884 = io_inAddr_20 == 6'h2a; // @[Switch.scala 30:53:@13594.4]
  assign valid_42_20 = io_inValid_20 & _T_33884; // @[Switch.scala 30:36:@13595.4]
  assign _T_33887 = io_inAddr_21 == 6'h2a; // @[Switch.scala 30:53:@13597.4]
  assign valid_42_21 = io_inValid_21 & _T_33887; // @[Switch.scala 30:36:@13598.4]
  assign _T_33890 = io_inAddr_22 == 6'h2a; // @[Switch.scala 30:53:@13600.4]
  assign valid_42_22 = io_inValid_22 & _T_33890; // @[Switch.scala 30:36:@13601.4]
  assign _T_33893 = io_inAddr_23 == 6'h2a; // @[Switch.scala 30:53:@13603.4]
  assign valid_42_23 = io_inValid_23 & _T_33893; // @[Switch.scala 30:36:@13604.4]
  assign _T_33896 = io_inAddr_24 == 6'h2a; // @[Switch.scala 30:53:@13606.4]
  assign valid_42_24 = io_inValid_24 & _T_33896; // @[Switch.scala 30:36:@13607.4]
  assign _T_33899 = io_inAddr_25 == 6'h2a; // @[Switch.scala 30:53:@13609.4]
  assign valid_42_25 = io_inValid_25 & _T_33899; // @[Switch.scala 30:36:@13610.4]
  assign _T_33902 = io_inAddr_26 == 6'h2a; // @[Switch.scala 30:53:@13612.4]
  assign valid_42_26 = io_inValid_26 & _T_33902; // @[Switch.scala 30:36:@13613.4]
  assign _T_33905 = io_inAddr_27 == 6'h2a; // @[Switch.scala 30:53:@13615.4]
  assign valid_42_27 = io_inValid_27 & _T_33905; // @[Switch.scala 30:36:@13616.4]
  assign _T_33908 = io_inAddr_28 == 6'h2a; // @[Switch.scala 30:53:@13618.4]
  assign valid_42_28 = io_inValid_28 & _T_33908; // @[Switch.scala 30:36:@13619.4]
  assign _T_33911 = io_inAddr_29 == 6'h2a; // @[Switch.scala 30:53:@13621.4]
  assign valid_42_29 = io_inValid_29 & _T_33911; // @[Switch.scala 30:36:@13622.4]
  assign _T_33914 = io_inAddr_30 == 6'h2a; // @[Switch.scala 30:53:@13624.4]
  assign valid_42_30 = io_inValid_30 & _T_33914; // @[Switch.scala 30:36:@13625.4]
  assign _T_33917 = io_inAddr_31 == 6'h2a; // @[Switch.scala 30:53:@13627.4]
  assign valid_42_31 = io_inValid_31 & _T_33917; // @[Switch.scala 30:36:@13628.4]
  assign _T_33920 = io_inAddr_32 == 6'h2a; // @[Switch.scala 30:53:@13630.4]
  assign valid_42_32 = io_inValid_32 & _T_33920; // @[Switch.scala 30:36:@13631.4]
  assign _T_33923 = io_inAddr_33 == 6'h2a; // @[Switch.scala 30:53:@13633.4]
  assign valid_42_33 = io_inValid_33 & _T_33923; // @[Switch.scala 30:36:@13634.4]
  assign _T_33926 = io_inAddr_34 == 6'h2a; // @[Switch.scala 30:53:@13636.4]
  assign valid_42_34 = io_inValid_34 & _T_33926; // @[Switch.scala 30:36:@13637.4]
  assign _T_33929 = io_inAddr_35 == 6'h2a; // @[Switch.scala 30:53:@13639.4]
  assign valid_42_35 = io_inValid_35 & _T_33929; // @[Switch.scala 30:36:@13640.4]
  assign _T_33932 = io_inAddr_36 == 6'h2a; // @[Switch.scala 30:53:@13642.4]
  assign valid_42_36 = io_inValid_36 & _T_33932; // @[Switch.scala 30:36:@13643.4]
  assign _T_33935 = io_inAddr_37 == 6'h2a; // @[Switch.scala 30:53:@13645.4]
  assign valid_42_37 = io_inValid_37 & _T_33935; // @[Switch.scala 30:36:@13646.4]
  assign _T_33938 = io_inAddr_38 == 6'h2a; // @[Switch.scala 30:53:@13648.4]
  assign valid_42_38 = io_inValid_38 & _T_33938; // @[Switch.scala 30:36:@13649.4]
  assign _T_33941 = io_inAddr_39 == 6'h2a; // @[Switch.scala 30:53:@13651.4]
  assign valid_42_39 = io_inValid_39 & _T_33941; // @[Switch.scala 30:36:@13652.4]
  assign _T_33944 = io_inAddr_40 == 6'h2a; // @[Switch.scala 30:53:@13654.4]
  assign valid_42_40 = io_inValid_40 & _T_33944; // @[Switch.scala 30:36:@13655.4]
  assign _T_33947 = io_inAddr_41 == 6'h2a; // @[Switch.scala 30:53:@13657.4]
  assign valid_42_41 = io_inValid_41 & _T_33947; // @[Switch.scala 30:36:@13658.4]
  assign _T_33950 = io_inAddr_42 == 6'h2a; // @[Switch.scala 30:53:@13660.4]
  assign valid_42_42 = io_inValid_42 & _T_33950; // @[Switch.scala 30:36:@13661.4]
  assign _T_33953 = io_inAddr_43 == 6'h2a; // @[Switch.scala 30:53:@13663.4]
  assign valid_42_43 = io_inValid_43 & _T_33953; // @[Switch.scala 30:36:@13664.4]
  assign _T_33956 = io_inAddr_44 == 6'h2a; // @[Switch.scala 30:53:@13666.4]
  assign valid_42_44 = io_inValid_44 & _T_33956; // @[Switch.scala 30:36:@13667.4]
  assign _T_33959 = io_inAddr_45 == 6'h2a; // @[Switch.scala 30:53:@13669.4]
  assign valid_42_45 = io_inValid_45 & _T_33959; // @[Switch.scala 30:36:@13670.4]
  assign _T_33962 = io_inAddr_46 == 6'h2a; // @[Switch.scala 30:53:@13672.4]
  assign valid_42_46 = io_inValid_46 & _T_33962; // @[Switch.scala 30:36:@13673.4]
  assign _T_33965 = io_inAddr_47 == 6'h2a; // @[Switch.scala 30:53:@13675.4]
  assign valid_42_47 = io_inValid_47 & _T_33965; // @[Switch.scala 30:36:@13676.4]
  assign _T_33968 = io_inAddr_48 == 6'h2a; // @[Switch.scala 30:53:@13678.4]
  assign valid_42_48 = io_inValid_48 & _T_33968; // @[Switch.scala 30:36:@13679.4]
  assign _T_33971 = io_inAddr_49 == 6'h2a; // @[Switch.scala 30:53:@13681.4]
  assign valid_42_49 = io_inValid_49 & _T_33971; // @[Switch.scala 30:36:@13682.4]
  assign _T_33974 = io_inAddr_50 == 6'h2a; // @[Switch.scala 30:53:@13684.4]
  assign valid_42_50 = io_inValid_50 & _T_33974; // @[Switch.scala 30:36:@13685.4]
  assign _T_33977 = io_inAddr_51 == 6'h2a; // @[Switch.scala 30:53:@13687.4]
  assign valid_42_51 = io_inValid_51 & _T_33977; // @[Switch.scala 30:36:@13688.4]
  assign _T_33980 = io_inAddr_52 == 6'h2a; // @[Switch.scala 30:53:@13690.4]
  assign valid_42_52 = io_inValid_52 & _T_33980; // @[Switch.scala 30:36:@13691.4]
  assign _T_33983 = io_inAddr_53 == 6'h2a; // @[Switch.scala 30:53:@13693.4]
  assign valid_42_53 = io_inValid_53 & _T_33983; // @[Switch.scala 30:36:@13694.4]
  assign _T_33986 = io_inAddr_54 == 6'h2a; // @[Switch.scala 30:53:@13696.4]
  assign valid_42_54 = io_inValid_54 & _T_33986; // @[Switch.scala 30:36:@13697.4]
  assign _T_33989 = io_inAddr_55 == 6'h2a; // @[Switch.scala 30:53:@13699.4]
  assign valid_42_55 = io_inValid_55 & _T_33989; // @[Switch.scala 30:36:@13700.4]
  assign _T_33992 = io_inAddr_56 == 6'h2a; // @[Switch.scala 30:53:@13702.4]
  assign valid_42_56 = io_inValid_56 & _T_33992; // @[Switch.scala 30:36:@13703.4]
  assign _T_33995 = io_inAddr_57 == 6'h2a; // @[Switch.scala 30:53:@13705.4]
  assign valid_42_57 = io_inValid_57 & _T_33995; // @[Switch.scala 30:36:@13706.4]
  assign _T_33998 = io_inAddr_58 == 6'h2a; // @[Switch.scala 30:53:@13708.4]
  assign valid_42_58 = io_inValid_58 & _T_33998; // @[Switch.scala 30:36:@13709.4]
  assign _T_34001 = io_inAddr_59 == 6'h2a; // @[Switch.scala 30:53:@13711.4]
  assign valid_42_59 = io_inValid_59 & _T_34001; // @[Switch.scala 30:36:@13712.4]
  assign _T_34004 = io_inAddr_60 == 6'h2a; // @[Switch.scala 30:53:@13714.4]
  assign valid_42_60 = io_inValid_60 & _T_34004; // @[Switch.scala 30:36:@13715.4]
  assign _T_34007 = io_inAddr_61 == 6'h2a; // @[Switch.scala 30:53:@13717.4]
  assign valid_42_61 = io_inValid_61 & _T_34007; // @[Switch.scala 30:36:@13718.4]
  assign _T_34010 = io_inAddr_62 == 6'h2a; // @[Switch.scala 30:53:@13720.4]
  assign valid_42_62 = io_inValid_62 & _T_34010; // @[Switch.scala 30:36:@13721.4]
  assign _T_34013 = io_inAddr_63 == 6'h2a; // @[Switch.scala 30:53:@13723.4]
  assign valid_42_63 = io_inValid_63 & _T_34013; // @[Switch.scala 30:36:@13724.4]
  assign _T_34079 = valid_42_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@13726.4]
  assign _T_34080 = valid_42_61 ? 6'h3d : _T_34079; // @[Mux.scala 31:69:@13727.4]
  assign _T_34081 = valid_42_60 ? 6'h3c : _T_34080; // @[Mux.scala 31:69:@13728.4]
  assign _T_34082 = valid_42_59 ? 6'h3b : _T_34081; // @[Mux.scala 31:69:@13729.4]
  assign _T_34083 = valid_42_58 ? 6'h3a : _T_34082; // @[Mux.scala 31:69:@13730.4]
  assign _T_34084 = valid_42_57 ? 6'h39 : _T_34083; // @[Mux.scala 31:69:@13731.4]
  assign _T_34085 = valid_42_56 ? 6'h38 : _T_34084; // @[Mux.scala 31:69:@13732.4]
  assign _T_34086 = valid_42_55 ? 6'h37 : _T_34085; // @[Mux.scala 31:69:@13733.4]
  assign _T_34087 = valid_42_54 ? 6'h36 : _T_34086; // @[Mux.scala 31:69:@13734.4]
  assign _T_34088 = valid_42_53 ? 6'h35 : _T_34087; // @[Mux.scala 31:69:@13735.4]
  assign _T_34089 = valid_42_52 ? 6'h34 : _T_34088; // @[Mux.scala 31:69:@13736.4]
  assign _T_34090 = valid_42_51 ? 6'h33 : _T_34089; // @[Mux.scala 31:69:@13737.4]
  assign _T_34091 = valid_42_50 ? 6'h32 : _T_34090; // @[Mux.scala 31:69:@13738.4]
  assign _T_34092 = valid_42_49 ? 6'h31 : _T_34091; // @[Mux.scala 31:69:@13739.4]
  assign _T_34093 = valid_42_48 ? 6'h30 : _T_34092; // @[Mux.scala 31:69:@13740.4]
  assign _T_34094 = valid_42_47 ? 6'h2f : _T_34093; // @[Mux.scala 31:69:@13741.4]
  assign _T_34095 = valid_42_46 ? 6'h2e : _T_34094; // @[Mux.scala 31:69:@13742.4]
  assign _T_34096 = valid_42_45 ? 6'h2d : _T_34095; // @[Mux.scala 31:69:@13743.4]
  assign _T_34097 = valid_42_44 ? 6'h2c : _T_34096; // @[Mux.scala 31:69:@13744.4]
  assign _T_34098 = valid_42_43 ? 6'h2b : _T_34097; // @[Mux.scala 31:69:@13745.4]
  assign _T_34099 = valid_42_42 ? 6'h2a : _T_34098; // @[Mux.scala 31:69:@13746.4]
  assign _T_34100 = valid_42_41 ? 6'h29 : _T_34099; // @[Mux.scala 31:69:@13747.4]
  assign _T_34101 = valid_42_40 ? 6'h28 : _T_34100; // @[Mux.scala 31:69:@13748.4]
  assign _T_34102 = valid_42_39 ? 6'h27 : _T_34101; // @[Mux.scala 31:69:@13749.4]
  assign _T_34103 = valid_42_38 ? 6'h26 : _T_34102; // @[Mux.scala 31:69:@13750.4]
  assign _T_34104 = valid_42_37 ? 6'h25 : _T_34103; // @[Mux.scala 31:69:@13751.4]
  assign _T_34105 = valid_42_36 ? 6'h24 : _T_34104; // @[Mux.scala 31:69:@13752.4]
  assign _T_34106 = valid_42_35 ? 6'h23 : _T_34105; // @[Mux.scala 31:69:@13753.4]
  assign _T_34107 = valid_42_34 ? 6'h22 : _T_34106; // @[Mux.scala 31:69:@13754.4]
  assign _T_34108 = valid_42_33 ? 6'h21 : _T_34107; // @[Mux.scala 31:69:@13755.4]
  assign _T_34109 = valid_42_32 ? 6'h20 : _T_34108; // @[Mux.scala 31:69:@13756.4]
  assign _T_34110 = valid_42_31 ? 6'h1f : _T_34109; // @[Mux.scala 31:69:@13757.4]
  assign _T_34111 = valid_42_30 ? 6'h1e : _T_34110; // @[Mux.scala 31:69:@13758.4]
  assign _T_34112 = valid_42_29 ? 6'h1d : _T_34111; // @[Mux.scala 31:69:@13759.4]
  assign _T_34113 = valid_42_28 ? 6'h1c : _T_34112; // @[Mux.scala 31:69:@13760.4]
  assign _T_34114 = valid_42_27 ? 6'h1b : _T_34113; // @[Mux.scala 31:69:@13761.4]
  assign _T_34115 = valid_42_26 ? 6'h1a : _T_34114; // @[Mux.scala 31:69:@13762.4]
  assign _T_34116 = valid_42_25 ? 6'h19 : _T_34115; // @[Mux.scala 31:69:@13763.4]
  assign _T_34117 = valid_42_24 ? 6'h18 : _T_34116; // @[Mux.scala 31:69:@13764.4]
  assign _T_34118 = valid_42_23 ? 6'h17 : _T_34117; // @[Mux.scala 31:69:@13765.4]
  assign _T_34119 = valid_42_22 ? 6'h16 : _T_34118; // @[Mux.scala 31:69:@13766.4]
  assign _T_34120 = valid_42_21 ? 6'h15 : _T_34119; // @[Mux.scala 31:69:@13767.4]
  assign _T_34121 = valid_42_20 ? 6'h14 : _T_34120; // @[Mux.scala 31:69:@13768.4]
  assign _T_34122 = valid_42_19 ? 6'h13 : _T_34121; // @[Mux.scala 31:69:@13769.4]
  assign _T_34123 = valid_42_18 ? 6'h12 : _T_34122; // @[Mux.scala 31:69:@13770.4]
  assign _T_34124 = valid_42_17 ? 6'h11 : _T_34123; // @[Mux.scala 31:69:@13771.4]
  assign _T_34125 = valid_42_16 ? 6'h10 : _T_34124; // @[Mux.scala 31:69:@13772.4]
  assign _T_34126 = valid_42_15 ? 6'hf : _T_34125; // @[Mux.scala 31:69:@13773.4]
  assign _T_34127 = valid_42_14 ? 6'he : _T_34126; // @[Mux.scala 31:69:@13774.4]
  assign _T_34128 = valid_42_13 ? 6'hd : _T_34127; // @[Mux.scala 31:69:@13775.4]
  assign _T_34129 = valid_42_12 ? 6'hc : _T_34128; // @[Mux.scala 31:69:@13776.4]
  assign _T_34130 = valid_42_11 ? 6'hb : _T_34129; // @[Mux.scala 31:69:@13777.4]
  assign _T_34131 = valid_42_10 ? 6'ha : _T_34130; // @[Mux.scala 31:69:@13778.4]
  assign _T_34132 = valid_42_9 ? 6'h9 : _T_34131; // @[Mux.scala 31:69:@13779.4]
  assign _T_34133 = valid_42_8 ? 6'h8 : _T_34132; // @[Mux.scala 31:69:@13780.4]
  assign _T_34134 = valid_42_7 ? 6'h7 : _T_34133; // @[Mux.scala 31:69:@13781.4]
  assign _T_34135 = valid_42_6 ? 6'h6 : _T_34134; // @[Mux.scala 31:69:@13782.4]
  assign _T_34136 = valid_42_5 ? 6'h5 : _T_34135; // @[Mux.scala 31:69:@13783.4]
  assign _T_34137 = valid_42_4 ? 6'h4 : _T_34136; // @[Mux.scala 31:69:@13784.4]
  assign _T_34138 = valid_42_3 ? 6'h3 : _T_34137; // @[Mux.scala 31:69:@13785.4]
  assign _T_34139 = valid_42_2 ? 6'h2 : _T_34138; // @[Mux.scala 31:69:@13786.4]
  assign _T_34140 = valid_42_1 ? 6'h1 : _T_34139; // @[Mux.scala 31:69:@13787.4]
  assign select_42 = valid_42_0 ? 6'h0 : _T_34140; // @[Mux.scala 31:69:@13788.4]
  assign _GEN_2689 = 6'h1 == select_42 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2690 = 6'h2 == select_42 ? io_inData_2 : _GEN_2689; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2691 = 6'h3 == select_42 ? io_inData_3 : _GEN_2690; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2692 = 6'h4 == select_42 ? io_inData_4 : _GEN_2691; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2693 = 6'h5 == select_42 ? io_inData_5 : _GEN_2692; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2694 = 6'h6 == select_42 ? io_inData_6 : _GEN_2693; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2695 = 6'h7 == select_42 ? io_inData_7 : _GEN_2694; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2696 = 6'h8 == select_42 ? io_inData_8 : _GEN_2695; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2697 = 6'h9 == select_42 ? io_inData_9 : _GEN_2696; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2698 = 6'ha == select_42 ? io_inData_10 : _GEN_2697; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2699 = 6'hb == select_42 ? io_inData_11 : _GEN_2698; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2700 = 6'hc == select_42 ? io_inData_12 : _GEN_2699; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2701 = 6'hd == select_42 ? io_inData_13 : _GEN_2700; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2702 = 6'he == select_42 ? io_inData_14 : _GEN_2701; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2703 = 6'hf == select_42 ? io_inData_15 : _GEN_2702; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2704 = 6'h10 == select_42 ? io_inData_16 : _GEN_2703; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2705 = 6'h11 == select_42 ? io_inData_17 : _GEN_2704; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2706 = 6'h12 == select_42 ? io_inData_18 : _GEN_2705; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2707 = 6'h13 == select_42 ? io_inData_19 : _GEN_2706; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2708 = 6'h14 == select_42 ? io_inData_20 : _GEN_2707; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2709 = 6'h15 == select_42 ? io_inData_21 : _GEN_2708; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2710 = 6'h16 == select_42 ? io_inData_22 : _GEN_2709; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2711 = 6'h17 == select_42 ? io_inData_23 : _GEN_2710; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2712 = 6'h18 == select_42 ? io_inData_24 : _GEN_2711; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2713 = 6'h19 == select_42 ? io_inData_25 : _GEN_2712; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2714 = 6'h1a == select_42 ? io_inData_26 : _GEN_2713; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2715 = 6'h1b == select_42 ? io_inData_27 : _GEN_2714; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2716 = 6'h1c == select_42 ? io_inData_28 : _GEN_2715; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2717 = 6'h1d == select_42 ? io_inData_29 : _GEN_2716; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2718 = 6'h1e == select_42 ? io_inData_30 : _GEN_2717; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2719 = 6'h1f == select_42 ? io_inData_31 : _GEN_2718; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2720 = 6'h20 == select_42 ? io_inData_32 : _GEN_2719; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2721 = 6'h21 == select_42 ? io_inData_33 : _GEN_2720; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2722 = 6'h22 == select_42 ? io_inData_34 : _GEN_2721; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2723 = 6'h23 == select_42 ? io_inData_35 : _GEN_2722; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2724 = 6'h24 == select_42 ? io_inData_36 : _GEN_2723; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2725 = 6'h25 == select_42 ? io_inData_37 : _GEN_2724; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2726 = 6'h26 == select_42 ? io_inData_38 : _GEN_2725; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2727 = 6'h27 == select_42 ? io_inData_39 : _GEN_2726; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2728 = 6'h28 == select_42 ? io_inData_40 : _GEN_2727; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2729 = 6'h29 == select_42 ? io_inData_41 : _GEN_2728; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2730 = 6'h2a == select_42 ? io_inData_42 : _GEN_2729; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2731 = 6'h2b == select_42 ? io_inData_43 : _GEN_2730; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2732 = 6'h2c == select_42 ? io_inData_44 : _GEN_2731; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2733 = 6'h2d == select_42 ? io_inData_45 : _GEN_2732; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2734 = 6'h2e == select_42 ? io_inData_46 : _GEN_2733; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2735 = 6'h2f == select_42 ? io_inData_47 : _GEN_2734; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2736 = 6'h30 == select_42 ? io_inData_48 : _GEN_2735; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2737 = 6'h31 == select_42 ? io_inData_49 : _GEN_2736; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2738 = 6'h32 == select_42 ? io_inData_50 : _GEN_2737; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2739 = 6'h33 == select_42 ? io_inData_51 : _GEN_2738; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2740 = 6'h34 == select_42 ? io_inData_52 : _GEN_2739; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2741 = 6'h35 == select_42 ? io_inData_53 : _GEN_2740; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2742 = 6'h36 == select_42 ? io_inData_54 : _GEN_2741; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2743 = 6'h37 == select_42 ? io_inData_55 : _GEN_2742; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2744 = 6'h38 == select_42 ? io_inData_56 : _GEN_2743; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2745 = 6'h39 == select_42 ? io_inData_57 : _GEN_2744; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2746 = 6'h3a == select_42 ? io_inData_58 : _GEN_2745; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2747 = 6'h3b == select_42 ? io_inData_59 : _GEN_2746; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2748 = 6'h3c == select_42 ? io_inData_60 : _GEN_2747; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2749 = 6'h3d == select_42 ? io_inData_61 : _GEN_2748; // @[Switch.scala 33:19:@13790.4]
  assign _GEN_2750 = 6'h3e == select_42 ? io_inData_62 : _GEN_2749; // @[Switch.scala 33:19:@13790.4]
  assign _T_34149 = {valid_42_7,valid_42_6,valid_42_5,valid_42_4,valid_42_3,valid_42_2,valid_42_1,valid_42_0}; // @[Switch.scala 34:32:@13797.4]
  assign _T_34157 = {valid_42_15,valid_42_14,valid_42_13,valid_42_12,valid_42_11,valid_42_10,valid_42_9,valid_42_8,_T_34149}; // @[Switch.scala 34:32:@13805.4]
  assign _T_34164 = {valid_42_23,valid_42_22,valid_42_21,valid_42_20,valid_42_19,valid_42_18,valid_42_17,valid_42_16}; // @[Switch.scala 34:32:@13812.4]
  assign _T_34173 = {valid_42_31,valid_42_30,valid_42_29,valid_42_28,valid_42_27,valid_42_26,valid_42_25,valid_42_24,_T_34164,_T_34157}; // @[Switch.scala 34:32:@13821.4]
  assign _T_34180 = {valid_42_39,valid_42_38,valid_42_37,valid_42_36,valid_42_35,valid_42_34,valid_42_33,valid_42_32}; // @[Switch.scala 34:32:@13828.4]
  assign _T_34188 = {valid_42_47,valid_42_46,valid_42_45,valid_42_44,valid_42_43,valid_42_42,valid_42_41,valid_42_40,_T_34180}; // @[Switch.scala 34:32:@13836.4]
  assign _T_34195 = {valid_42_55,valid_42_54,valid_42_53,valid_42_52,valid_42_51,valid_42_50,valid_42_49,valid_42_48}; // @[Switch.scala 34:32:@13843.4]
  assign _T_34204 = {valid_42_63,valid_42_62,valid_42_61,valid_42_60,valid_42_59,valid_42_58,valid_42_57,valid_42_56,_T_34195,_T_34188}; // @[Switch.scala 34:32:@13852.4]
  assign _T_34205 = {_T_34204,_T_34173}; // @[Switch.scala 34:32:@13853.4]
  assign _T_34209 = io_inAddr_0 == 6'h2b; // @[Switch.scala 30:53:@13856.4]
  assign valid_43_0 = io_inValid_0 & _T_34209; // @[Switch.scala 30:36:@13857.4]
  assign _T_34212 = io_inAddr_1 == 6'h2b; // @[Switch.scala 30:53:@13859.4]
  assign valid_43_1 = io_inValid_1 & _T_34212; // @[Switch.scala 30:36:@13860.4]
  assign _T_34215 = io_inAddr_2 == 6'h2b; // @[Switch.scala 30:53:@13862.4]
  assign valid_43_2 = io_inValid_2 & _T_34215; // @[Switch.scala 30:36:@13863.4]
  assign _T_34218 = io_inAddr_3 == 6'h2b; // @[Switch.scala 30:53:@13865.4]
  assign valid_43_3 = io_inValid_3 & _T_34218; // @[Switch.scala 30:36:@13866.4]
  assign _T_34221 = io_inAddr_4 == 6'h2b; // @[Switch.scala 30:53:@13868.4]
  assign valid_43_4 = io_inValid_4 & _T_34221; // @[Switch.scala 30:36:@13869.4]
  assign _T_34224 = io_inAddr_5 == 6'h2b; // @[Switch.scala 30:53:@13871.4]
  assign valid_43_5 = io_inValid_5 & _T_34224; // @[Switch.scala 30:36:@13872.4]
  assign _T_34227 = io_inAddr_6 == 6'h2b; // @[Switch.scala 30:53:@13874.4]
  assign valid_43_6 = io_inValid_6 & _T_34227; // @[Switch.scala 30:36:@13875.4]
  assign _T_34230 = io_inAddr_7 == 6'h2b; // @[Switch.scala 30:53:@13877.4]
  assign valid_43_7 = io_inValid_7 & _T_34230; // @[Switch.scala 30:36:@13878.4]
  assign _T_34233 = io_inAddr_8 == 6'h2b; // @[Switch.scala 30:53:@13880.4]
  assign valid_43_8 = io_inValid_8 & _T_34233; // @[Switch.scala 30:36:@13881.4]
  assign _T_34236 = io_inAddr_9 == 6'h2b; // @[Switch.scala 30:53:@13883.4]
  assign valid_43_9 = io_inValid_9 & _T_34236; // @[Switch.scala 30:36:@13884.4]
  assign _T_34239 = io_inAddr_10 == 6'h2b; // @[Switch.scala 30:53:@13886.4]
  assign valid_43_10 = io_inValid_10 & _T_34239; // @[Switch.scala 30:36:@13887.4]
  assign _T_34242 = io_inAddr_11 == 6'h2b; // @[Switch.scala 30:53:@13889.4]
  assign valid_43_11 = io_inValid_11 & _T_34242; // @[Switch.scala 30:36:@13890.4]
  assign _T_34245 = io_inAddr_12 == 6'h2b; // @[Switch.scala 30:53:@13892.4]
  assign valid_43_12 = io_inValid_12 & _T_34245; // @[Switch.scala 30:36:@13893.4]
  assign _T_34248 = io_inAddr_13 == 6'h2b; // @[Switch.scala 30:53:@13895.4]
  assign valid_43_13 = io_inValid_13 & _T_34248; // @[Switch.scala 30:36:@13896.4]
  assign _T_34251 = io_inAddr_14 == 6'h2b; // @[Switch.scala 30:53:@13898.4]
  assign valid_43_14 = io_inValid_14 & _T_34251; // @[Switch.scala 30:36:@13899.4]
  assign _T_34254 = io_inAddr_15 == 6'h2b; // @[Switch.scala 30:53:@13901.4]
  assign valid_43_15 = io_inValid_15 & _T_34254; // @[Switch.scala 30:36:@13902.4]
  assign _T_34257 = io_inAddr_16 == 6'h2b; // @[Switch.scala 30:53:@13904.4]
  assign valid_43_16 = io_inValid_16 & _T_34257; // @[Switch.scala 30:36:@13905.4]
  assign _T_34260 = io_inAddr_17 == 6'h2b; // @[Switch.scala 30:53:@13907.4]
  assign valid_43_17 = io_inValid_17 & _T_34260; // @[Switch.scala 30:36:@13908.4]
  assign _T_34263 = io_inAddr_18 == 6'h2b; // @[Switch.scala 30:53:@13910.4]
  assign valid_43_18 = io_inValid_18 & _T_34263; // @[Switch.scala 30:36:@13911.4]
  assign _T_34266 = io_inAddr_19 == 6'h2b; // @[Switch.scala 30:53:@13913.4]
  assign valid_43_19 = io_inValid_19 & _T_34266; // @[Switch.scala 30:36:@13914.4]
  assign _T_34269 = io_inAddr_20 == 6'h2b; // @[Switch.scala 30:53:@13916.4]
  assign valid_43_20 = io_inValid_20 & _T_34269; // @[Switch.scala 30:36:@13917.4]
  assign _T_34272 = io_inAddr_21 == 6'h2b; // @[Switch.scala 30:53:@13919.4]
  assign valid_43_21 = io_inValid_21 & _T_34272; // @[Switch.scala 30:36:@13920.4]
  assign _T_34275 = io_inAddr_22 == 6'h2b; // @[Switch.scala 30:53:@13922.4]
  assign valid_43_22 = io_inValid_22 & _T_34275; // @[Switch.scala 30:36:@13923.4]
  assign _T_34278 = io_inAddr_23 == 6'h2b; // @[Switch.scala 30:53:@13925.4]
  assign valid_43_23 = io_inValid_23 & _T_34278; // @[Switch.scala 30:36:@13926.4]
  assign _T_34281 = io_inAddr_24 == 6'h2b; // @[Switch.scala 30:53:@13928.4]
  assign valid_43_24 = io_inValid_24 & _T_34281; // @[Switch.scala 30:36:@13929.4]
  assign _T_34284 = io_inAddr_25 == 6'h2b; // @[Switch.scala 30:53:@13931.4]
  assign valid_43_25 = io_inValid_25 & _T_34284; // @[Switch.scala 30:36:@13932.4]
  assign _T_34287 = io_inAddr_26 == 6'h2b; // @[Switch.scala 30:53:@13934.4]
  assign valid_43_26 = io_inValid_26 & _T_34287; // @[Switch.scala 30:36:@13935.4]
  assign _T_34290 = io_inAddr_27 == 6'h2b; // @[Switch.scala 30:53:@13937.4]
  assign valid_43_27 = io_inValid_27 & _T_34290; // @[Switch.scala 30:36:@13938.4]
  assign _T_34293 = io_inAddr_28 == 6'h2b; // @[Switch.scala 30:53:@13940.4]
  assign valid_43_28 = io_inValid_28 & _T_34293; // @[Switch.scala 30:36:@13941.4]
  assign _T_34296 = io_inAddr_29 == 6'h2b; // @[Switch.scala 30:53:@13943.4]
  assign valid_43_29 = io_inValid_29 & _T_34296; // @[Switch.scala 30:36:@13944.4]
  assign _T_34299 = io_inAddr_30 == 6'h2b; // @[Switch.scala 30:53:@13946.4]
  assign valid_43_30 = io_inValid_30 & _T_34299; // @[Switch.scala 30:36:@13947.4]
  assign _T_34302 = io_inAddr_31 == 6'h2b; // @[Switch.scala 30:53:@13949.4]
  assign valid_43_31 = io_inValid_31 & _T_34302; // @[Switch.scala 30:36:@13950.4]
  assign _T_34305 = io_inAddr_32 == 6'h2b; // @[Switch.scala 30:53:@13952.4]
  assign valid_43_32 = io_inValid_32 & _T_34305; // @[Switch.scala 30:36:@13953.4]
  assign _T_34308 = io_inAddr_33 == 6'h2b; // @[Switch.scala 30:53:@13955.4]
  assign valid_43_33 = io_inValid_33 & _T_34308; // @[Switch.scala 30:36:@13956.4]
  assign _T_34311 = io_inAddr_34 == 6'h2b; // @[Switch.scala 30:53:@13958.4]
  assign valid_43_34 = io_inValid_34 & _T_34311; // @[Switch.scala 30:36:@13959.4]
  assign _T_34314 = io_inAddr_35 == 6'h2b; // @[Switch.scala 30:53:@13961.4]
  assign valid_43_35 = io_inValid_35 & _T_34314; // @[Switch.scala 30:36:@13962.4]
  assign _T_34317 = io_inAddr_36 == 6'h2b; // @[Switch.scala 30:53:@13964.4]
  assign valid_43_36 = io_inValid_36 & _T_34317; // @[Switch.scala 30:36:@13965.4]
  assign _T_34320 = io_inAddr_37 == 6'h2b; // @[Switch.scala 30:53:@13967.4]
  assign valid_43_37 = io_inValid_37 & _T_34320; // @[Switch.scala 30:36:@13968.4]
  assign _T_34323 = io_inAddr_38 == 6'h2b; // @[Switch.scala 30:53:@13970.4]
  assign valid_43_38 = io_inValid_38 & _T_34323; // @[Switch.scala 30:36:@13971.4]
  assign _T_34326 = io_inAddr_39 == 6'h2b; // @[Switch.scala 30:53:@13973.4]
  assign valid_43_39 = io_inValid_39 & _T_34326; // @[Switch.scala 30:36:@13974.4]
  assign _T_34329 = io_inAddr_40 == 6'h2b; // @[Switch.scala 30:53:@13976.4]
  assign valid_43_40 = io_inValid_40 & _T_34329; // @[Switch.scala 30:36:@13977.4]
  assign _T_34332 = io_inAddr_41 == 6'h2b; // @[Switch.scala 30:53:@13979.4]
  assign valid_43_41 = io_inValid_41 & _T_34332; // @[Switch.scala 30:36:@13980.4]
  assign _T_34335 = io_inAddr_42 == 6'h2b; // @[Switch.scala 30:53:@13982.4]
  assign valid_43_42 = io_inValid_42 & _T_34335; // @[Switch.scala 30:36:@13983.4]
  assign _T_34338 = io_inAddr_43 == 6'h2b; // @[Switch.scala 30:53:@13985.4]
  assign valid_43_43 = io_inValid_43 & _T_34338; // @[Switch.scala 30:36:@13986.4]
  assign _T_34341 = io_inAddr_44 == 6'h2b; // @[Switch.scala 30:53:@13988.4]
  assign valid_43_44 = io_inValid_44 & _T_34341; // @[Switch.scala 30:36:@13989.4]
  assign _T_34344 = io_inAddr_45 == 6'h2b; // @[Switch.scala 30:53:@13991.4]
  assign valid_43_45 = io_inValid_45 & _T_34344; // @[Switch.scala 30:36:@13992.4]
  assign _T_34347 = io_inAddr_46 == 6'h2b; // @[Switch.scala 30:53:@13994.4]
  assign valid_43_46 = io_inValid_46 & _T_34347; // @[Switch.scala 30:36:@13995.4]
  assign _T_34350 = io_inAddr_47 == 6'h2b; // @[Switch.scala 30:53:@13997.4]
  assign valid_43_47 = io_inValid_47 & _T_34350; // @[Switch.scala 30:36:@13998.4]
  assign _T_34353 = io_inAddr_48 == 6'h2b; // @[Switch.scala 30:53:@14000.4]
  assign valid_43_48 = io_inValid_48 & _T_34353; // @[Switch.scala 30:36:@14001.4]
  assign _T_34356 = io_inAddr_49 == 6'h2b; // @[Switch.scala 30:53:@14003.4]
  assign valid_43_49 = io_inValid_49 & _T_34356; // @[Switch.scala 30:36:@14004.4]
  assign _T_34359 = io_inAddr_50 == 6'h2b; // @[Switch.scala 30:53:@14006.4]
  assign valid_43_50 = io_inValid_50 & _T_34359; // @[Switch.scala 30:36:@14007.4]
  assign _T_34362 = io_inAddr_51 == 6'h2b; // @[Switch.scala 30:53:@14009.4]
  assign valid_43_51 = io_inValid_51 & _T_34362; // @[Switch.scala 30:36:@14010.4]
  assign _T_34365 = io_inAddr_52 == 6'h2b; // @[Switch.scala 30:53:@14012.4]
  assign valid_43_52 = io_inValid_52 & _T_34365; // @[Switch.scala 30:36:@14013.4]
  assign _T_34368 = io_inAddr_53 == 6'h2b; // @[Switch.scala 30:53:@14015.4]
  assign valid_43_53 = io_inValid_53 & _T_34368; // @[Switch.scala 30:36:@14016.4]
  assign _T_34371 = io_inAddr_54 == 6'h2b; // @[Switch.scala 30:53:@14018.4]
  assign valid_43_54 = io_inValid_54 & _T_34371; // @[Switch.scala 30:36:@14019.4]
  assign _T_34374 = io_inAddr_55 == 6'h2b; // @[Switch.scala 30:53:@14021.4]
  assign valid_43_55 = io_inValid_55 & _T_34374; // @[Switch.scala 30:36:@14022.4]
  assign _T_34377 = io_inAddr_56 == 6'h2b; // @[Switch.scala 30:53:@14024.4]
  assign valid_43_56 = io_inValid_56 & _T_34377; // @[Switch.scala 30:36:@14025.4]
  assign _T_34380 = io_inAddr_57 == 6'h2b; // @[Switch.scala 30:53:@14027.4]
  assign valid_43_57 = io_inValid_57 & _T_34380; // @[Switch.scala 30:36:@14028.4]
  assign _T_34383 = io_inAddr_58 == 6'h2b; // @[Switch.scala 30:53:@14030.4]
  assign valid_43_58 = io_inValid_58 & _T_34383; // @[Switch.scala 30:36:@14031.4]
  assign _T_34386 = io_inAddr_59 == 6'h2b; // @[Switch.scala 30:53:@14033.4]
  assign valid_43_59 = io_inValid_59 & _T_34386; // @[Switch.scala 30:36:@14034.4]
  assign _T_34389 = io_inAddr_60 == 6'h2b; // @[Switch.scala 30:53:@14036.4]
  assign valid_43_60 = io_inValid_60 & _T_34389; // @[Switch.scala 30:36:@14037.4]
  assign _T_34392 = io_inAddr_61 == 6'h2b; // @[Switch.scala 30:53:@14039.4]
  assign valid_43_61 = io_inValid_61 & _T_34392; // @[Switch.scala 30:36:@14040.4]
  assign _T_34395 = io_inAddr_62 == 6'h2b; // @[Switch.scala 30:53:@14042.4]
  assign valid_43_62 = io_inValid_62 & _T_34395; // @[Switch.scala 30:36:@14043.4]
  assign _T_34398 = io_inAddr_63 == 6'h2b; // @[Switch.scala 30:53:@14045.4]
  assign valid_43_63 = io_inValid_63 & _T_34398; // @[Switch.scala 30:36:@14046.4]
  assign _T_34464 = valid_43_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@14048.4]
  assign _T_34465 = valid_43_61 ? 6'h3d : _T_34464; // @[Mux.scala 31:69:@14049.4]
  assign _T_34466 = valid_43_60 ? 6'h3c : _T_34465; // @[Mux.scala 31:69:@14050.4]
  assign _T_34467 = valid_43_59 ? 6'h3b : _T_34466; // @[Mux.scala 31:69:@14051.4]
  assign _T_34468 = valid_43_58 ? 6'h3a : _T_34467; // @[Mux.scala 31:69:@14052.4]
  assign _T_34469 = valid_43_57 ? 6'h39 : _T_34468; // @[Mux.scala 31:69:@14053.4]
  assign _T_34470 = valid_43_56 ? 6'h38 : _T_34469; // @[Mux.scala 31:69:@14054.4]
  assign _T_34471 = valid_43_55 ? 6'h37 : _T_34470; // @[Mux.scala 31:69:@14055.4]
  assign _T_34472 = valid_43_54 ? 6'h36 : _T_34471; // @[Mux.scala 31:69:@14056.4]
  assign _T_34473 = valid_43_53 ? 6'h35 : _T_34472; // @[Mux.scala 31:69:@14057.4]
  assign _T_34474 = valid_43_52 ? 6'h34 : _T_34473; // @[Mux.scala 31:69:@14058.4]
  assign _T_34475 = valid_43_51 ? 6'h33 : _T_34474; // @[Mux.scala 31:69:@14059.4]
  assign _T_34476 = valid_43_50 ? 6'h32 : _T_34475; // @[Mux.scala 31:69:@14060.4]
  assign _T_34477 = valid_43_49 ? 6'h31 : _T_34476; // @[Mux.scala 31:69:@14061.4]
  assign _T_34478 = valid_43_48 ? 6'h30 : _T_34477; // @[Mux.scala 31:69:@14062.4]
  assign _T_34479 = valid_43_47 ? 6'h2f : _T_34478; // @[Mux.scala 31:69:@14063.4]
  assign _T_34480 = valid_43_46 ? 6'h2e : _T_34479; // @[Mux.scala 31:69:@14064.4]
  assign _T_34481 = valid_43_45 ? 6'h2d : _T_34480; // @[Mux.scala 31:69:@14065.4]
  assign _T_34482 = valid_43_44 ? 6'h2c : _T_34481; // @[Mux.scala 31:69:@14066.4]
  assign _T_34483 = valid_43_43 ? 6'h2b : _T_34482; // @[Mux.scala 31:69:@14067.4]
  assign _T_34484 = valid_43_42 ? 6'h2a : _T_34483; // @[Mux.scala 31:69:@14068.4]
  assign _T_34485 = valid_43_41 ? 6'h29 : _T_34484; // @[Mux.scala 31:69:@14069.4]
  assign _T_34486 = valid_43_40 ? 6'h28 : _T_34485; // @[Mux.scala 31:69:@14070.4]
  assign _T_34487 = valid_43_39 ? 6'h27 : _T_34486; // @[Mux.scala 31:69:@14071.4]
  assign _T_34488 = valid_43_38 ? 6'h26 : _T_34487; // @[Mux.scala 31:69:@14072.4]
  assign _T_34489 = valid_43_37 ? 6'h25 : _T_34488; // @[Mux.scala 31:69:@14073.4]
  assign _T_34490 = valid_43_36 ? 6'h24 : _T_34489; // @[Mux.scala 31:69:@14074.4]
  assign _T_34491 = valid_43_35 ? 6'h23 : _T_34490; // @[Mux.scala 31:69:@14075.4]
  assign _T_34492 = valid_43_34 ? 6'h22 : _T_34491; // @[Mux.scala 31:69:@14076.4]
  assign _T_34493 = valid_43_33 ? 6'h21 : _T_34492; // @[Mux.scala 31:69:@14077.4]
  assign _T_34494 = valid_43_32 ? 6'h20 : _T_34493; // @[Mux.scala 31:69:@14078.4]
  assign _T_34495 = valid_43_31 ? 6'h1f : _T_34494; // @[Mux.scala 31:69:@14079.4]
  assign _T_34496 = valid_43_30 ? 6'h1e : _T_34495; // @[Mux.scala 31:69:@14080.4]
  assign _T_34497 = valid_43_29 ? 6'h1d : _T_34496; // @[Mux.scala 31:69:@14081.4]
  assign _T_34498 = valid_43_28 ? 6'h1c : _T_34497; // @[Mux.scala 31:69:@14082.4]
  assign _T_34499 = valid_43_27 ? 6'h1b : _T_34498; // @[Mux.scala 31:69:@14083.4]
  assign _T_34500 = valid_43_26 ? 6'h1a : _T_34499; // @[Mux.scala 31:69:@14084.4]
  assign _T_34501 = valid_43_25 ? 6'h19 : _T_34500; // @[Mux.scala 31:69:@14085.4]
  assign _T_34502 = valid_43_24 ? 6'h18 : _T_34501; // @[Mux.scala 31:69:@14086.4]
  assign _T_34503 = valid_43_23 ? 6'h17 : _T_34502; // @[Mux.scala 31:69:@14087.4]
  assign _T_34504 = valid_43_22 ? 6'h16 : _T_34503; // @[Mux.scala 31:69:@14088.4]
  assign _T_34505 = valid_43_21 ? 6'h15 : _T_34504; // @[Mux.scala 31:69:@14089.4]
  assign _T_34506 = valid_43_20 ? 6'h14 : _T_34505; // @[Mux.scala 31:69:@14090.4]
  assign _T_34507 = valid_43_19 ? 6'h13 : _T_34506; // @[Mux.scala 31:69:@14091.4]
  assign _T_34508 = valid_43_18 ? 6'h12 : _T_34507; // @[Mux.scala 31:69:@14092.4]
  assign _T_34509 = valid_43_17 ? 6'h11 : _T_34508; // @[Mux.scala 31:69:@14093.4]
  assign _T_34510 = valid_43_16 ? 6'h10 : _T_34509; // @[Mux.scala 31:69:@14094.4]
  assign _T_34511 = valid_43_15 ? 6'hf : _T_34510; // @[Mux.scala 31:69:@14095.4]
  assign _T_34512 = valid_43_14 ? 6'he : _T_34511; // @[Mux.scala 31:69:@14096.4]
  assign _T_34513 = valid_43_13 ? 6'hd : _T_34512; // @[Mux.scala 31:69:@14097.4]
  assign _T_34514 = valid_43_12 ? 6'hc : _T_34513; // @[Mux.scala 31:69:@14098.4]
  assign _T_34515 = valid_43_11 ? 6'hb : _T_34514; // @[Mux.scala 31:69:@14099.4]
  assign _T_34516 = valid_43_10 ? 6'ha : _T_34515; // @[Mux.scala 31:69:@14100.4]
  assign _T_34517 = valid_43_9 ? 6'h9 : _T_34516; // @[Mux.scala 31:69:@14101.4]
  assign _T_34518 = valid_43_8 ? 6'h8 : _T_34517; // @[Mux.scala 31:69:@14102.4]
  assign _T_34519 = valid_43_7 ? 6'h7 : _T_34518; // @[Mux.scala 31:69:@14103.4]
  assign _T_34520 = valid_43_6 ? 6'h6 : _T_34519; // @[Mux.scala 31:69:@14104.4]
  assign _T_34521 = valid_43_5 ? 6'h5 : _T_34520; // @[Mux.scala 31:69:@14105.4]
  assign _T_34522 = valid_43_4 ? 6'h4 : _T_34521; // @[Mux.scala 31:69:@14106.4]
  assign _T_34523 = valid_43_3 ? 6'h3 : _T_34522; // @[Mux.scala 31:69:@14107.4]
  assign _T_34524 = valid_43_2 ? 6'h2 : _T_34523; // @[Mux.scala 31:69:@14108.4]
  assign _T_34525 = valid_43_1 ? 6'h1 : _T_34524; // @[Mux.scala 31:69:@14109.4]
  assign select_43 = valid_43_0 ? 6'h0 : _T_34525; // @[Mux.scala 31:69:@14110.4]
  assign _GEN_2753 = 6'h1 == select_43 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2754 = 6'h2 == select_43 ? io_inData_2 : _GEN_2753; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2755 = 6'h3 == select_43 ? io_inData_3 : _GEN_2754; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2756 = 6'h4 == select_43 ? io_inData_4 : _GEN_2755; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2757 = 6'h5 == select_43 ? io_inData_5 : _GEN_2756; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2758 = 6'h6 == select_43 ? io_inData_6 : _GEN_2757; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2759 = 6'h7 == select_43 ? io_inData_7 : _GEN_2758; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2760 = 6'h8 == select_43 ? io_inData_8 : _GEN_2759; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2761 = 6'h9 == select_43 ? io_inData_9 : _GEN_2760; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2762 = 6'ha == select_43 ? io_inData_10 : _GEN_2761; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2763 = 6'hb == select_43 ? io_inData_11 : _GEN_2762; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2764 = 6'hc == select_43 ? io_inData_12 : _GEN_2763; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2765 = 6'hd == select_43 ? io_inData_13 : _GEN_2764; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2766 = 6'he == select_43 ? io_inData_14 : _GEN_2765; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2767 = 6'hf == select_43 ? io_inData_15 : _GEN_2766; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2768 = 6'h10 == select_43 ? io_inData_16 : _GEN_2767; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2769 = 6'h11 == select_43 ? io_inData_17 : _GEN_2768; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2770 = 6'h12 == select_43 ? io_inData_18 : _GEN_2769; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2771 = 6'h13 == select_43 ? io_inData_19 : _GEN_2770; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2772 = 6'h14 == select_43 ? io_inData_20 : _GEN_2771; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2773 = 6'h15 == select_43 ? io_inData_21 : _GEN_2772; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2774 = 6'h16 == select_43 ? io_inData_22 : _GEN_2773; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2775 = 6'h17 == select_43 ? io_inData_23 : _GEN_2774; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2776 = 6'h18 == select_43 ? io_inData_24 : _GEN_2775; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2777 = 6'h19 == select_43 ? io_inData_25 : _GEN_2776; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2778 = 6'h1a == select_43 ? io_inData_26 : _GEN_2777; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2779 = 6'h1b == select_43 ? io_inData_27 : _GEN_2778; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2780 = 6'h1c == select_43 ? io_inData_28 : _GEN_2779; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2781 = 6'h1d == select_43 ? io_inData_29 : _GEN_2780; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2782 = 6'h1e == select_43 ? io_inData_30 : _GEN_2781; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2783 = 6'h1f == select_43 ? io_inData_31 : _GEN_2782; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2784 = 6'h20 == select_43 ? io_inData_32 : _GEN_2783; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2785 = 6'h21 == select_43 ? io_inData_33 : _GEN_2784; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2786 = 6'h22 == select_43 ? io_inData_34 : _GEN_2785; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2787 = 6'h23 == select_43 ? io_inData_35 : _GEN_2786; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2788 = 6'h24 == select_43 ? io_inData_36 : _GEN_2787; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2789 = 6'h25 == select_43 ? io_inData_37 : _GEN_2788; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2790 = 6'h26 == select_43 ? io_inData_38 : _GEN_2789; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2791 = 6'h27 == select_43 ? io_inData_39 : _GEN_2790; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2792 = 6'h28 == select_43 ? io_inData_40 : _GEN_2791; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2793 = 6'h29 == select_43 ? io_inData_41 : _GEN_2792; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2794 = 6'h2a == select_43 ? io_inData_42 : _GEN_2793; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2795 = 6'h2b == select_43 ? io_inData_43 : _GEN_2794; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2796 = 6'h2c == select_43 ? io_inData_44 : _GEN_2795; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2797 = 6'h2d == select_43 ? io_inData_45 : _GEN_2796; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2798 = 6'h2e == select_43 ? io_inData_46 : _GEN_2797; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2799 = 6'h2f == select_43 ? io_inData_47 : _GEN_2798; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2800 = 6'h30 == select_43 ? io_inData_48 : _GEN_2799; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2801 = 6'h31 == select_43 ? io_inData_49 : _GEN_2800; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2802 = 6'h32 == select_43 ? io_inData_50 : _GEN_2801; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2803 = 6'h33 == select_43 ? io_inData_51 : _GEN_2802; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2804 = 6'h34 == select_43 ? io_inData_52 : _GEN_2803; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2805 = 6'h35 == select_43 ? io_inData_53 : _GEN_2804; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2806 = 6'h36 == select_43 ? io_inData_54 : _GEN_2805; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2807 = 6'h37 == select_43 ? io_inData_55 : _GEN_2806; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2808 = 6'h38 == select_43 ? io_inData_56 : _GEN_2807; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2809 = 6'h39 == select_43 ? io_inData_57 : _GEN_2808; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2810 = 6'h3a == select_43 ? io_inData_58 : _GEN_2809; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2811 = 6'h3b == select_43 ? io_inData_59 : _GEN_2810; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2812 = 6'h3c == select_43 ? io_inData_60 : _GEN_2811; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2813 = 6'h3d == select_43 ? io_inData_61 : _GEN_2812; // @[Switch.scala 33:19:@14112.4]
  assign _GEN_2814 = 6'h3e == select_43 ? io_inData_62 : _GEN_2813; // @[Switch.scala 33:19:@14112.4]
  assign _T_34534 = {valid_43_7,valid_43_6,valid_43_5,valid_43_4,valid_43_3,valid_43_2,valid_43_1,valid_43_0}; // @[Switch.scala 34:32:@14119.4]
  assign _T_34542 = {valid_43_15,valid_43_14,valid_43_13,valid_43_12,valid_43_11,valid_43_10,valid_43_9,valid_43_8,_T_34534}; // @[Switch.scala 34:32:@14127.4]
  assign _T_34549 = {valid_43_23,valid_43_22,valid_43_21,valid_43_20,valid_43_19,valid_43_18,valid_43_17,valid_43_16}; // @[Switch.scala 34:32:@14134.4]
  assign _T_34558 = {valid_43_31,valid_43_30,valid_43_29,valid_43_28,valid_43_27,valid_43_26,valid_43_25,valid_43_24,_T_34549,_T_34542}; // @[Switch.scala 34:32:@14143.4]
  assign _T_34565 = {valid_43_39,valid_43_38,valid_43_37,valid_43_36,valid_43_35,valid_43_34,valid_43_33,valid_43_32}; // @[Switch.scala 34:32:@14150.4]
  assign _T_34573 = {valid_43_47,valid_43_46,valid_43_45,valid_43_44,valid_43_43,valid_43_42,valid_43_41,valid_43_40,_T_34565}; // @[Switch.scala 34:32:@14158.4]
  assign _T_34580 = {valid_43_55,valid_43_54,valid_43_53,valid_43_52,valid_43_51,valid_43_50,valid_43_49,valid_43_48}; // @[Switch.scala 34:32:@14165.4]
  assign _T_34589 = {valid_43_63,valid_43_62,valid_43_61,valid_43_60,valid_43_59,valid_43_58,valid_43_57,valid_43_56,_T_34580,_T_34573}; // @[Switch.scala 34:32:@14174.4]
  assign _T_34590 = {_T_34589,_T_34558}; // @[Switch.scala 34:32:@14175.4]
  assign _T_34594 = io_inAddr_0 == 6'h2c; // @[Switch.scala 30:53:@14178.4]
  assign valid_44_0 = io_inValid_0 & _T_34594; // @[Switch.scala 30:36:@14179.4]
  assign _T_34597 = io_inAddr_1 == 6'h2c; // @[Switch.scala 30:53:@14181.4]
  assign valid_44_1 = io_inValid_1 & _T_34597; // @[Switch.scala 30:36:@14182.4]
  assign _T_34600 = io_inAddr_2 == 6'h2c; // @[Switch.scala 30:53:@14184.4]
  assign valid_44_2 = io_inValid_2 & _T_34600; // @[Switch.scala 30:36:@14185.4]
  assign _T_34603 = io_inAddr_3 == 6'h2c; // @[Switch.scala 30:53:@14187.4]
  assign valid_44_3 = io_inValid_3 & _T_34603; // @[Switch.scala 30:36:@14188.4]
  assign _T_34606 = io_inAddr_4 == 6'h2c; // @[Switch.scala 30:53:@14190.4]
  assign valid_44_4 = io_inValid_4 & _T_34606; // @[Switch.scala 30:36:@14191.4]
  assign _T_34609 = io_inAddr_5 == 6'h2c; // @[Switch.scala 30:53:@14193.4]
  assign valid_44_5 = io_inValid_5 & _T_34609; // @[Switch.scala 30:36:@14194.4]
  assign _T_34612 = io_inAddr_6 == 6'h2c; // @[Switch.scala 30:53:@14196.4]
  assign valid_44_6 = io_inValid_6 & _T_34612; // @[Switch.scala 30:36:@14197.4]
  assign _T_34615 = io_inAddr_7 == 6'h2c; // @[Switch.scala 30:53:@14199.4]
  assign valid_44_7 = io_inValid_7 & _T_34615; // @[Switch.scala 30:36:@14200.4]
  assign _T_34618 = io_inAddr_8 == 6'h2c; // @[Switch.scala 30:53:@14202.4]
  assign valid_44_8 = io_inValid_8 & _T_34618; // @[Switch.scala 30:36:@14203.4]
  assign _T_34621 = io_inAddr_9 == 6'h2c; // @[Switch.scala 30:53:@14205.4]
  assign valid_44_9 = io_inValid_9 & _T_34621; // @[Switch.scala 30:36:@14206.4]
  assign _T_34624 = io_inAddr_10 == 6'h2c; // @[Switch.scala 30:53:@14208.4]
  assign valid_44_10 = io_inValid_10 & _T_34624; // @[Switch.scala 30:36:@14209.4]
  assign _T_34627 = io_inAddr_11 == 6'h2c; // @[Switch.scala 30:53:@14211.4]
  assign valid_44_11 = io_inValid_11 & _T_34627; // @[Switch.scala 30:36:@14212.4]
  assign _T_34630 = io_inAddr_12 == 6'h2c; // @[Switch.scala 30:53:@14214.4]
  assign valid_44_12 = io_inValid_12 & _T_34630; // @[Switch.scala 30:36:@14215.4]
  assign _T_34633 = io_inAddr_13 == 6'h2c; // @[Switch.scala 30:53:@14217.4]
  assign valid_44_13 = io_inValid_13 & _T_34633; // @[Switch.scala 30:36:@14218.4]
  assign _T_34636 = io_inAddr_14 == 6'h2c; // @[Switch.scala 30:53:@14220.4]
  assign valid_44_14 = io_inValid_14 & _T_34636; // @[Switch.scala 30:36:@14221.4]
  assign _T_34639 = io_inAddr_15 == 6'h2c; // @[Switch.scala 30:53:@14223.4]
  assign valid_44_15 = io_inValid_15 & _T_34639; // @[Switch.scala 30:36:@14224.4]
  assign _T_34642 = io_inAddr_16 == 6'h2c; // @[Switch.scala 30:53:@14226.4]
  assign valid_44_16 = io_inValid_16 & _T_34642; // @[Switch.scala 30:36:@14227.4]
  assign _T_34645 = io_inAddr_17 == 6'h2c; // @[Switch.scala 30:53:@14229.4]
  assign valid_44_17 = io_inValid_17 & _T_34645; // @[Switch.scala 30:36:@14230.4]
  assign _T_34648 = io_inAddr_18 == 6'h2c; // @[Switch.scala 30:53:@14232.4]
  assign valid_44_18 = io_inValid_18 & _T_34648; // @[Switch.scala 30:36:@14233.4]
  assign _T_34651 = io_inAddr_19 == 6'h2c; // @[Switch.scala 30:53:@14235.4]
  assign valid_44_19 = io_inValid_19 & _T_34651; // @[Switch.scala 30:36:@14236.4]
  assign _T_34654 = io_inAddr_20 == 6'h2c; // @[Switch.scala 30:53:@14238.4]
  assign valid_44_20 = io_inValid_20 & _T_34654; // @[Switch.scala 30:36:@14239.4]
  assign _T_34657 = io_inAddr_21 == 6'h2c; // @[Switch.scala 30:53:@14241.4]
  assign valid_44_21 = io_inValid_21 & _T_34657; // @[Switch.scala 30:36:@14242.4]
  assign _T_34660 = io_inAddr_22 == 6'h2c; // @[Switch.scala 30:53:@14244.4]
  assign valid_44_22 = io_inValid_22 & _T_34660; // @[Switch.scala 30:36:@14245.4]
  assign _T_34663 = io_inAddr_23 == 6'h2c; // @[Switch.scala 30:53:@14247.4]
  assign valid_44_23 = io_inValid_23 & _T_34663; // @[Switch.scala 30:36:@14248.4]
  assign _T_34666 = io_inAddr_24 == 6'h2c; // @[Switch.scala 30:53:@14250.4]
  assign valid_44_24 = io_inValid_24 & _T_34666; // @[Switch.scala 30:36:@14251.4]
  assign _T_34669 = io_inAddr_25 == 6'h2c; // @[Switch.scala 30:53:@14253.4]
  assign valid_44_25 = io_inValid_25 & _T_34669; // @[Switch.scala 30:36:@14254.4]
  assign _T_34672 = io_inAddr_26 == 6'h2c; // @[Switch.scala 30:53:@14256.4]
  assign valid_44_26 = io_inValid_26 & _T_34672; // @[Switch.scala 30:36:@14257.4]
  assign _T_34675 = io_inAddr_27 == 6'h2c; // @[Switch.scala 30:53:@14259.4]
  assign valid_44_27 = io_inValid_27 & _T_34675; // @[Switch.scala 30:36:@14260.4]
  assign _T_34678 = io_inAddr_28 == 6'h2c; // @[Switch.scala 30:53:@14262.4]
  assign valid_44_28 = io_inValid_28 & _T_34678; // @[Switch.scala 30:36:@14263.4]
  assign _T_34681 = io_inAddr_29 == 6'h2c; // @[Switch.scala 30:53:@14265.4]
  assign valid_44_29 = io_inValid_29 & _T_34681; // @[Switch.scala 30:36:@14266.4]
  assign _T_34684 = io_inAddr_30 == 6'h2c; // @[Switch.scala 30:53:@14268.4]
  assign valid_44_30 = io_inValid_30 & _T_34684; // @[Switch.scala 30:36:@14269.4]
  assign _T_34687 = io_inAddr_31 == 6'h2c; // @[Switch.scala 30:53:@14271.4]
  assign valid_44_31 = io_inValid_31 & _T_34687; // @[Switch.scala 30:36:@14272.4]
  assign _T_34690 = io_inAddr_32 == 6'h2c; // @[Switch.scala 30:53:@14274.4]
  assign valid_44_32 = io_inValid_32 & _T_34690; // @[Switch.scala 30:36:@14275.4]
  assign _T_34693 = io_inAddr_33 == 6'h2c; // @[Switch.scala 30:53:@14277.4]
  assign valid_44_33 = io_inValid_33 & _T_34693; // @[Switch.scala 30:36:@14278.4]
  assign _T_34696 = io_inAddr_34 == 6'h2c; // @[Switch.scala 30:53:@14280.4]
  assign valid_44_34 = io_inValid_34 & _T_34696; // @[Switch.scala 30:36:@14281.4]
  assign _T_34699 = io_inAddr_35 == 6'h2c; // @[Switch.scala 30:53:@14283.4]
  assign valid_44_35 = io_inValid_35 & _T_34699; // @[Switch.scala 30:36:@14284.4]
  assign _T_34702 = io_inAddr_36 == 6'h2c; // @[Switch.scala 30:53:@14286.4]
  assign valid_44_36 = io_inValid_36 & _T_34702; // @[Switch.scala 30:36:@14287.4]
  assign _T_34705 = io_inAddr_37 == 6'h2c; // @[Switch.scala 30:53:@14289.4]
  assign valid_44_37 = io_inValid_37 & _T_34705; // @[Switch.scala 30:36:@14290.4]
  assign _T_34708 = io_inAddr_38 == 6'h2c; // @[Switch.scala 30:53:@14292.4]
  assign valid_44_38 = io_inValid_38 & _T_34708; // @[Switch.scala 30:36:@14293.4]
  assign _T_34711 = io_inAddr_39 == 6'h2c; // @[Switch.scala 30:53:@14295.4]
  assign valid_44_39 = io_inValid_39 & _T_34711; // @[Switch.scala 30:36:@14296.4]
  assign _T_34714 = io_inAddr_40 == 6'h2c; // @[Switch.scala 30:53:@14298.4]
  assign valid_44_40 = io_inValid_40 & _T_34714; // @[Switch.scala 30:36:@14299.4]
  assign _T_34717 = io_inAddr_41 == 6'h2c; // @[Switch.scala 30:53:@14301.4]
  assign valid_44_41 = io_inValid_41 & _T_34717; // @[Switch.scala 30:36:@14302.4]
  assign _T_34720 = io_inAddr_42 == 6'h2c; // @[Switch.scala 30:53:@14304.4]
  assign valid_44_42 = io_inValid_42 & _T_34720; // @[Switch.scala 30:36:@14305.4]
  assign _T_34723 = io_inAddr_43 == 6'h2c; // @[Switch.scala 30:53:@14307.4]
  assign valid_44_43 = io_inValid_43 & _T_34723; // @[Switch.scala 30:36:@14308.4]
  assign _T_34726 = io_inAddr_44 == 6'h2c; // @[Switch.scala 30:53:@14310.4]
  assign valid_44_44 = io_inValid_44 & _T_34726; // @[Switch.scala 30:36:@14311.4]
  assign _T_34729 = io_inAddr_45 == 6'h2c; // @[Switch.scala 30:53:@14313.4]
  assign valid_44_45 = io_inValid_45 & _T_34729; // @[Switch.scala 30:36:@14314.4]
  assign _T_34732 = io_inAddr_46 == 6'h2c; // @[Switch.scala 30:53:@14316.4]
  assign valid_44_46 = io_inValid_46 & _T_34732; // @[Switch.scala 30:36:@14317.4]
  assign _T_34735 = io_inAddr_47 == 6'h2c; // @[Switch.scala 30:53:@14319.4]
  assign valid_44_47 = io_inValid_47 & _T_34735; // @[Switch.scala 30:36:@14320.4]
  assign _T_34738 = io_inAddr_48 == 6'h2c; // @[Switch.scala 30:53:@14322.4]
  assign valid_44_48 = io_inValid_48 & _T_34738; // @[Switch.scala 30:36:@14323.4]
  assign _T_34741 = io_inAddr_49 == 6'h2c; // @[Switch.scala 30:53:@14325.4]
  assign valid_44_49 = io_inValid_49 & _T_34741; // @[Switch.scala 30:36:@14326.4]
  assign _T_34744 = io_inAddr_50 == 6'h2c; // @[Switch.scala 30:53:@14328.4]
  assign valid_44_50 = io_inValid_50 & _T_34744; // @[Switch.scala 30:36:@14329.4]
  assign _T_34747 = io_inAddr_51 == 6'h2c; // @[Switch.scala 30:53:@14331.4]
  assign valid_44_51 = io_inValid_51 & _T_34747; // @[Switch.scala 30:36:@14332.4]
  assign _T_34750 = io_inAddr_52 == 6'h2c; // @[Switch.scala 30:53:@14334.4]
  assign valid_44_52 = io_inValid_52 & _T_34750; // @[Switch.scala 30:36:@14335.4]
  assign _T_34753 = io_inAddr_53 == 6'h2c; // @[Switch.scala 30:53:@14337.4]
  assign valid_44_53 = io_inValid_53 & _T_34753; // @[Switch.scala 30:36:@14338.4]
  assign _T_34756 = io_inAddr_54 == 6'h2c; // @[Switch.scala 30:53:@14340.4]
  assign valid_44_54 = io_inValid_54 & _T_34756; // @[Switch.scala 30:36:@14341.4]
  assign _T_34759 = io_inAddr_55 == 6'h2c; // @[Switch.scala 30:53:@14343.4]
  assign valid_44_55 = io_inValid_55 & _T_34759; // @[Switch.scala 30:36:@14344.4]
  assign _T_34762 = io_inAddr_56 == 6'h2c; // @[Switch.scala 30:53:@14346.4]
  assign valid_44_56 = io_inValid_56 & _T_34762; // @[Switch.scala 30:36:@14347.4]
  assign _T_34765 = io_inAddr_57 == 6'h2c; // @[Switch.scala 30:53:@14349.4]
  assign valid_44_57 = io_inValid_57 & _T_34765; // @[Switch.scala 30:36:@14350.4]
  assign _T_34768 = io_inAddr_58 == 6'h2c; // @[Switch.scala 30:53:@14352.4]
  assign valid_44_58 = io_inValid_58 & _T_34768; // @[Switch.scala 30:36:@14353.4]
  assign _T_34771 = io_inAddr_59 == 6'h2c; // @[Switch.scala 30:53:@14355.4]
  assign valid_44_59 = io_inValid_59 & _T_34771; // @[Switch.scala 30:36:@14356.4]
  assign _T_34774 = io_inAddr_60 == 6'h2c; // @[Switch.scala 30:53:@14358.4]
  assign valid_44_60 = io_inValid_60 & _T_34774; // @[Switch.scala 30:36:@14359.4]
  assign _T_34777 = io_inAddr_61 == 6'h2c; // @[Switch.scala 30:53:@14361.4]
  assign valid_44_61 = io_inValid_61 & _T_34777; // @[Switch.scala 30:36:@14362.4]
  assign _T_34780 = io_inAddr_62 == 6'h2c; // @[Switch.scala 30:53:@14364.4]
  assign valid_44_62 = io_inValid_62 & _T_34780; // @[Switch.scala 30:36:@14365.4]
  assign _T_34783 = io_inAddr_63 == 6'h2c; // @[Switch.scala 30:53:@14367.4]
  assign valid_44_63 = io_inValid_63 & _T_34783; // @[Switch.scala 30:36:@14368.4]
  assign _T_34849 = valid_44_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@14370.4]
  assign _T_34850 = valid_44_61 ? 6'h3d : _T_34849; // @[Mux.scala 31:69:@14371.4]
  assign _T_34851 = valid_44_60 ? 6'h3c : _T_34850; // @[Mux.scala 31:69:@14372.4]
  assign _T_34852 = valid_44_59 ? 6'h3b : _T_34851; // @[Mux.scala 31:69:@14373.4]
  assign _T_34853 = valid_44_58 ? 6'h3a : _T_34852; // @[Mux.scala 31:69:@14374.4]
  assign _T_34854 = valid_44_57 ? 6'h39 : _T_34853; // @[Mux.scala 31:69:@14375.4]
  assign _T_34855 = valid_44_56 ? 6'h38 : _T_34854; // @[Mux.scala 31:69:@14376.4]
  assign _T_34856 = valid_44_55 ? 6'h37 : _T_34855; // @[Mux.scala 31:69:@14377.4]
  assign _T_34857 = valid_44_54 ? 6'h36 : _T_34856; // @[Mux.scala 31:69:@14378.4]
  assign _T_34858 = valid_44_53 ? 6'h35 : _T_34857; // @[Mux.scala 31:69:@14379.4]
  assign _T_34859 = valid_44_52 ? 6'h34 : _T_34858; // @[Mux.scala 31:69:@14380.4]
  assign _T_34860 = valid_44_51 ? 6'h33 : _T_34859; // @[Mux.scala 31:69:@14381.4]
  assign _T_34861 = valid_44_50 ? 6'h32 : _T_34860; // @[Mux.scala 31:69:@14382.4]
  assign _T_34862 = valid_44_49 ? 6'h31 : _T_34861; // @[Mux.scala 31:69:@14383.4]
  assign _T_34863 = valid_44_48 ? 6'h30 : _T_34862; // @[Mux.scala 31:69:@14384.4]
  assign _T_34864 = valid_44_47 ? 6'h2f : _T_34863; // @[Mux.scala 31:69:@14385.4]
  assign _T_34865 = valid_44_46 ? 6'h2e : _T_34864; // @[Mux.scala 31:69:@14386.4]
  assign _T_34866 = valid_44_45 ? 6'h2d : _T_34865; // @[Mux.scala 31:69:@14387.4]
  assign _T_34867 = valid_44_44 ? 6'h2c : _T_34866; // @[Mux.scala 31:69:@14388.4]
  assign _T_34868 = valid_44_43 ? 6'h2b : _T_34867; // @[Mux.scala 31:69:@14389.4]
  assign _T_34869 = valid_44_42 ? 6'h2a : _T_34868; // @[Mux.scala 31:69:@14390.4]
  assign _T_34870 = valid_44_41 ? 6'h29 : _T_34869; // @[Mux.scala 31:69:@14391.4]
  assign _T_34871 = valid_44_40 ? 6'h28 : _T_34870; // @[Mux.scala 31:69:@14392.4]
  assign _T_34872 = valid_44_39 ? 6'h27 : _T_34871; // @[Mux.scala 31:69:@14393.4]
  assign _T_34873 = valid_44_38 ? 6'h26 : _T_34872; // @[Mux.scala 31:69:@14394.4]
  assign _T_34874 = valid_44_37 ? 6'h25 : _T_34873; // @[Mux.scala 31:69:@14395.4]
  assign _T_34875 = valid_44_36 ? 6'h24 : _T_34874; // @[Mux.scala 31:69:@14396.4]
  assign _T_34876 = valid_44_35 ? 6'h23 : _T_34875; // @[Mux.scala 31:69:@14397.4]
  assign _T_34877 = valid_44_34 ? 6'h22 : _T_34876; // @[Mux.scala 31:69:@14398.4]
  assign _T_34878 = valid_44_33 ? 6'h21 : _T_34877; // @[Mux.scala 31:69:@14399.4]
  assign _T_34879 = valid_44_32 ? 6'h20 : _T_34878; // @[Mux.scala 31:69:@14400.4]
  assign _T_34880 = valid_44_31 ? 6'h1f : _T_34879; // @[Mux.scala 31:69:@14401.4]
  assign _T_34881 = valid_44_30 ? 6'h1e : _T_34880; // @[Mux.scala 31:69:@14402.4]
  assign _T_34882 = valid_44_29 ? 6'h1d : _T_34881; // @[Mux.scala 31:69:@14403.4]
  assign _T_34883 = valid_44_28 ? 6'h1c : _T_34882; // @[Mux.scala 31:69:@14404.4]
  assign _T_34884 = valid_44_27 ? 6'h1b : _T_34883; // @[Mux.scala 31:69:@14405.4]
  assign _T_34885 = valid_44_26 ? 6'h1a : _T_34884; // @[Mux.scala 31:69:@14406.4]
  assign _T_34886 = valid_44_25 ? 6'h19 : _T_34885; // @[Mux.scala 31:69:@14407.4]
  assign _T_34887 = valid_44_24 ? 6'h18 : _T_34886; // @[Mux.scala 31:69:@14408.4]
  assign _T_34888 = valid_44_23 ? 6'h17 : _T_34887; // @[Mux.scala 31:69:@14409.4]
  assign _T_34889 = valid_44_22 ? 6'h16 : _T_34888; // @[Mux.scala 31:69:@14410.4]
  assign _T_34890 = valid_44_21 ? 6'h15 : _T_34889; // @[Mux.scala 31:69:@14411.4]
  assign _T_34891 = valid_44_20 ? 6'h14 : _T_34890; // @[Mux.scala 31:69:@14412.4]
  assign _T_34892 = valid_44_19 ? 6'h13 : _T_34891; // @[Mux.scala 31:69:@14413.4]
  assign _T_34893 = valid_44_18 ? 6'h12 : _T_34892; // @[Mux.scala 31:69:@14414.4]
  assign _T_34894 = valid_44_17 ? 6'h11 : _T_34893; // @[Mux.scala 31:69:@14415.4]
  assign _T_34895 = valid_44_16 ? 6'h10 : _T_34894; // @[Mux.scala 31:69:@14416.4]
  assign _T_34896 = valid_44_15 ? 6'hf : _T_34895; // @[Mux.scala 31:69:@14417.4]
  assign _T_34897 = valid_44_14 ? 6'he : _T_34896; // @[Mux.scala 31:69:@14418.4]
  assign _T_34898 = valid_44_13 ? 6'hd : _T_34897; // @[Mux.scala 31:69:@14419.4]
  assign _T_34899 = valid_44_12 ? 6'hc : _T_34898; // @[Mux.scala 31:69:@14420.4]
  assign _T_34900 = valid_44_11 ? 6'hb : _T_34899; // @[Mux.scala 31:69:@14421.4]
  assign _T_34901 = valid_44_10 ? 6'ha : _T_34900; // @[Mux.scala 31:69:@14422.4]
  assign _T_34902 = valid_44_9 ? 6'h9 : _T_34901; // @[Mux.scala 31:69:@14423.4]
  assign _T_34903 = valid_44_8 ? 6'h8 : _T_34902; // @[Mux.scala 31:69:@14424.4]
  assign _T_34904 = valid_44_7 ? 6'h7 : _T_34903; // @[Mux.scala 31:69:@14425.4]
  assign _T_34905 = valid_44_6 ? 6'h6 : _T_34904; // @[Mux.scala 31:69:@14426.4]
  assign _T_34906 = valid_44_5 ? 6'h5 : _T_34905; // @[Mux.scala 31:69:@14427.4]
  assign _T_34907 = valid_44_4 ? 6'h4 : _T_34906; // @[Mux.scala 31:69:@14428.4]
  assign _T_34908 = valid_44_3 ? 6'h3 : _T_34907; // @[Mux.scala 31:69:@14429.4]
  assign _T_34909 = valid_44_2 ? 6'h2 : _T_34908; // @[Mux.scala 31:69:@14430.4]
  assign _T_34910 = valid_44_1 ? 6'h1 : _T_34909; // @[Mux.scala 31:69:@14431.4]
  assign select_44 = valid_44_0 ? 6'h0 : _T_34910; // @[Mux.scala 31:69:@14432.4]
  assign _GEN_2817 = 6'h1 == select_44 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2818 = 6'h2 == select_44 ? io_inData_2 : _GEN_2817; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2819 = 6'h3 == select_44 ? io_inData_3 : _GEN_2818; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2820 = 6'h4 == select_44 ? io_inData_4 : _GEN_2819; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2821 = 6'h5 == select_44 ? io_inData_5 : _GEN_2820; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2822 = 6'h6 == select_44 ? io_inData_6 : _GEN_2821; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2823 = 6'h7 == select_44 ? io_inData_7 : _GEN_2822; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2824 = 6'h8 == select_44 ? io_inData_8 : _GEN_2823; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2825 = 6'h9 == select_44 ? io_inData_9 : _GEN_2824; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2826 = 6'ha == select_44 ? io_inData_10 : _GEN_2825; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2827 = 6'hb == select_44 ? io_inData_11 : _GEN_2826; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2828 = 6'hc == select_44 ? io_inData_12 : _GEN_2827; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2829 = 6'hd == select_44 ? io_inData_13 : _GEN_2828; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2830 = 6'he == select_44 ? io_inData_14 : _GEN_2829; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2831 = 6'hf == select_44 ? io_inData_15 : _GEN_2830; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2832 = 6'h10 == select_44 ? io_inData_16 : _GEN_2831; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2833 = 6'h11 == select_44 ? io_inData_17 : _GEN_2832; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2834 = 6'h12 == select_44 ? io_inData_18 : _GEN_2833; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2835 = 6'h13 == select_44 ? io_inData_19 : _GEN_2834; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2836 = 6'h14 == select_44 ? io_inData_20 : _GEN_2835; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2837 = 6'h15 == select_44 ? io_inData_21 : _GEN_2836; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2838 = 6'h16 == select_44 ? io_inData_22 : _GEN_2837; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2839 = 6'h17 == select_44 ? io_inData_23 : _GEN_2838; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2840 = 6'h18 == select_44 ? io_inData_24 : _GEN_2839; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2841 = 6'h19 == select_44 ? io_inData_25 : _GEN_2840; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2842 = 6'h1a == select_44 ? io_inData_26 : _GEN_2841; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2843 = 6'h1b == select_44 ? io_inData_27 : _GEN_2842; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2844 = 6'h1c == select_44 ? io_inData_28 : _GEN_2843; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2845 = 6'h1d == select_44 ? io_inData_29 : _GEN_2844; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2846 = 6'h1e == select_44 ? io_inData_30 : _GEN_2845; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2847 = 6'h1f == select_44 ? io_inData_31 : _GEN_2846; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2848 = 6'h20 == select_44 ? io_inData_32 : _GEN_2847; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2849 = 6'h21 == select_44 ? io_inData_33 : _GEN_2848; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2850 = 6'h22 == select_44 ? io_inData_34 : _GEN_2849; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2851 = 6'h23 == select_44 ? io_inData_35 : _GEN_2850; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2852 = 6'h24 == select_44 ? io_inData_36 : _GEN_2851; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2853 = 6'h25 == select_44 ? io_inData_37 : _GEN_2852; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2854 = 6'h26 == select_44 ? io_inData_38 : _GEN_2853; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2855 = 6'h27 == select_44 ? io_inData_39 : _GEN_2854; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2856 = 6'h28 == select_44 ? io_inData_40 : _GEN_2855; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2857 = 6'h29 == select_44 ? io_inData_41 : _GEN_2856; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2858 = 6'h2a == select_44 ? io_inData_42 : _GEN_2857; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2859 = 6'h2b == select_44 ? io_inData_43 : _GEN_2858; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2860 = 6'h2c == select_44 ? io_inData_44 : _GEN_2859; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2861 = 6'h2d == select_44 ? io_inData_45 : _GEN_2860; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2862 = 6'h2e == select_44 ? io_inData_46 : _GEN_2861; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2863 = 6'h2f == select_44 ? io_inData_47 : _GEN_2862; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2864 = 6'h30 == select_44 ? io_inData_48 : _GEN_2863; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2865 = 6'h31 == select_44 ? io_inData_49 : _GEN_2864; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2866 = 6'h32 == select_44 ? io_inData_50 : _GEN_2865; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2867 = 6'h33 == select_44 ? io_inData_51 : _GEN_2866; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2868 = 6'h34 == select_44 ? io_inData_52 : _GEN_2867; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2869 = 6'h35 == select_44 ? io_inData_53 : _GEN_2868; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2870 = 6'h36 == select_44 ? io_inData_54 : _GEN_2869; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2871 = 6'h37 == select_44 ? io_inData_55 : _GEN_2870; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2872 = 6'h38 == select_44 ? io_inData_56 : _GEN_2871; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2873 = 6'h39 == select_44 ? io_inData_57 : _GEN_2872; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2874 = 6'h3a == select_44 ? io_inData_58 : _GEN_2873; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2875 = 6'h3b == select_44 ? io_inData_59 : _GEN_2874; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2876 = 6'h3c == select_44 ? io_inData_60 : _GEN_2875; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2877 = 6'h3d == select_44 ? io_inData_61 : _GEN_2876; // @[Switch.scala 33:19:@14434.4]
  assign _GEN_2878 = 6'h3e == select_44 ? io_inData_62 : _GEN_2877; // @[Switch.scala 33:19:@14434.4]
  assign _T_34919 = {valid_44_7,valid_44_6,valid_44_5,valid_44_4,valid_44_3,valid_44_2,valid_44_1,valid_44_0}; // @[Switch.scala 34:32:@14441.4]
  assign _T_34927 = {valid_44_15,valid_44_14,valid_44_13,valid_44_12,valid_44_11,valid_44_10,valid_44_9,valid_44_8,_T_34919}; // @[Switch.scala 34:32:@14449.4]
  assign _T_34934 = {valid_44_23,valid_44_22,valid_44_21,valid_44_20,valid_44_19,valid_44_18,valid_44_17,valid_44_16}; // @[Switch.scala 34:32:@14456.4]
  assign _T_34943 = {valid_44_31,valid_44_30,valid_44_29,valid_44_28,valid_44_27,valid_44_26,valid_44_25,valid_44_24,_T_34934,_T_34927}; // @[Switch.scala 34:32:@14465.4]
  assign _T_34950 = {valid_44_39,valid_44_38,valid_44_37,valid_44_36,valid_44_35,valid_44_34,valid_44_33,valid_44_32}; // @[Switch.scala 34:32:@14472.4]
  assign _T_34958 = {valid_44_47,valid_44_46,valid_44_45,valid_44_44,valid_44_43,valid_44_42,valid_44_41,valid_44_40,_T_34950}; // @[Switch.scala 34:32:@14480.4]
  assign _T_34965 = {valid_44_55,valid_44_54,valid_44_53,valid_44_52,valid_44_51,valid_44_50,valid_44_49,valid_44_48}; // @[Switch.scala 34:32:@14487.4]
  assign _T_34974 = {valid_44_63,valid_44_62,valid_44_61,valid_44_60,valid_44_59,valid_44_58,valid_44_57,valid_44_56,_T_34965,_T_34958}; // @[Switch.scala 34:32:@14496.4]
  assign _T_34975 = {_T_34974,_T_34943}; // @[Switch.scala 34:32:@14497.4]
  assign _T_34979 = io_inAddr_0 == 6'h2d; // @[Switch.scala 30:53:@14500.4]
  assign valid_45_0 = io_inValid_0 & _T_34979; // @[Switch.scala 30:36:@14501.4]
  assign _T_34982 = io_inAddr_1 == 6'h2d; // @[Switch.scala 30:53:@14503.4]
  assign valid_45_1 = io_inValid_1 & _T_34982; // @[Switch.scala 30:36:@14504.4]
  assign _T_34985 = io_inAddr_2 == 6'h2d; // @[Switch.scala 30:53:@14506.4]
  assign valid_45_2 = io_inValid_2 & _T_34985; // @[Switch.scala 30:36:@14507.4]
  assign _T_34988 = io_inAddr_3 == 6'h2d; // @[Switch.scala 30:53:@14509.4]
  assign valid_45_3 = io_inValid_3 & _T_34988; // @[Switch.scala 30:36:@14510.4]
  assign _T_34991 = io_inAddr_4 == 6'h2d; // @[Switch.scala 30:53:@14512.4]
  assign valid_45_4 = io_inValid_4 & _T_34991; // @[Switch.scala 30:36:@14513.4]
  assign _T_34994 = io_inAddr_5 == 6'h2d; // @[Switch.scala 30:53:@14515.4]
  assign valid_45_5 = io_inValid_5 & _T_34994; // @[Switch.scala 30:36:@14516.4]
  assign _T_34997 = io_inAddr_6 == 6'h2d; // @[Switch.scala 30:53:@14518.4]
  assign valid_45_6 = io_inValid_6 & _T_34997; // @[Switch.scala 30:36:@14519.4]
  assign _T_35000 = io_inAddr_7 == 6'h2d; // @[Switch.scala 30:53:@14521.4]
  assign valid_45_7 = io_inValid_7 & _T_35000; // @[Switch.scala 30:36:@14522.4]
  assign _T_35003 = io_inAddr_8 == 6'h2d; // @[Switch.scala 30:53:@14524.4]
  assign valid_45_8 = io_inValid_8 & _T_35003; // @[Switch.scala 30:36:@14525.4]
  assign _T_35006 = io_inAddr_9 == 6'h2d; // @[Switch.scala 30:53:@14527.4]
  assign valid_45_9 = io_inValid_9 & _T_35006; // @[Switch.scala 30:36:@14528.4]
  assign _T_35009 = io_inAddr_10 == 6'h2d; // @[Switch.scala 30:53:@14530.4]
  assign valid_45_10 = io_inValid_10 & _T_35009; // @[Switch.scala 30:36:@14531.4]
  assign _T_35012 = io_inAddr_11 == 6'h2d; // @[Switch.scala 30:53:@14533.4]
  assign valid_45_11 = io_inValid_11 & _T_35012; // @[Switch.scala 30:36:@14534.4]
  assign _T_35015 = io_inAddr_12 == 6'h2d; // @[Switch.scala 30:53:@14536.4]
  assign valid_45_12 = io_inValid_12 & _T_35015; // @[Switch.scala 30:36:@14537.4]
  assign _T_35018 = io_inAddr_13 == 6'h2d; // @[Switch.scala 30:53:@14539.4]
  assign valid_45_13 = io_inValid_13 & _T_35018; // @[Switch.scala 30:36:@14540.4]
  assign _T_35021 = io_inAddr_14 == 6'h2d; // @[Switch.scala 30:53:@14542.4]
  assign valid_45_14 = io_inValid_14 & _T_35021; // @[Switch.scala 30:36:@14543.4]
  assign _T_35024 = io_inAddr_15 == 6'h2d; // @[Switch.scala 30:53:@14545.4]
  assign valid_45_15 = io_inValid_15 & _T_35024; // @[Switch.scala 30:36:@14546.4]
  assign _T_35027 = io_inAddr_16 == 6'h2d; // @[Switch.scala 30:53:@14548.4]
  assign valid_45_16 = io_inValid_16 & _T_35027; // @[Switch.scala 30:36:@14549.4]
  assign _T_35030 = io_inAddr_17 == 6'h2d; // @[Switch.scala 30:53:@14551.4]
  assign valid_45_17 = io_inValid_17 & _T_35030; // @[Switch.scala 30:36:@14552.4]
  assign _T_35033 = io_inAddr_18 == 6'h2d; // @[Switch.scala 30:53:@14554.4]
  assign valid_45_18 = io_inValid_18 & _T_35033; // @[Switch.scala 30:36:@14555.4]
  assign _T_35036 = io_inAddr_19 == 6'h2d; // @[Switch.scala 30:53:@14557.4]
  assign valid_45_19 = io_inValid_19 & _T_35036; // @[Switch.scala 30:36:@14558.4]
  assign _T_35039 = io_inAddr_20 == 6'h2d; // @[Switch.scala 30:53:@14560.4]
  assign valid_45_20 = io_inValid_20 & _T_35039; // @[Switch.scala 30:36:@14561.4]
  assign _T_35042 = io_inAddr_21 == 6'h2d; // @[Switch.scala 30:53:@14563.4]
  assign valid_45_21 = io_inValid_21 & _T_35042; // @[Switch.scala 30:36:@14564.4]
  assign _T_35045 = io_inAddr_22 == 6'h2d; // @[Switch.scala 30:53:@14566.4]
  assign valid_45_22 = io_inValid_22 & _T_35045; // @[Switch.scala 30:36:@14567.4]
  assign _T_35048 = io_inAddr_23 == 6'h2d; // @[Switch.scala 30:53:@14569.4]
  assign valid_45_23 = io_inValid_23 & _T_35048; // @[Switch.scala 30:36:@14570.4]
  assign _T_35051 = io_inAddr_24 == 6'h2d; // @[Switch.scala 30:53:@14572.4]
  assign valid_45_24 = io_inValid_24 & _T_35051; // @[Switch.scala 30:36:@14573.4]
  assign _T_35054 = io_inAddr_25 == 6'h2d; // @[Switch.scala 30:53:@14575.4]
  assign valid_45_25 = io_inValid_25 & _T_35054; // @[Switch.scala 30:36:@14576.4]
  assign _T_35057 = io_inAddr_26 == 6'h2d; // @[Switch.scala 30:53:@14578.4]
  assign valid_45_26 = io_inValid_26 & _T_35057; // @[Switch.scala 30:36:@14579.4]
  assign _T_35060 = io_inAddr_27 == 6'h2d; // @[Switch.scala 30:53:@14581.4]
  assign valid_45_27 = io_inValid_27 & _T_35060; // @[Switch.scala 30:36:@14582.4]
  assign _T_35063 = io_inAddr_28 == 6'h2d; // @[Switch.scala 30:53:@14584.4]
  assign valid_45_28 = io_inValid_28 & _T_35063; // @[Switch.scala 30:36:@14585.4]
  assign _T_35066 = io_inAddr_29 == 6'h2d; // @[Switch.scala 30:53:@14587.4]
  assign valid_45_29 = io_inValid_29 & _T_35066; // @[Switch.scala 30:36:@14588.4]
  assign _T_35069 = io_inAddr_30 == 6'h2d; // @[Switch.scala 30:53:@14590.4]
  assign valid_45_30 = io_inValid_30 & _T_35069; // @[Switch.scala 30:36:@14591.4]
  assign _T_35072 = io_inAddr_31 == 6'h2d; // @[Switch.scala 30:53:@14593.4]
  assign valid_45_31 = io_inValid_31 & _T_35072; // @[Switch.scala 30:36:@14594.4]
  assign _T_35075 = io_inAddr_32 == 6'h2d; // @[Switch.scala 30:53:@14596.4]
  assign valid_45_32 = io_inValid_32 & _T_35075; // @[Switch.scala 30:36:@14597.4]
  assign _T_35078 = io_inAddr_33 == 6'h2d; // @[Switch.scala 30:53:@14599.4]
  assign valid_45_33 = io_inValid_33 & _T_35078; // @[Switch.scala 30:36:@14600.4]
  assign _T_35081 = io_inAddr_34 == 6'h2d; // @[Switch.scala 30:53:@14602.4]
  assign valid_45_34 = io_inValid_34 & _T_35081; // @[Switch.scala 30:36:@14603.4]
  assign _T_35084 = io_inAddr_35 == 6'h2d; // @[Switch.scala 30:53:@14605.4]
  assign valid_45_35 = io_inValid_35 & _T_35084; // @[Switch.scala 30:36:@14606.4]
  assign _T_35087 = io_inAddr_36 == 6'h2d; // @[Switch.scala 30:53:@14608.4]
  assign valid_45_36 = io_inValid_36 & _T_35087; // @[Switch.scala 30:36:@14609.4]
  assign _T_35090 = io_inAddr_37 == 6'h2d; // @[Switch.scala 30:53:@14611.4]
  assign valid_45_37 = io_inValid_37 & _T_35090; // @[Switch.scala 30:36:@14612.4]
  assign _T_35093 = io_inAddr_38 == 6'h2d; // @[Switch.scala 30:53:@14614.4]
  assign valid_45_38 = io_inValid_38 & _T_35093; // @[Switch.scala 30:36:@14615.4]
  assign _T_35096 = io_inAddr_39 == 6'h2d; // @[Switch.scala 30:53:@14617.4]
  assign valid_45_39 = io_inValid_39 & _T_35096; // @[Switch.scala 30:36:@14618.4]
  assign _T_35099 = io_inAddr_40 == 6'h2d; // @[Switch.scala 30:53:@14620.4]
  assign valid_45_40 = io_inValid_40 & _T_35099; // @[Switch.scala 30:36:@14621.4]
  assign _T_35102 = io_inAddr_41 == 6'h2d; // @[Switch.scala 30:53:@14623.4]
  assign valid_45_41 = io_inValid_41 & _T_35102; // @[Switch.scala 30:36:@14624.4]
  assign _T_35105 = io_inAddr_42 == 6'h2d; // @[Switch.scala 30:53:@14626.4]
  assign valid_45_42 = io_inValid_42 & _T_35105; // @[Switch.scala 30:36:@14627.4]
  assign _T_35108 = io_inAddr_43 == 6'h2d; // @[Switch.scala 30:53:@14629.4]
  assign valid_45_43 = io_inValid_43 & _T_35108; // @[Switch.scala 30:36:@14630.4]
  assign _T_35111 = io_inAddr_44 == 6'h2d; // @[Switch.scala 30:53:@14632.4]
  assign valid_45_44 = io_inValid_44 & _T_35111; // @[Switch.scala 30:36:@14633.4]
  assign _T_35114 = io_inAddr_45 == 6'h2d; // @[Switch.scala 30:53:@14635.4]
  assign valid_45_45 = io_inValid_45 & _T_35114; // @[Switch.scala 30:36:@14636.4]
  assign _T_35117 = io_inAddr_46 == 6'h2d; // @[Switch.scala 30:53:@14638.4]
  assign valid_45_46 = io_inValid_46 & _T_35117; // @[Switch.scala 30:36:@14639.4]
  assign _T_35120 = io_inAddr_47 == 6'h2d; // @[Switch.scala 30:53:@14641.4]
  assign valid_45_47 = io_inValid_47 & _T_35120; // @[Switch.scala 30:36:@14642.4]
  assign _T_35123 = io_inAddr_48 == 6'h2d; // @[Switch.scala 30:53:@14644.4]
  assign valid_45_48 = io_inValid_48 & _T_35123; // @[Switch.scala 30:36:@14645.4]
  assign _T_35126 = io_inAddr_49 == 6'h2d; // @[Switch.scala 30:53:@14647.4]
  assign valid_45_49 = io_inValid_49 & _T_35126; // @[Switch.scala 30:36:@14648.4]
  assign _T_35129 = io_inAddr_50 == 6'h2d; // @[Switch.scala 30:53:@14650.4]
  assign valid_45_50 = io_inValid_50 & _T_35129; // @[Switch.scala 30:36:@14651.4]
  assign _T_35132 = io_inAddr_51 == 6'h2d; // @[Switch.scala 30:53:@14653.4]
  assign valid_45_51 = io_inValid_51 & _T_35132; // @[Switch.scala 30:36:@14654.4]
  assign _T_35135 = io_inAddr_52 == 6'h2d; // @[Switch.scala 30:53:@14656.4]
  assign valid_45_52 = io_inValid_52 & _T_35135; // @[Switch.scala 30:36:@14657.4]
  assign _T_35138 = io_inAddr_53 == 6'h2d; // @[Switch.scala 30:53:@14659.4]
  assign valid_45_53 = io_inValid_53 & _T_35138; // @[Switch.scala 30:36:@14660.4]
  assign _T_35141 = io_inAddr_54 == 6'h2d; // @[Switch.scala 30:53:@14662.4]
  assign valid_45_54 = io_inValid_54 & _T_35141; // @[Switch.scala 30:36:@14663.4]
  assign _T_35144 = io_inAddr_55 == 6'h2d; // @[Switch.scala 30:53:@14665.4]
  assign valid_45_55 = io_inValid_55 & _T_35144; // @[Switch.scala 30:36:@14666.4]
  assign _T_35147 = io_inAddr_56 == 6'h2d; // @[Switch.scala 30:53:@14668.4]
  assign valid_45_56 = io_inValid_56 & _T_35147; // @[Switch.scala 30:36:@14669.4]
  assign _T_35150 = io_inAddr_57 == 6'h2d; // @[Switch.scala 30:53:@14671.4]
  assign valid_45_57 = io_inValid_57 & _T_35150; // @[Switch.scala 30:36:@14672.4]
  assign _T_35153 = io_inAddr_58 == 6'h2d; // @[Switch.scala 30:53:@14674.4]
  assign valid_45_58 = io_inValid_58 & _T_35153; // @[Switch.scala 30:36:@14675.4]
  assign _T_35156 = io_inAddr_59 == 6'h2d; // @[Switch.scala 30:53:@14677.4]
  assign valid_45_59 = io_inValid_59 & _T_35156; // @[Switch.scala 30:36:@14678.4]
  assign _T_35159 = io_inAddr_60 == 6'h2d; // @[Switch.scala 30:53:@14680.4]
  assign valid_45_60 = io_inValid_60 & _T_35159; // @[Switch.scala 30:36:@14681.4]
  assign _T_35162 = io_inAddr_61 == 6'h2d; // @[Switch.scala 30:53:@14683.4]
  assign valid_45_61 = io_inValid_61 & _T_35162; // @[Switch.scala 30:36:@14684.4]
  assign _T_35165 = io_inAddr_62 == 6'h2d; // @[Switch.scala 30:53:@14686.4]
  assign valid_45_62 = io_inValid_62 & _T_35165; // @[Switch.scala 30:36:@14687.4]
  assign _T_35168 = io_inAddr_63 == 6'h2d; // @[Switch.scala 30:53:@14689.4]
  assign valid_45_63 = io_inValid_63 & _T_35168; // @[Switch.scala 30:36:@14690.4]
  assign _T_35234 = valid_45_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@14692.4]
  assign _T_35235 = valid_45_61 ? 6'h3d : _T_35234; // @[Mux.scala 31:69:@14693.4]
  assign _T_35236 = valid_45_60 ? 6'h3c : _T_35235; // @[Mux.scala 31:69:@14694.4]
  assign _T_35237 = valid_45_59 ? 6'h3b : _T_35236; // @[Mux.scala 31:69:@14695.4]
  assign _T_35238 = valid_45_58 ? 6'h3a : _T_35237; // @[Mux.scala 31:69:@14696.4]
  assign _T_35239 = valid_45_57 ? 6'h39 : _T_35238; // @[Mux.scala 31:69:@14697.4]
  assign _T_35240 = valid_45_56 ? 6'h38 : _T_35239; // @[Mux.scala 31:69:@14698.4]
  assign _T_35241 = valid_45_55 ? 6'h37 : _T_35240; // @[Mux.scala 31:69:@14699.4]
  assign _T_35242 = valid_45_54 ? 6'h36 : _T_35241; // @[Mux.scala 31:69:@14700.4]
  assign _T_35243 = valid_45_53 ? 6'h35 : _T_35242; // @[Mux.scala 31:69:@14701.4]
  assign _T_35244 = valid_45_52 ? 6'h34 : _T_35243; // @[Mux.scala 31:69:@14702.4]
  assign _T_35245 = valid_45_51 ? 6'h33 : _T_35244; // @[Mux.scala 31:69:@14703.4]
  assign _T_35246 = valid_45_50 ? 6'h32 : _T_35245; // @[Mux.scala 31:69:@14704.4]
  assign _T_35247 = valid_45_49 ? 6'h31 : _T_35246; // @[Mux.scala 31:69:@14705.4]
  assign _T_35248 = valid_45_48 ? 6'h30 : _T_35247; // @[Mux.scala 31:69:@14706.4]
  assign _T_35249 = valid_45_47 ? 6'h2f : _T_35248; // @[Mux.scala 31:69:@14707.4]
  assign _T_35250 = valid_45_46 ? 6'h2e : _T_35249; // @[Mux.scala 31:69:@14708.4]
  assign _T_35251 = valid_45_45 ? 6'h2d : _T_35250; // @[Mux.scala 31:69:@14709.4]
  assign _T_35252 = valid_45_44 ? 6'h2c : _T_35251; // @[Mux.scala 31:69:@14710.4]
  assign _T_35253 = valid_45_43 ? 6'h2b : _T_35252; // @[Mux.scala 31:69:@14711.4]
  assign _T_35254 = valid_45_42 ? 6'h2a : _T_35253; // @[Mux.scala 31:69:@14712.4]
  assign _T_35255 = valid_45_41 ? 6'h29 : _T_35254; // @[Mux.scala 31:69:@14713.4]
  assign _T_35256 = valid_45_40 ? 6'h28 : _T_35255; // @[Mux.scala 31:69:@14714.4]
  assign _T_35257 = valid_45_39 ? 6'h27 : _T_35256; // @[Mux.scala 31:69:@14715.4]
  assign _T_35258 = valid_45_38 ? 6'h26 : _T_35257; // @[Mux.scala 31:69:@14716.4]
  assign _T_35259 = valid_45_37 ? 6'h25 : _T_35258; // @[Mux.scala 31:69:@14717.4]
  assign _T_35260 = valid_45_36 ? 6'h24 : _T_35259; // @[Mux.scala 31:69:@14718.4]
  assign _T_35261 = valid_45_35 ? 6'h23 : _T_35260; // @[Mux.scala 31:69:@14719.4]
  assign _T_35262 = valid_45_34 ? 6'h22 : _T_35261; // @[Mux.scala 31:69:@14720.4]
  assign _T_35263 = valid_45_33 ? 6'h21 : _T_35262; // @[Mux.scala 31:69:@14721.4]
  assign _T_35264 = valid_45_32 ? 6'h20 : _T_35263; // @[Mux.scala 31:69:@14722.4]
  assign _T_35265 = valid_45_31 ? 6'h1f : _T_35264; // @[Mux.scala 31:69:@14723.4]
  assign _T_35266 = valid_45_30 ? 6'h1e : _T_35265; // @[Mux.scala 31:69:@14724.4]
  assign _T_35267 = valid_45_29 ? 6'h1d : _T_35266; // @[Mux.scala 31:69:@14725.4]
  assign _T_35268 = valid_45_28 ? 6'h1c : _T_35267; // @[Mux.scala 31:69:@14726.4]
  assign _T_35269 = valid_45_27 ? 6'h1b : _T_35268; // @[Mux.scala 31:69:@14727.4]
  assign _T_35270 = valid_45_26 ? 6'h1a : _T_35269; // @[Mux.scala 31:69:@14728.4]
  assign _T_35271 = valid_45_25 ? 6'h19 : _T_35270; // @[Mux.scala 31:69:@14729.4]
  assign _T_35272 = valid_45_24 ? 6'h18 : _T_35271; // @[Mux.scala 31:69:@14730.4]
  assign _T_35273 = valid_45_23 ? 6'h17 : _T_35272; // @[Mux.scala 31:69:@14731.4]
  assign _T_35274 = valid_45_22 ? 6'h16 : _T_35273; // @[Mux.scala 31:69:@14732.4]
  assign _T_35275 = valid_45_21 ? 6'h15 : _T_35274; // @[Mux.scala 31:69:@14733.4]
  assign _T_35276 = valid_45_20 ? 6'h14 : _T_35275; // @[Mux.scala 31:69:@14734.4]
  assign _T_35277 = valid_45_19 ? 6'h13 : _T_35276; // @[Mux.scala 31:69:@14735.4]
  assign _T_35278 = valid_45_18 ? 6'h12 : _T_35277; // @[Mux.scala 31:69:@14736.4]
  assign _T_35279 = valid_45_17 ? 6'h11 : _T_35278; // @[Mux.scala 31:69:@14737.4]
  assign _T_35280 = valid_45_16 ? 6'h10 : _T_35279; // @[Mux.scala 31:69:@14738.4]
  assign _T_35281 = valid_45_15 ? 6'hf : _T_35280; // @[Mux.scala 31:69:@14739.4]
  assign _T_35282 = valid_45_14 ? 6'he : _T_35281; // @[Mux.scala 31:69:@14740.4]
  assign _T_35283 = valid_45_13 ? 6'hd : _T_35282; // @[Mux.scala 31:69:@14741.4]
  assign _T_35284 = valid_45_12 ? 6'hc : _T_35283; // @[Mux.scala 31:69:@14742.4]
  assign _T_35285 = valid_45_11 ? 6'hb : _T_35284; // @[Mux.scala 31:69:@14743.4]
  assign _T_35286 = valid_45_10 ? 6'ha : _T_35285; // @[Mux.scala 31:69:@14744.4]
  assign _T_35287 = valid_45_9 ? 6'h9 : _T_35286; // @[Mux.scala 31:69:@14745.4]
  assign _T_35288 = valid_45_8 ? 6'h8 : _T_35287; // @[Mux.scala 31:69:@14746.4]
  assign _T_35289 = valid_45_7 ? 6'h7 : _T_35288; // @[Mux.scala 31:69:@14747.4]
  assign _T_35290 = valid_45_6 ? 6'h6 : _T_35289; // @[Mux.scala 31:69:@14748.4]
  assign _T_35291 = valid_45_5 ? 6'h5 : _T_35290; // @[Mux.scala 31:69:@14749.4]
  assign _T_35292 = valid_45_4 ? 6'h4 : _T_35291; // @[Mux.scala 31:69:@14750.4]
  assign _T_35293 = valid_45_3 ? 6'h3 : _T_35292; // @[Mux.scala 31:69:@14751.4]
  assign _T_35294 = valid_45_2 ? 6'h2 : _T_35293; // @[Mux.scala 31:69:@14752.4]
  assign _T_35295 = valid_45_1 ? 6'h1 : _T_35294; // @[Mux.scala 31:69:@14753.4]
  assign select_45 = valid_45_0 ? 6'h0 : _T_35295; // @[Mux.scala 31:69:@14754.4]
  assign _GEN_2881 = 6'h1 == select_45 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2882 = 6'h2 == select_45 ? io_inData_2 : _GEN_2881; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2883 = 6'h3 == select_45 ? io_inData_3 : _GEN_2882; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2884 = 6'h4 == select_45 ? io_inData_4 : _GEN_2883; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2885 = 6'h5 == select_45 ? io_inData_5 : _GEN_2884; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2886 = 6'h6 == select_45 ? io_inData_6 : _GEN_2885; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2887 = 6'h7 == select_45 ? io_inData_7 : _GEN_2886; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2888 = 6'h8 == select_45 ? io_inData_8 : _GEN_2887; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2889 = 6'h9 == select_45 ? io_inData_9 : _GEN_2888; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2890 = 6'ha == select_45 ? io_inData_10 : _GEN_2889; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2891 = 6'hb == select_45 ? io_inData_11 : _GEN_2890; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2892 = 6'hc == select_45 ? io_inData_12 : _GEN_2891; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2893 = 6'hd == select_45 ? io_inData_13 : _GEN_2892; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2894 = 6'he == select_45 ? io_inData_14 : _GEN_2893; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2895 = 6'hf == select_45 ? io_inData_15 : _GEN_2894; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2896 = 6'h10 == select_45 ? io_inData_16 : _GEN_2895; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2897 = 6'h11 == select_45 ? io_inData_17 : _GEN_2896; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2898 = 6'h12 == select_45 ? io_inData_18 : _GEN_2897; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2899 = 6'h13 == select_45 ? io_inData_19 : _GEN_2898; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2900 = 6'h14 == select_45 ? io_inData_20 : _GEN_2899; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2901 = 6'h15 == select_45 ? io_inData_21 : _GEN_2900; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2902 = 6'h16 == select_45 ? io_inData_22 : _GEN_2901; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2903 = 6'h17 == select_45 ? io_inData_23 : _GEN_2902; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2904 = 6'h18 == select_45 ? io_inData_24 : _GEN_2903; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2905 = 6'h19 == select_45 ? io_inData_25 : _GEN_2904; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2906 = 6'h1a == select_45 ? io_inData_26 : _GEN_2905; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2907 = 6'h1b == select_45 ? io_inData_27 : _GEN_2906; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2908 = 6'h1c == select_45 ? io_inData_28 : _GEN_2907; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2909 = 6'h1d == select_45 ? io_inData_29 : _GEN_2908; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2910 = 6'h1e == select_45 ? io_inData_30 : _GEN_2909; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2911 = 6'h1f == select_45 ? io_inData_31 : _GEN_2910; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2912 = 6'h20 == select_45 ? io_inData_32 : _GEN_2911; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2913 = 6'h21 == select_45 ? io_inData_33 : _GEN_2912; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2914 = 6'h22 == select_45 ? io_inData_34 : _GEN_2913; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2915 = 6'h23 == select_45 ? io_inData_35 : _GEN_2914; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2916 = 6'h24 == select_45 ? io_inData_36 : _GEN_2915; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2917 = 6'h25 == select_45 ? io_inData_37 : _GEN_2916; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2918 = 6'h26 == select_45 ? io_inData_38 : _GEN_2917; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2919 = 6'h27 == select_45 ? io_inData_39 : _GEN_2918; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2920 = 6'h28 == select_45 ? io_inData_40 : _GEN_2919; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2921 = 6'h29 == select_45 ? io_inData_41 : _GEN_2920; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2922 = 6'h2a == select_45 ? io_inData_42 : _GEN_2921; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2923 = 6'h2b == select_45 ? io_inData_43 : _GEN_2922; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2924 = 6'h2c == select_45 ? io_inData_44 : _GEN_2923; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2925 = 6'h2d == select_45 ? io_inData_45 : _GEN_2924; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2926 = 6'h2e == select_45 ? io_inData_46 : _GEN_2925; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2927 = 6'h2f == select_45 ? io_inData_47 : _GEN_2926; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2928 = 6'h30 == select_45 ? io_inData_48 : _GEN_2927; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2929 = 6'h31 == select_45 ? io_inData_49 : _GEN_2928; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2930 = 6'h32 == select_45 ? io_inData_50 : _GEN_2929; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2931 = 6'h33 == select_45 ? io_inData_51 : _GEN_2930; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2932 = 6'h34 == select_45 ? io_inData_52 : _GEN_2931; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2933 = 6'h35 == select_45 ? io_inData_53 : _GEN_2932; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2934 = 6'h36 == select_45 ? io_inData_54 : _GEN_2933; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2935 = 6'h37 == select_45 ? io_inData_55 : _GEN_2934; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2936 = 6'h38 == select_45 ? io_inData_56 : _GEN_2935; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2937 = 6'h39 == select_45 ? io_inData_57 : _GEN_2936; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2938 = 6'h3a == select_45 ? io_inData_58 : _GEN_2937; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2939 = 6'h3b == select_45 ? io_inData_59 : _GEN_2938; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2940 = 6'h3c == select_45 ? io_inData_60 : _GEN_2939; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2941 = 6'h3d == select_45 ? io_inData_61 : _GEN_2940; // @[Switch.scala 33:19:@14756.4]
  assign _GEN_2942 = 6'h3e == select_45 ? io_inData_62 : _GEN_2941; // @[Switch.scala 33:19:@14756.4]
  assign _T_35304 = {valid_45_7,valid_45_6,valid_45_5,valid_45_4,valid_45_3,valid_45_2,valid_45_1,valid_45_0}; // @[Switch.scala 34:32:@14763.4]
  assign _T_35312 = {valid_45_15,valid_45_14,valid_45_13,valid_45_12,valid_45_11,valid_45_10,valid_45_9,valid_45_8,_T_35304}; // @[Switch.scala 34:32:@14771.4]
  assign _T_35319 = {valid_45_23,valid_45_22,valid_45_21,valid_45_20,valid_45_19,valid_45_18,valid_45_17,valid_45_16}; // @[Switch.scala 34:32:@14778.4]
  assign _T_35328 = {valid_45_31,valid_45_30,valid_45_29,valid_45_28,valid_45_27,valid_45_26,valid_45_25,valid_45_24,_T_35319,_T_35312}; // @[Switch.scala 34:32:@14787.4]
  assign _T_35335 = {valid_45_39,valid_45_38,valid_45_37,valid_45_36,valid_45_35,valid_45_34,valid_45_33,valid_45_32}; // @[Switch.scala 34:32:@14794.4]
  assign _T_35343 = {valid_45_47,valid_45_46,valid_45_45,valid_45_44,valid_45_43,valid_45_42,valid_45_41,valid_45_40,_T_35335}; // @[Switch.scala 34:32:@14802.4]
  assign _T_35350 = {valid_45_55,valid_45_54,valid_45_53,valid_45_52,valid_45_51,valid_45_50,valid_45_49,valid_45_48}; // @[Switch.scala 34:32:@14809.4]
  assign _T_35359 = {valid_45_63,valid_45_62,valid_45_61,valid_45_60,valid_45_59,valid_45_58,valid_45_57,valid_45_56,_T_35350,_T_35343}; // @[Switch.scala 34:32:@14818.4]
  assign _T_35360 = {_T_35359,_T_35328}; // @[Switch.scala 34:32:@14819.4]
  assign _T_35364 = io_inAddr_0 == 6'h2e; // @[Switch.scala 30:53:@14822.4]
  assign valid_46_0 = io_inValid_0 & _T_35364; // @[Switch.scala 30:36:@14823.4]
  assign _T_35367 = io_inAddr_1 == 6'h2e; // @[Switch.scala 30:53:@14825.4]
  assign valid_46_1 = io_inValid_1 & _T_35367; // @[Switch.scala 30:36:@14826.4]
  assign _T_35370 = io_inAddr_2 == 6'h2e; // @[Switch.scala 30:53:@14828.4]
  assign valid_46_2 = io_inValid_2 & _T_35370; // @[Switch.scala 30:36:@14829.4]
  assign _T_35373 = io_inAddr_3 == 6'h2e; // @[Switch.scala 30:53:@14831.4]
  assign valid_46_3 = io_inValid_3 & _T_35373; // @[Switch.scala 30:36:@14832.4]
  assign _T_35376 = io_inAddr_4 == 6'h2e; // @[Switch.scala 30:53:@14834.4]
  assign valid_46_4 = io_inValid_4 & _T_35376; // @[Switch.scala 30:36:@14835.4]
  assign _T_35379 = io_inAddr_5 == 6'h2e; // @[Switch.scala 30:53:@14837.4]
  assign valid_46_5 = io_inValid_5 & _T_35379; // @[Switch.scala 30:36:@14838.4]
  assign _T_35382 = io_inAddr_6 == 6'h2e; // @[Switch.scala 30:53:@14840.4]
  assign valid_46_6 = io_inValid_6 & _T_35382; // @[Switch.scala 30:36:@14841.4]
  assign _T_35385 = io_inAddr_7 == 6'h2e; // @[Switch.scala 30:53:@14843.4]
  assign valid_46_7 = io_inValid_7 & _T_35385; // @[Switch.scala 30:36:@14844.4]
  assign _T_35388 = io_inAddr_8 == 6'h2e; // @[Switch.scala 30:53:@14846.4]
  assign valid_46_8 = io_inValid_8 & _T_35388; // @[Switch.scala 30:36:@14847.4]
  assign _T_35391 = io_inAddr_9 == 6'h2e; // @[Switch.scala 30:53:@14849.4]
  assign valid_46_9 = io_inValid_9 & _T_35391; // @[Switch.scala 30:36:@14850.4]
  assign _T_35394 = io_inAddr_10 == 6'h2e; // @[Switch.scala 30:53:@14852.4]
  assign valid_46_10 = io_inValid_10 & _T_35394; // @[Switch.scala 30:36:@14853.4]
  assign _T_35397 = io_inAddr_11 == 6'h2e; // @[Switch.scala 30:53:@14855.4]
  assign valid_46_11 = io_inValid_11 & _T_35397; // @[Switch.scala 30:36:@14856.4]
  assign _T_35400 = io_inAddr_12 == 6'h2e; // @[Switch.scala 30:53:@14858.4]
  assign valid_46_12 = io_inValid_12 & _T_35400; // @[Switch.scala 30:36:@14859.4]
  assign _T_35403 = io_inAddr_13 == 6'h2e; // @[Switch.scala 30:53:@14861.4]
  assign valid_46_13 = io_inValid_13 & _T_35403; // @[Switch.scala 30:36:@14862.4]
  assign _T_35406 = io_inAddr_14 == 6'h2e; // @[Switch.scala 30:53:@14864.4]
  assign valid_46_14 = io_inValid_14 & _T_35406; // @[Switch.scala 30:36:@14865.4]
  assign _T_35409 = io_inAddr_15 == 6'h2e; // @[Switch.scala 30:53:@14867.4]
  assign valid_46_15 = io_inValid_15 & _T_35409; // @[Switch.scala 30:36:@14868.4]
  assign _T_35412 = io_inAddr_16 == 6'h2e; // @[Switch.scala 30:53:@14870.4]
  assign valid_46_16 = io_inValid_16 & _T_35412; // @[Switch.scala 30:36:@14871.4]
  assign _T_35415 = io_inAddr_17 == 6'h2e; // @[Switch.scala 30:53:@14873.4]
  assign valid_46_17 = io_inValid_17 & _T_35415; // @[Switch.scala 30:36:@14874.4]
  assign _T_35418 = io_inAddr_18 == 6'h2e; // @[Switch.scala 30:53:@14876.4]
  assign valid_46_18 = io_inValid_18 & _T_35418; // @[Switch.scala 30:36:@14877.4]
  assign _T_35421 = io_inAddr_19 == 6'h2e; // @[Switch.scala 30:53:@14879.4]
  assign valid_46_19 = io_inValid_19 & _T_35421; // @[Switch.scala 30:36:@14880.4]
  assign _T_35424 = io_inAddr_20 == 6'h2e; // @[Switch.scala 30:53:@14882.4]
  assign valid_46_20 = io_inValid_20 & _T_35424; // @[Switch.scala 30:36:@14883.4]
  assign _T_35427 = io_inAddr_21 == 6'h2e; // @[Switch.scala 30:53:@14885.4]
  assign valid_46_21 = io_inValid_21 & _T_35427; // @[Switch.scala 30:36:@14886.4]
  assign _T_35430 = io_inAddr_22 == 6'h2e; // @[Switch.scala 30:53:@14888.4]
  assign valid_46_22 = io_inValid_22 & _T_35430; // @[Switch.scala 30:36:@14889.4]
  assign _T_35433 = io_inAddr_23 == 6'h2e; // @[Switch.scala 30:53:@14891.4]
  assign valid_46_23 = io_inValid_23 & _T_35433; // @[Switch.scala 30:36:@14892.4]
  assign _T_35436 = io_inAddr_24 == 6'h2e; // @[Switch.scala 30:53:@14894.4]
  assign valid_46_24 = io_inValid_24 & _T_35436; // @[Switch.scala 30:36:@14895.4]
  assign _T_35439 = io_inAddr_25 == 6'h2e; // @[Switch.scala 30:53:@14897.4]
  assign valid_46_25 = io_inValid_25 & _T_35439; // @[Switch.scala 30:36:@14898.4]
  assign _T_35442 = io_inAddr_26 == 6'h2e; // @[Switch.scala 30:53:@14900.4]
  assign valid_46_26 = io_inValid_26 & _T_35442; // @[Switch.scala 30:36:@14901.4]
  assign _T_35445 = io_inAddr_27 == 6'h2e; // @[Switch.scala 30:53:@14903.4]
  assign valid_46_27 = io_inValid_27 & _T_35445; // @[Switch.scala 30:36:@14904.4]
  assign _T_35448 = io_inAddr_28 == 6'h2e; // @[Switch.scala 30:53:@14906.4]
  assign valid_46_28 = io_inValid_28 & _T_35448; // @[Switch.scala 30:36:@14907.4]
  assign _T_35451 = io_inAddr_29 == 6'h2e; // @[Switch.scala 30:53:@14909.4]
  assign valid_46_29 = io_inValid_29 & _T_35451; // @[Switch.scala 30:36:@14910.4]
  assign _T_35454 = io_inAddr_30 == 6'h2e; // @[Switch.scala 30:53:@14912.4]
  assign valid_46_30 = io_inValid_30 & _T_35454; // @[Switch.scala 30:36:@14913.4]
  assign _T_35457 = io_inAddr_31 == 6'h2e; // @[Switch.scala 30:53:@14915.4]
  assign valid_46_31 = io_inValid_31 & _T_35457; // @[Switch.scala 30:36:@14916.4]
  assign _T_35460 = io_inAddr_32 == 6'h2e; // @[Switch.scala 30:53:@14918.4]
  assign valid_46_32 = io_inValid_32 & _T_35460; // @[Switch.scala 30:36:@14919.4]
  assign _T_35463 = io_inAddr_33 == 6'h2e; // @[Switch.scala 30:53:@14921.4]
  assign valid_46_33 = io_inValid_33 & _T_35463; // @[Switch.scala 30:36:@14922.4]
  assign _T_35466 = io_inAddr_34 == 6'h2e; // @[Switch.scala 30:53:@14924.4]
  assign valid_46_34 = io_inValid_34 & _T_35466; // @[Switch.scala 30:36:@14925.4]
  assign _T_35469 = io_inAddr_35 == 6'h2e; // @[Switch.scala 30:53:@14927.4]
  assign valid_46_35 = io_inValid_35 & _T_35469; // @[Switch.scala 30:36:@14928.4]
  assign _T_35472 = io_inAddr_36 == 6'h2e; // @[Switch.scala 30:53:@14930.4]
  assign valid_46_36 = io_inValid_36 & _T_35472; // @[Switch.scala 30:36:@14931.4]
  assign _T_35475 = io_inAddr_37 == 6'h2e; // @[Switch.scala 30:53:@14933.4]
  assign valid_46_37 = io_inValid_37 & _T_35475; // @[Switch.scala 30:36:@14934.4]
  assign _T_35478 = io_inAddr_38 == 6'h2e; // @[Switch.scala 30:53:@14936.4]
  assign valid_46_38 = io_inValid_38 & _T_35478; // @[Switch.scala 30:36:@14937.4]
  assign _T_35481 = io_inAddr_39 == 6'h2e; // @[Switch.scala 30:53:@14939.4]
  assign valid_46_39 = io_inValid_39 & _T_35481; // @[Switch.scala 30:36:@14940.4]
  assign _T_35484 = io_inAddr_40 == 6'h2e; // @[Switch.scala 30:53:@14942.4]
  assign valid_46_40 = io_inValid_40 & _T_35484; // @[Switch.scala 30:36:@14943.4]
  assign _T_35487 = io_inAddr_41 == 6'h2e; // @[Switch.scala 30:53:@14945.4]
  assign valid_46_41 = io_inValid_41 & _T_35487; // @[Switch.scala 30:36:@14946.4]
  assign _T_35490 = io_inAddr_42 == 6'h2e; // @[Switch.scala 30:53:@14948.4]
  assign valid_46_42 = io_inValid_42 & _T_35490; // @[Switch.scala 30:36:@14949.4]
  assign _T_35493 = io_inAddr_43 == 6'h2e; // @[Switch.scala 30:53:@14951.4]
  assign valid_46_43 = io_inValid_43 & _T_35493; // @[Switch.scala 30:36:@14952.4]
  assign _T_35496 = io_inAddr_44 == 6'h2e; // @[Switch.scala 30:53:@14954.4]
  assign valid_46_44 = io_inValid_44 & _T_35496; // @[Switch.scala 30:36:@14955.4]
  assign _T_35499 = io_inAddr_45 == 6'h2e; // @[Switch.scala 30:53:@14957.4]
  assign valid_46_45 = io_inValid_45 & _T_35499; // @[Switch.scala 30:36:@14958.4]
  assign _T_35502 = io_inAddr_46 == 6'h2e; // @[Switch.scala 30:53:@14960.4]
  assign valid_46_46 = io_inValid_46 & _T_35502; // @[Switch.scala 30:36:@14961.4]
  assign _T_35505 = io_inAddr_47 == 6'h2e; // @[Switch.scala 30:53:@14963.4]
  assign valid_46_47 = io_inValid_47 & _T_35505; // @[Switch.scala 30:36:@14964.4]
  assign _T_35508 = io_inAddr_48 == 6'h2e; // @[Switch.scala 30:53:@14966.4]
  assign valid_46_48 = io_inValid_48 & _T_35508; // @[Switch.scala 30:36:@14967.4]
  assign _T_35511 = io_inAddr_49 == 6'h2e; // @[Switch.scala 30:53:@14969.4]
  assign valid_46_49 = io_inValid_49 & _T_35511; // @[Switch.scala 30:36:@14970.4]
  assign _T_35514 = io_inAddr_50 == 6'h2e; // @[Switch.scala 30:53:@14972.4]
  assign valid_46_50 = io_inValid_50 & _T_35514; // @[Switch.scala 30:36:@14973.4]
  assign _T_35517 = io_inAddr_51 == 6'h2e; // @[Switch.scala 30:53:@14975.4]
  assign valid_46_51 = io_inValid_51 & _T_35517; // @[Switch.scala 30:36:@14976.4]
  assign _T_35520 = io_inAddr_52 == 6'h2e; // @[Switch.scala 30:53:@14978.4]
  assign valid_46_52 = io_inValid_52 & _T_35520; // @[Switch.scala 30:36:@14979.4]
  assign _T_35523 = io_inAddr_53 == 6'h2e; // @[Switch.scala 30:53:@14981.4]
  assign valid_46_53 = io_inValid_53 & _T_35523; // @[Switch.scala 30:36:@14982.4]
  assign _T_35526 = io_inAddr_54 == 6'h2e; // @[Switch.scala 30:53:@14984.4]
  assign valid_46_54 = io_inValid_54 & _T_35526; // @[Switch.scala 30:36:@14985.4]
  assign _T_35529 = io_inAddr_55 == 6'h2e; // @[Switch.scala 30:53:@14987.4]
  assign valid_46_55 = io_inValid_55 & _T_35529; // @[Switch.scala 30:36:@14988.4]
  assign _T_35532 = io_inAddr_56 == 6'h2e; // @[Switch.scala 30:53:@14990.4]
  assign valid_46_56 = io_inValid_56 & _T_35532; // @[Switch.scala 30:36:@14991.4]
  assign _T_35535 = io_inAddr_57 == 6'h2e; // @[Switch.scala 30:53:@14993.4]
  assign valid_46_57 = io_inValid_57 & _T_35535; // @[Switch.scala 30:36:@14994.4]
  assign _T_35538 = io_inAddr_58 == 6'h2e; // @[Switch.scala 30:53:@14996.4]
  assign valid_46_58 = io_inValid_58 & _T_35538; // @[Switch.scala 30:36:@14997.4]
  assign _T_35541 = io_inAddr_59 == 6'h2e; // @[Switch.scala 30:53:@14999.4]
  assign valid_46_59 = io_inValid_59 & _T_35541; // @[Switch.scala 30:36:@15000.4]
  assign _T_35544 = io_inAddr_60 == 6'h2e; // @[Switch.scala 30:53:@15002.4]
  assign valid_46_60 = io_inValid_60 & _T_35544; // @[Switch.scala 30:36:@15003.4]
  assign _T_35547 = io_inAddr_61 == 6'h2e; // @[Switch.scala 30:53:@15005.4]
  assign valid_46_61 = io_inValid_61 & _T_35547; // @[Switch.scala 30:36:@15006.4]
  assign _T_35550 = io_inAddr_62 == 6'h2e; // @[Switch.scala 30:53:@15008.4]
  assign valid_46_62 = io_inValid_62 & _T_35550; // @[Switch.scala 30:36:@15009.4]
  assign _T_35553 = io_inAddr_63 == 6'h2e; // @[Switch.scala 30:53:@15011.4]
  assign valid_46_63 = io_inValid_63 & _T_35553; // @[Switch.scala 30:36:@15012.4]
  assign _T_35619 = valid_46_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@15014.4]
  assign _T_35620 = valid_46_61 ? 6'h3d : _T_35619; // @[Mux.scala 31:69:@15015.4]
  assign _T_35621 = valid_46_60 ? 6'h3c : _T_35620; // @[Mux.scala 31:69:@15016.4]
  assign _T_35622 = valid_46_59 ? 6'h3b : _T_35621; // @[Mux.scala 31:69:@15017.4]
  assign _T_35623 = valid_46_58 ? 6'h3a : _T_35622; // @[Mux.scala 31:69:@15018.4]
  assign _T_35624 = valid_46_57 ? 6'h39 : _T_35623; // @[Mux.scala 31:69:@15019.4]
  assign _T_35625 = valid_46_56 ? 6'h38 : _T_35624; // @[Mux.scala 31:69:@15020.4]
  assign _T_35626 = valid_46_55 ? 6'h37 : _T_35625; // @[Mux.scala 31:69:@15021.4]
  assign _T_35627 = valid_46_54 ? 6'h36 : _T_35626; // @[Mux.scala 31:69:@15022.4]
  assign _T_35628 = valid_46_53 ? 6'h35 : _T_35627; // @[Mux.scala 31:69:@15023.4]
  assign _T_35629 = valid_46_52 ? 6'h34 : _T_35628; // @[Mux.scala 31:69:@15024.4]
  assign _T_35630 = valid_46_51 ? 6'h33 : _T_35629; // @[Mux.scala 31:69:@15025.4]
  assign _T_35631 = valid_46_50 ? 6'h32 : _T_35630; // @[Mux.scala 31:69:@15026.4]
  assign _T_35632 = valid_46_49 ? 6'h31 : _T_35631; // @[Mux.scala 31:69:@15027.4]
  assign _T_35633 = valid_46_48 ? 6'h30 : _T_35632; // @[Mux.scala 31:69:@15028.4]
  assign _T_35634 = valid_46_47 ? 6'h2f : _T_35633; // @[Mux.scala 31:69:@15029.4]
  assign _T_35635 = valid_46_46 ? 6'h2e : _T_35634; // @[Mux.scala 31:69:@15030.4]
  assign _T_35636 = valid_46_45 ? 6'h2d : _T_35635; // @[Mux.scala 31:69:@15031.4]
  assign _T_35637 = valid_46_44 ? 6'h2c : _T_35636; // @[Mux.scala 31:69:@15032.4]
  assign _T_35638 = valid_46_43 ? 6'h2b : _T_35637; // @[Mux.scala 31:69:@15033.4]
  assign _T_35639 = valid_46_42 ? 6'h2a : _T_35638; // @[Mux.scala 31:69:@15034.4]
  assign _T_35640 = valid_46_41 ? 6'h29 : _T_35639; // @[Mux.scala 31:69:@15035.4]
  assign _T_35641 = valid_46_40 ? 6'h28 : _T_35640; // @[Mux.scala 31:69:@15036.4]
  assign _T_35642 = valid_46_39 ? 6'h27 : _T_35641; // @[Mux.scala 31:69:@15037.4]
  assign _T_35643 = valid_46_38 ? 6'h26 : _T_35642; // @[Mux.scala 31:69:@15038.4]
  assign _T_35644 = valid_46_37 ? 6'h25 : _T_35643; // @[Mux.scala 31:69:@15039.4]
  assign _T_35645 = valid_46_36 ? 6'h24 : _T_35644; // @[Mux.scala 31:69:@15040.4]
  assign _T_35646 = valid_46_35 ? 6'h23 : _T_35645; // @[Mux.scala 31:69:@15041.4]
  assign _T_35647 = valid_46_34 ? 6'h22 : _T_35646; // @[Mux.scala 31:69:@15042.4]
  assign _T_35648 = valid_46_33 ? 6'h21 : _T_35647; // @[Mux.scala 31:69:@15043.4]
  assign _T_35649 = valid_46_32 ? 6'h20 : _T_35648; // @[Mux.scala 31:69:@15044.4]
  assign _T_35650 = valid_46_31 ? 6'h1f : _T_35649; // @[Mux.scala 31:69:@15045.4]
  assign _T_35651 = valid_46_30 ? 6'h1e : _T_35650; // @[Mux.scala 31:69:@15046.4]
  assign _T_35652 = valid_46_29 ? 6'h1d : _T_35651; // @[Mux.scala 31:69:@15047.4]
  assign _T_35653 = valid_46_28 ? 6'h1c : _T_35652; // @[Mux.scala 31:69:@15048.4]
  assign _T_35654 = valid_46_27 ? 6'h1b : _T_35653; // @[Mux.scala 31:69:@15049.4]
  assign _T_35655 = valid_46_26 ? 6'h1a : _T_35654; // @[Mux.scala 31:69:@15050.4]
  assign _T_35656 = valid_46_25 ? 6'h19 : _T_35655; // @[Mux.scala 31:69:@15051.4]
  assign _T_35657 = valid_46_24 ? 6'h18 : _T_35656; // @[Mux.scala 31:69:@15052.4]
  assign _T_35658 = valid_46_23 ? 6'h17 : _T_35657; // @[Mux.scala 31:69:@15053.4]
  assign _T_35659 = valid_46_22 ? 6'h16 : _T_35658; // @[Mux.scala 31:69:@15054.4]
  assign _T_35660 = valid_46_21 ? 6'h15 : _T_35659; // @[Mux.scala 31:69:@15055.4]
  assign _T_35661 = valid_46_20 ? 6'h14 : _T_35660; // @[Mux.scala 31:69:@15056.4]
  assign _T_35662 = valid_46_19 ? 6'h13 : _T_35661; // @[Mux.scala 31:69:@15057.4]
  assign _T_35663 = valid_46_18 ? 6'h12 : _T_35662; // @[Mux.scala 31:69:@15058.4]
  assign _T_35664 = valid_46_17 ? 6'h11 : _T_35663; // @[Mux.scala 31:69:@15059.4]
  assign _T_35665 = valid_46_16 ? 6'h10 : _T_35664; // @[Mux.scala 31:69:@15060.4]
  assign _T_35666 = valid_46_15 ? 6'hf : _T_35665; // @[Mux.scala 31:69:@15061.4]
  assign _T_35667 = valid_46_14 ? 6'he : _T_35666; // @[Mux.scala 31:69:@15062.4]
  assign _T_35668 = valid_46_13 ? 6'hd : _T_35667; // @[Mux.scala 31:69:@15063.4]
  assign _T_35669 = valid_46_12 ? 6'hc : _T_35668; // @[Mux.scala 31:69:@15064.4]
  assign _T_35670 = valid_46_11 ? 6'hb : _T_35669; // @[Mux.scala 31:69:@15065.4]
  assign _T_35671 = valid_46_10 ? 6'ha : _T_35670; // @[Mux.scala 31:69:@15066.4]
  assign _T_35672 = valid_46_9 ? 6'h9 : _T_35671; // @[Mux.scala 31:69:@15067.4]
  assign _T_35673 = valid_46_8 ? 6'h8 : _T_35672; // @[Mux.scala 31:69:@15068.4]
  assign _T_35674 = valid_46_7 ? 6'h7 : _T_35673; // @[Mux.scala 31:69:@15069.4]
  assign _T_35675 = valid_46_6 ? 6'h6 : _T_35674; // @[Mux.scala 31:69:@15070.4]
  assign _T_35676 = valid_46_5 ? 6'h5 : _T_35675; // @[Mux.scala 31:69:@15071.4]
  assign _T_35677 = valid_46_4 ? 6'h4 : _T_35676; // @[Mux.scala 31:69:@15072.4]
  assign _T_35678 = valid_46_3 ? 6'h3 : _T_35677; // @[Mux.scala 31:69:@15073.4]
  assign _T_35679 = valid_46_2 ? 6'h2 : _T_35678; // @[Mux.scala 31:69:@15074.4]
  assign _T_35680 = valid_46_1 ? 6'h1 : _T_35679; // @[Mux.scala 31:69:@15075.4]
  assign select_46 = valid_46_0 ? 6'h0 : _T_35680; // @[Mux.scala 31:69:@15076.4]
  assign _GEN_2945 = 6'h1 == select_46 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2946 = 6'h2 == select_46 ? io_inData_2 : _GEN_2945; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2947 = 6'h3 == select_46 ? io_inData_3 : _GEN_2946; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2948 = 6'h4 == select_46 ? io_inData_4 : _GEN_2947; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2949 = 6'h5 == select_46 ? io_inData_5 : _GEN_2948; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2950 = 6'h6 == select_46 ? io_inData_6 : _GEN_2949; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2951 = 6'h7 == select_46 ? io_inData_7 : _GEN_2950; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2952 = 6'h8 == select_46 ? io_inData_8 : _GEN_2951; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2953 = 6'h9 == select_46 ? io_inData_9 : _GEN_2952; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2954 = 6'ha == select_46 ? io_inData_10 : _GEN_2953; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2955 = 6'hb == select_46 ? io_inData_11 : _GEN_2954; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2956 = 6'hc == select_46 ? io_inData_12 : _GEN_2955; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2957 = 6'hd == select_46 ? io_inData_13 : _GEN_2956; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2958 = 6'he == select_46 ? io_inData_14 : _GEN_2957; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2959 = 6'hf == select_46 ? io_inData_15 : _GEN_2958; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2960 = 6'h10 == select_46 ? io_inData_16 : _GEN_2959; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2961 = 6'h11 == select_46 ? io_inData_17 : _GEN_2960; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2962 = 6'h12 == select_46 ? io_inData_18 : _GEN_2961; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2963 = 6'h13 == select_46 ? io_inData_19 : _GEN_2962; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2964 = 6'h14 == select_46 ? io_inData_20 : _GEN_2963; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2965 = 6'h15 == select_46 ? io_inData_21 : _GEN_2964; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2966 = 6'h16 == select_46 ? io_inData_22 : _GEN_2965; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2967 = 6'h17 == select_46 ? io_inData_23 : _GEN_2966; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2968 = 6'h18 == select_46 ? io_inData_24 : _GEN_2967; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2969 = 6'h19 == select_46 ? io_inData_25 : _GEN_2968; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2970 = 6'h1a == select_46 ? io_inData_26 : _GEN_2969; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2971 = 6'h1b == select_46 ? io_inData_27 : _GEN_2970; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2972 = 6'h1c == select_46 ? io_inData_28 : _GEN_2971; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2973 = 6'h1d == select_46 ? io_inData_29 : _GEN_2972; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2974 = 6'h1e == select_46 ? io_inData_30 : _GEN_2973; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2975 = 6'h1f == select_46 ? io_inData_31 : _GEN_2974; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2976 = 6'h20 == select_46 ? io_inData_32 : _GEN_2975; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2977 = 6'h21 == select_46 ? io_inData_33 : _GEN_2976; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2978 = 6'h22 == select_46 ? io_inData_34 : _GEN_2977; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2979 = 6'h23 == select_46 ? io_inData_35 : _GEN_2978; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2980 = 6'h24 == select_46 ? io_inData_36 : _GEN_2979; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2981 = 6'h25 == select_46 ? io_inData_37 : _GEN_2980; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2982 = 6'h26 == select_46 ? io_inData_38 : _GEN_2981; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2983 = 6'h27 == select_46 ? io_inData_39 : _GEN_2982; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2984 = 6'h28 == select_46 ? io_inData_40 : _GEN_2983; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2985 = 6'h29 == select_46 ? io_inData_41 : _GEN_2984; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2986 = 6'h2a == select_46 ? io_inData_42 : _GEN_2985; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2987 = 6'h2b == select_46 ? io_inData_43 : _GEN_2986; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2988 = 6'h2c == select_46 ? io_inData_44 : _GEN_2987; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2989 = 6'h2d == select_46 ? io_inData_45 : _GEN_2988; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2990 = 6'h2e == select_46 ? io_inData_46 : _GEN_2989; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2991 = 6'h2f == select_46 ? io_inData_47 : _GEN_2990; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2992 = 6'h30 == select_46 ? io_inData_48 : _GEN_2991; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2993 = 6'h31 == select_46 ? io_inData_49 : _GEN_2992; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2994 = 6'h32 == select_46 ? io_inData_50 : _GEN_2993; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2995 = 6'h33 == select_46 ? io_inData_51 : _GEN_2994; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2996 = 6'h34 == select_46 ? io_inData_52 : _GEN_2995; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2997 = 6'h35 == select_46 ? io_inData_53 : _GEN_2996; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2998 = 6'h36 == select_46 ? io_inData_54 : _GEN_2997; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_2999 = 6'h37 == select_46 ? io_inData_55 : _GEN_2998; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_3000 = 6'h38 == select_46 ? io_inData_56 : _GEN_2999; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_3001 = 6'h39 == select_46 ? io_inData_57 : _GEN_3000; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_3002 = 6'h3a == select_46 ? io_inData_58 : _GEN_3001; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_3003 = 6'h3b == select_46 ? io_inData_59 : _GEN_3002; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_3004 = 6'h3c == select_46 ? io_inData_60 : _GEN_3003; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_3005 = 6'h3d == select_46 ? io_inData_61 : _GEN_3004; // @[Switch.scala 33:19:@15078.4]
  assign _GEN_3006 = 6'h3e == select_46 ? io_inData_62 : _GEN_3005; // @[Switch.scala 33:19:@15078.4]
  assign _T_35689 = {valid_46_7,valid_46_6,valid_46_5,valid_46_4,valid_46_3,valid_46_2,valid_46_1,valid_46_0}; // @[Switch.scala 34:32:@15085.4]
  assign _T_35697 = {valid_46_15,valid_46_14,valid_46_13,valid_46_12,valid_46_11,valid_46_10,valid_46_9,valid_46_8,_T_35689}; // @[Switch.scala 34:32:@15093.4]
  assign _T_35704 = {valid_46_23,valid_46_22,valid_46_21,valid_46_20,valid_46_19,valid_46_18,valid_46_17,valid_46_16}; // @[Switch.scala 34:32:@15100.4]
  assign _T_35713 = {valid_46_31,valid_46_30,valid_46_29,valid_46_28,valid_46_27,valid_46_26,valid_46_25,valid_46_24,_T_35704,_T_35697}; // @[Switch.scala 34:32:@15109.4]
  assign _T_35720 = {valid_46_39,valid_46_38,valid_46_37,valid_46_36,valid_46_35,valid_46_34,valid_46_33,valid_46_32}; // @[Switch.scala 34:32:@15116.4]
  assign _T_35728 = {valid_46_47,valid_46_46,valid_46_45,valid_46_44,valid_46_43,valid_46_42,valid_46_41,valid_46_40,_T_35720}; // @[Switch.scala 34:32:@15124.4]
  assign _T_35735 = {valid_46_55,valid_46_54,valid_46_53,valid_46_52,valid_46_51,valid_46_50,valid_46_49,valid_46_48}; // @[Switch.scala 34:32:@15131.4]
  assign _T_35744 = {valid_46_63,valid_46_62,valid_46_61,valid_46_60,valid_46_59,valid_46_58,valid_46_57,valid_46_56,_T_35735,_T_35728}; // @[Switch.scala 34:32:@15140.4]
  assign _T_35745 = {_T_35744,_T_35713}; // @[Switch.scala 34:32:@15141.4]
  assign _T_35749 = io_inAddr_0 == 6'h2f; // @[Switch.scala 30:53:@15144.4]
  assign valid_47_0 = io_inValid_0 & _T_35749; // @[Switch.scala 30:36:@15145.4]
  assign _T_35752 = io_inAddr_1 == 6'h2f; // @[Switch.scala 30:53:@15147.4]
  assign valid_47_1 = io_inValid_1 & _T_35752; // @[Switch.scala 30:36:@15148.4]
  assign _T_35755 = io_inAddr_2 == 6'h2f; // @[Switch.scala 30:53:@15150.4]
  assign valid_47_2 = io_inValid_2 & _T_35755; // @[Switch.scala 30:36:@15151.4]
  assign _T_35758 = io_inAddr_3 == 6'h2f; // @[Switch.scala 30:53:@15153.4]
  assign valid_47_3 = io_inValid_3 & _T_35758; // @[Switch.scala 30:36:@15154.4]
  assign _T_35761 = io_inAddr_4 == 6'h2f; // @[Switch.scala 30:53:@15156.4]
  assign valid_47_4 = io_inValid_4 & _T_35761; // @[Switch.scala 30:36:@15157.4]
  assign _T_35764 = io_inAddr_5 == 6'h2f; // @[Switch.scala 30:53:@15159.4]
  assign valid_47_5 = io_inValid_5 & _T_35764; // @[Switch.scala 30:36:@15160.4]
  assign _T_35767 = io_inAddr_6 == 6'h2f; // @[Switch.scala 30:53:@15162.4]
  assign valid_47_6 = io_inValid_6 & _T_35767; // @[Switch.scala 30:36:@15163.4]
  assign _T_35770 = io_inAddr_7 == 6'h2f; // @[Switch.scala 30:53:@15165.4]
  assign valid_47_7 = io_inValid_7 & _T_35770; // @[Switch.scala 30:36:@15166.4]
  assign _T_35773 = io_inAddr_8 == 6'h2f; // @[Switch.scala 30:53:@15168.4]
  assign valid_47_8 = io_inValid_8 & _T_35773; // @[Switch.scala 30:36:@15169.4]
  assign _T_35776 = io_inAddr_9 == 6'h2f; // @[Switch.scala 30:53:@15171.4]
  assign valid_47_9 = io_inValid_9 & _T_35776; // @[Switch.scala 30:36:@15172.4]
  assign _T_35779 = io_inAddr_10 == 6'h2f; // @[Switch.scala 30:53:@15174.4]
  assign valid_47_10 = io_inValid_10 & _T_35779; // @[Switch.scala 30:36:@15175.4]
  assign _T_35782 = io_inAddr_11 == 6'h2f; // @[Switch.scala 30:53:@15177.4]
  assign valid_47_11 = io_inValid_11 & _T_35782; // @[Switch.scala 30:36:@15178.4]
  assign _T_35785 = io_inAddr_12 == 6'h2f; // @[Switch.scala 30:53:@15180.4]
  assign valid_47_12 = io_inValid_12 & _T_35785; // @[Switch.scala 30:36:@15181.4]
  assign _T_35788 = io_inAddr_13 == 6'h2f; // @[Switch.scala 30:53:@15183.4]
  assign valid_47_13 = io_inValid_13 & _T_35788; // @[Switch.scala 30:36:@15184.4]
  assign _T_35791 = io_inAddr_14 == 6'h2f; // @[Switch.scala 30:53:@15186.4]
  assign valid_47_14 = io_inValid_14 & _T_35791; // @[Switch.scala 30:36:@15187.4]
  assign _T_35794 = io_inAddr_15 == 6'h2f; // @[Switch.scala 30:53:@15189.4]
  assign valid_47_15 = io_inValid_15 & _T_35794; // @[Switch.scala 30:36:@15190.4]
  assign _T_35797 = io_inAddr_16 == 6'h2f; // @[Switch.scala 30:53:@15192.4]
  assign valid_47_16 = io_inValid_16 & _T_35797; // @[Switch.scala 30:36:@15193.4]
  assign _T_35800 = io_inAddr_17 == 6'h2f; // @[Switch.scala 30:53:@15195.4]
  assign valid_47_17 = io_inValid_17 & _T_35800; // @[Switch.scala 30:36:@15196.4]
  assign _T_35803 = io_inAddr_18 == 6'h2f; // @[Switch.scala 30:53:@15198.4]
  assign valid_47_18 = io_inValid_18 & _T_35803; // @[Switch.scala 30:36:@15199.4]
  assign _T_35806 = io_inAddr_19 == 6'h2f; // @[Switch.scala 30:53:@15201.4]
  assign valid_47_19 = io_inValid_19 & _T_35806; // @[Switch.scala 30:36:@15202.4]
  assign _T_35809 = io_inAddr_20 == 6'h2f; // @[Switch.scala 30:53:@15204.4]
  assign valid_47_20 = io_inValid_20 & _T_35809; // @[Switch.scala 30:36:@15205.4]
  assign _T_35812 = io_inAddr_21 == 6'h2f; // @[Switch.scala 30:53:@15207.4]
  assign valid_47_21 = io_inValid_21 & _T_35812; // @[Switch.scala 30:36:@15208.4]
  assign _T_35815 = io_inAddr_22 == 6'h2f; // @[Switch.scala 30:53:@15210.4]
  assign valid_47_22 = io_inValid_22 & _T_35815; // @[Switch.scala 30:36:@15211.4]
  assign _T_35818 = io_inAddr_23 == 6'h2f; // @[Switch.scala 30:53:@15213.4]
  assign valid_47_23 = io_inValid_23 & _T_35818; // @[Switch.scala 30:36:@15214.4]
  assign _T_35821 = io_inAddr_24 == 6'h2f; // @[Switch.scala 30:53:@15216.4]
  assign valid_47_24 = io_inValid_24 & _T_35821; // @[Switch.scala 30:36:@15217.4]
  assign _T_35824 = io_inAddr_25 == 6'h2f; // @[Switch.scala 30:53:@15219.4]
  assign valid_47_25 = io_inValid_25 & _T_35824; // @[Switch.scala 30:36:@15220.4]
  assign _T_35827 = io_inAddr_26 == 6'h2f; // @[Switch.scala 30:53:@15222.4]
  assign valid_47_26 = io_inValid_26 & _T_35827; // @[Switch.scala 30:36:@15223.4]
  assign _T_35830 = io_inAddr_27 == 6'h2f; // @[Switch.scala 30:53:@15225.4]
  assign valid_47_27 = io_inValid_27 & _T_35830; // @[Switch.scala 30:36:@15226.4]
  assign _T_35833 = io_inAddr_28 == 6'h2f; // @[Switch.scala 30:53:@15228.4]
  assign valid_47_28 = io_inValid_28 & _T_35833; // @[Switch.scala 30:36:@15229.4]
  assign _T_35836 = io_inAddr_29 == 6'h2f; // @[Switch.scala 30:53:@15231.4]
  assign valid_47_29 = io_inValid_29 & _T_35836; // @[Switch.scala 30:36:@15232.4]
  assign _T_35839 = io_inAddr_30 == 6'h2f; // @[Switch.scala 30:53:@15234.4]
  assign valid_47_30 = io_inValid_30 & _T_35839; // @[Switch.scala 30:36:@15235.4]
  assign _T_35842 = io_inAddr_31 == 6'h2f; // @[Switch.scala 30:53:@15237.4]
  assign valid_47_31 = io_inValid_31 & _T_35842; // @[Switch.scala 30:36:@15238.4]
  assign _T_35845 = io_inAddr_32 == 6'h2f; // @[Switch.scala 30:53:@15240.4]
  assign valid_47_32 = io_inValid_32 & _T_35845; // @[Switch.scala 30:36:@15241.4]
  assign _T_35848 = io_inAddr_33 == 6'h2f; // @[Switch.scala 30:53:@15243.4]
  assign valid_47_33 = io_inValid_33 & _T_35848; // @[Switch.scala 30:36:@15244.4]
  assign _T_35851 = io_inAddr_34 == 6'h2f; // @[Switch.scala 30:53:@15246.4]
  assign valid_47_34 = io_inValid_34 & _T_35851; // @[Switch.scala 30:36:@15247.4]
  assign _T_35854 = io_inAddr_35 == 6'h2f; // @[Switch.scala 30:53:@15249.4]
  assign valid_47_35 = io_inValid_35 & _T_35854; // @[Switch.scala 30:36:@15250.4]
  assign _T_35857 = io_inAddr_36 == 6'h2f; // @[Switch.scala 30:53:@15252.4]
  assign valid_47_36 = io_inValid_36 & _T_35857; // @[Switch.scala 30:36:@15253.4]
  assign _T_35860 = io_inAddr_37 == 6'h2f; // @[Switch.scala 30:53:@15255.4]
  assign valid_47_37 = io_inValid_37 & _T_35860; // @[Switch.scala 30:36:@15256.4]
  assign _T_35863 = io_inAddr_38 == 6'h2f; // @[Switch.scala 30:53:@15258.4]
  assign valid_47_38 = io_inValid_38 & _T_35863; // @[Switch.scala 30:36:@15259.4]
  assign _T_35866 = io_inAddr_39 == 6'h2f; // @[Switch.scala 30:53:@15261.4]
  assign valid_47_39 = io_inValid_39 & _T_35866; // @[Switch.scala 30:36:@15262.4]
  assign _T_35869 = io_inAddr_40 == 6'h2f; // @[Switch.scala 30:53:@15264.4]
  assign valid_47_40 = io_inValid_40 & _T_35869; // @[Switch.scala 30:36:@15265.4]
  assign _T_35872 = io_inAddr_41 == 6'h2f; // @[Switch.scala 30:53:@15267.4]
  assign valid_47_41 = io_inValid_41 & _T_35872; // @[Switch.scala 30:36:@15268.4]
  assign _T_35875 = io_inAddr_42 == 6'h2f; // @[Switch.scala 30:53:@15270.4]
  assign valid_47_42 = io_inValid_42 & _T_35875; // @[Switch.scala 30:36:@15271.4]
  assign _T_35878 = io_inAddr_43 == 6'h2f; // @[Switch.scala 30:53:@15273.4]
  assign valid_47_43 = io_inValid_43 & _T_35878; // @[Switch.scala 30:36:@15274.4]
  assign _T_35881 = io_inAddr_44 == 6'h2f; // @[Switch.scala 30:53:@15276.4]
  assign valid_47_44 = io_inValid_44 & _T_35881; // @[Switch.scala 30:36:@15277.4]
  assign _T_35884 = io_inAddr_45 == 6'h2f; // @[Switch.scala 30:53:@15279.4]
  assign valid_47_45 = io_inValid_45 & _T_35884; // @[Switch.scala 30:36:@15280.4]
  assign _T_35887 = io_inAddr_46 == 6'h2f; // @[Switch.scala 30:53:@15282.4]
  assign valid_47_46 = io_inValid_46 & _T_35887; // @[Switch.scala 30:36:@15283.4]
  assign _T_35890 = io_inAddr_47 == 6'h2f; // @[Switch.scala 30:53:@15285.4]
  assign valid_47_47 = io_inValid_47 & _T_35890; // @[Switch.scala 30:36:@15286.4]
  assign _T_35893 = io_inAddr_48 == 6'h2f; // @[Switch.scala 30:53:@15288.4]
  assign valid_47_48 = io_inValid_48 & _T_35893; // @[Switch.scala 30:36:@15289.4]
  assign _T_35896 = io_inAddr_49 == 6'h2f; // @[Switch.scala 30:53:@15291.4]
  assign valid_47_49 = io_inValid_49 & _T_35896; // @[Switch.scala 30:36:@15292.4]
  assign _T_35899 = io_inAddr_50 == 6'h2f; // @[Switch.scala 30:53:@15294.4]
  assign valid_47_50 = io_inValid_50 & _T_35899; // @[Switch.scala 30:36:@15295.4]
  assign _T_35902 = io_inAddr_51 == 6'h2f; // @[Switch.scala 30:53:@15297.4]
  assign valid_47_51 = io_inValid_51 & _T_35902; // @[Switch.scala 30:36:@15298.4]
  assign _T_35905 = io_inAddr_52 == 6'h2f; // @[Switch.scala 30:53:@15300.4]
  assign valid_47_52 = io_inValid_52 & _T_35905; // @[Switch.scala 30:36:@15301.4]
  assign _T_35908 = io_inAddr_53 == 6'h2f; // @[Switch.scala 30:53:@15303.4]
  assign valid_47_53 = io_inValid_53 & _T_35908; // @[Switch.scala 30:36:@15304.4]
  assign _T_35911 = io_inAddr_54 == 6'h2f; // @[Switch.scala 30:53:@15306.4]
  assign valid_47_54 = io_inValid_54 & _T_35911; // @[Switch.scala 30:36:@15307.4]
  assign _T_35914 = io_inAddr_55 == 6'h2f; // @[Switch.scala 30:53:@15309.4]
  assign valid_47_55 = io_inValid_55 & _T_35914; // @[Switch.scala 30:36:@15310.4]
  assign _T_35917 = io_inAddr_56 == 6'h2f; // @[Switch.scala 30:53:@15312.4]
  assign valid_47_56 = io_inValid_56 & _T_35917; // @[Switch.scala 30:36:@15313.4]
  assign _T_35920 = io_inAddr_57 == 6'h2f; // @[Switch.scala 30:53:@15315.4]
  assign valid_47_57 = io_inValid_57 & _T_35920; // @[Switch.scala 30:36:@15316.4]
  assign _T_35923 = io_inAddr_58 == 6'h2f; // @[Switch.scala 30:53:@15318.4]
  assign valid_47_58 = io_inValid_58 & _T_35923; // @[Switch.scala 30:36:@15319.4]
  assign _T_35926 = io_inAddr_59 == 6'h2f; // @[Switch.scala 30:53:@15321.4]
  assign valid_47_59 = io_inValid_59 & _T_35926; // @[Switch.scala 30:36:@15322.4]
  assign _T_35929 = io_inAddr_60 == 6'h2f; // @[Switch.scala 30:53:@15324.4]
  assign valid_47_60 = io_inValid_60 & _T_35929; // @[Switch.scala 30:36:@15325.4]
  assign _T_35932 = io_inAddr_61 == 6'h2f; // @[Switch.scala 30:53:@15327.4]
  assign valid_47_61 = io_inValid_61 & _T_35932; // @[Switch.scala 30:36:@15328.4]
  assign _T_35935 = io_inAddr_62 == 6'h2f; // @[Switch.scala 30:53:@15330.4]
  assign valid_47_62 = io_inValid_62 & _T_35935; // @[Switch.scala 30:36:@15331.4]
  assign _T_35938 = io_inAddr_63 == 6'h2f; // @[Switch.scala 30:53:@15333.4]
  assign valid_47_63 = io_inValid_63 & _T_35938; // @[Switch.scala 30:36:@15334.4]
  assign _T_36004 = valid_47_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@15336.4]
  assign _T_36005 = valid_47_61 ? 6'h3d : _T_36004; // @[Mux.scala 31:69:@15337.4]
  assign _T_36006 = valid_47_60 ? 6'h3c : _T_36005; // @[Mux.scala 31:69:@15338.4]
  assign _T_36007 = valid_47_59 ? 6'h3b : _T_36006; // @[Mux.scala 31:69:@15339.4]
  assign _T_36008 = valid_47_58 ? 6'h3a : _T_36007; // @[Mux.scala 31:69:@15340.4]
  assign _T_36009 = valid_47_57 ? 6'h39 : _T_36008; // @[Mux.scala 31:69:@15341.4]
  assign _T_36010 = valid_47_56 ? 6'h38 : _T_36009; // @[Mux.scala 31:69:@15342.4]
  assign _T_36011 = valid_47_55 ? 6'h37 : _T_36010; // @[Mux.scala 31:69:@15343.4]
  assign _T_36012 = valid_47_54 ? 6'h36 : _T_36011; // @[Mux.scala 31:69:@15344.4]
  assign _T_36013 = valid_47_53 ? 6'h35 : _T_36012; // @[Mux.scala 31:69:@15345.4]
  assign _T_36014 = valid_47_52 ? 6'h34 : _T_36013; // @[Mux.scala 31:69:@15346.4]
  assign _T_36015 = valid_47_51 ? 6'h33 : _T_36014; // @[Mux.scala 31:69:@15347.4]
  assign _T_36016 = valid_47_50 ? 6'h32 : _T_36015; // @[Mux.scala 31:69:@15348.4]
  assign _T_36017 = valid_47_49 ? 6'h31 : _T_36016; // @[Mux.scala 31:69:@15349.4]
  assign _T_36018 = valid_47_48 ? 6'h30 : _T_36017; // @[Mux.scala 31:69:@15350.4]
  assign _T_36019 = valid_47_47 ? 6'h2f : _T_36018; // @[Mux.scala 31:69:@15351.4]
  assign _T_36020 = valid_47_46 ? 6'h2e : _T_36019; // @[Mux.scala 31:69:@15352.4]
  assign _T_36021 = valid_47_45 ? 6'h2d : _T_36020; // @[Mux.scala 31:69:@15353.4]
  assign _T_36022 = valid_47_44 ? 6'h2c : _T_36021; // @[Mux.scala 31:69:@15354.4]
  assign _T_36023 = valid_47_43 ? 6'h2b : _T_36022; // @[Mux.scala 31:69:@15355.4]
  assign _T_36024 = valid_47_42 ? 6'h2a : _T_36023; // @[Mux.scala 31:69:@15356.4]
  assign _T_36025 = valid_47_41 ? 6'h29 : _T_36024; // @[Mux.scala 31:69:@15357.4]
  assign _T_36026 = valid_47_40 ? 6'h28 : _T_36025; // @[Mux.scala 31:69:@15358.4]
  assign _T_36027 = valid_47_39 ? 6'h27 : _T_36026; // @[Mux.scala 31:69:@15359.4]
  assign _T_36028 = valid_47_38 ? 6'h26 : _T_36027; // @[Mux.scala 31:69:@15360.4]
  assign _T_36029 = valid_47_37 ? 6'h25 : _T_36028; // @[Mux.scala 31:69:@15361.4]
  assign _T_36030 = valid_47_36 ? 6'h24 : _T_36029; // @[Mux.scala 31:69:@15362.4]
  assign _T_36031 = valid_47_35 ? 6'h23 : _T_36030; // @[Mux.scala 31:69:@15363.4]
  assign _T_36032 = valid_47_34 ? 6'h22 : _T_36031; // @[Mux.scala 31:69:@15364.4]
  assign _T_36033 = valid_47_33 ? 6'h21 : _T_36032; // @[Mux.scala 31:69:@15365.4]
  assign _T_36034 = valid_47_32 ? 6'h20 : _T_36033; // @[Mux.scala 31:69:@15366.4]
  assign _T_36035 = valid_47_31 ? 6'h1f : _T_36034; // @[Mux.scala 31:69:@15367.4]
  assign _T_36036 = valid_47_30 ? 6'h1e : _T_36035; // @[Mux.scala 31:69:@15368.4]
  assign _T_36037 = valid_47_29 ? 6'h1d : _T_36036; // @[Mux.scala 31:69:@15369.4]
  assign _T_36038 = valid_47_28 ? 6'h1c : _T_36037; // @[Mux.scala 31:69:@15370.4]
  assign _T_36039 = valid_47_27 ? 6'h1b : _T_36038; // @[Mux.scala 31:69:@15371.4]
  assign _T_36040 = valid_47_26 ? 6'h1a : _T_36039; // @[Mux.scala 31:69:@15372.4]
  assign _T_36041 = valid_47_25 ? 6'h19 : _T_36040; // @[Mux.scala 31:69:@15373.4]
  assign _T_36042 = valid_47_24 ? 6'h18 : _T_36041; // @[Mux.scala 31:69:@15374.4]
  assign _T_36043 = valid_47_23 ? 6'h17 : _T_36042; // @[Mux.scala 31:69:@15375.4]
  assign _T_36044 = valid_47_22 ? 6'h16 : _T_36043; // @[Mux.scala 31:69:@15376.4]
  assign _T_36045 = valid_47_21 ? 6'h15 : _T_36044; // @[Mux.scala 31:69:@15377.4]
  assign _T_36046 = valid_47_20 ? 6'h14 : _T_36045; // @[Mux.scala 31:69:@15378.4]
  assign _T_36047 = valid_47_19 ? 6'h13 : _T_36046; // @[Mux.scala 31:69:@15379.4]
  assign _T_36048 = valid_47_18 ? 6'h12 : _T_36047; // @[Mux.scala 31:69:@15380.4]
  assign _T_36049 = valid_47_17 ? 6'h11 : _T_36048; // @[Mux.scala 31:69:@15381.4]
  assign _T_36050 = valid_47_16 ? 6'h10 : _T_36049; // @[Mux.scala 31:69:@15382.4]
  assign _T_36051 = valid_47_15 ? 6'hf : _T_36050; // @[Mux.scala 31:69:@15383.4]
  assign _T_36052 = valid_47_14 ? 6'he : _T_36051; // @[Mux.scala 31:69:@15384.4]
  assign _T_36053 = valid_47_13 ? 6'hd : _T_36052; // @[Mux.scala 31:69:@15385.4]
  assign _T_36054 = valid_47_12 ? 6'hc : _T_36053; // @[Mux.scala 31:69:@15386.4]
  assign _T_36055 = valid_47_11 ? 6'hb : _T_36054; // @[Mux.scala 31:69:@15387.4]
  assign _T_36056 = valid_47_10 ? 6'ha : _T_36055; // @[Mux.scala 31:69:@15388.4]
  assign _T_36057 = valid_47_9 ? 6'h9 : _T_36056; // @[Mux.scala 31:69:@15389.4]
  assign _T_36058 = valid_47_8 ? 6'h8 : _T_36057; // @[Mux.scala 31:69:@15390.4]
  assign _T_36059 = valid_47_7 ? 6'h7 : _T_36058; // @[Mux.scala 31:69:@15391.4]
  assign _T_36060 = valid_47_6 ? 6'h6 : _T_36059; // @[Mux.scala 31:69:@15392.4]
  assign _T_36061 = valid_47_5 ? 6'h5 : _T_36060; // @[Mux.scala 31:69:@15393.4]
  assign _T_36062 = valid_47_4 ? 6'h4 : _T_36061; // @[Mux.scala 31:69:@15394.4]
  assign _T_36063 = valid_47_3 ? 6'h3 : _T_36062; // @[Mux.scala 31:69:@15395.4]
  assign _T_36064 = valid_47_2 ? 6'h2 : _T_36063; // @[Mux.scala 31:69:@15396.4]
  assign _T_36065 = valid_47_1 ? 6'h1 : _T_36064; // @[Mux.scala 31:69:@15397.4]
  assign select_47 = valid_47_0 ? 6'h0 : _T_36065; // @[Mux.scala 31:69:@15398.4]
  assign _GEN_3009 = 6'h1 == select_47 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3010 = 6'h2 == select_47 ? io_inData_2 : _GEN_3009; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3011 = 6'h3 == select_47 ? io_inData_3 : _GEN_3010; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3012 = 6'h4 == select_47 ? io_inData_4 : _GEN_3011; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3013 = 6'h5 == select_47 ? io_inData_5 : _GEN_3012; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3014 = 6'h6 == select_47 ? io_inData_6 : _GEN_3013; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3015 = 6'h7 == select_47 ? io_inData_7 : _GEN_3014; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3016 = 6'h8 == select_47 ? io_inData_8 : _GEN_3015; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3017 = 6'h9 == select_47 ? io_inData_9 : _GEN_3016; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3018 = 6'ha == select_47 ? io_inData_10 : _GEN_3017; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3019 = 6'hb == select_47 ? io_inData_11 : _GEN_3018; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3020 = 6'hc == select_47 ? io_inData_12 : _GEN_3019; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3021 = 6'hd == select_47 ? io_inData_13 : _GEN_3020; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3022 = 6'he == select_47 ? io_inData_14 : _GEN_3021; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3023 = 6'hf == select_47 ? io_inData_15 : _GEN_3022; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3024 = 6'h10 == select_47 ? io_inData_16 : _GEN_3023; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3025 = 6'h11 == select_47 ? io_inData_17 : _GEN_3024; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3026 = 6'h12 == select_47 ? io_inData_18 : _GEN_3025; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3027 = 6'h13 == select_47 ? io_inData_19 : _GEN_3026; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3028 = 6'h14 == select_47 ? io_inData_20 : _GEN_3027; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3029 = 6'h15 == select_47 ? io_inData_21 : _GEN_3028; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3030 = 6'h16 == select_47 ? io_inData_22 : _GEN_3029; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3031 = 6'h17 == select_47 ? io_inData_23 : _GEN_3030; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3032 = 6'h18 == select_47 ? io_inData_24 : _GEN_3031; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3033 = 6'h19 == select_47 ? io_inData_25 : _GEN_3032; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3034 = 6'h1a == select_47 ? io_inData_26 : _GEN_3033; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3035 = 6'h1b == select_47 ? io_inData_27 : _GEN_3034; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3036 = 6'h1c == select_47 ? io_inData_28 : _GEN_3035; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3037 = 6'h1d == select_47 ? io_inData_29 : _GEN_3036; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3038 = 6'h1e == select_47 ? io_inData_30 : _GEN_3037; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3039 = 6'h1f == select_47 ? io_inData_31 : _GEN_3038; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3040 = 6'h20 == select_47 ? io_inData_32 : _GEN_3039; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3041 = 6'h21 == select_47 ? io_inData_33 : _GEN_3040; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3042 = 6'h22 == select_47 ? io_inData_34 : _GEN_3041; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3043 = 6'h23 == select_47 ? io_inData_35 : _GEN_3042; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3044 = 6'h24 == select_47 ? io_inData_36 : _GEN_3043; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3045 = 6'h25 == select_47 ? io_inData_37 : _GEN_3044; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3046 = 6'h26 == select_47 ? io_inData_38 : _GEN_3045; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3047 = 6'h27 == select_47 ? io_inData_39 : _GEN_3046; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3048 = 6'h28 == select_47 ? io_inData_40 : _GEN_3047; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3049 = 6'h29 == select_47 ? io_inData_41 : _GEN_3048; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3050 = 6'h2a == select_47 ? io_inData_42 : _GEN_3049; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3051 = 6'h2b == select_47 ? io_inData_43 : _GEN_3050; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3052 = 6'h2c == select_47 ? io_inData_44 : _GEN_3051; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3053 = 6'h2d == select_47 ? io_inData_45 : _GEN_3052; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3054 = 6'h2e == select_47 ? io_inData_46 : _GEN_3053; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3055 = 6'h2f == select_47 ? io_inData_47 : _GEN_3054; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3056 = 6'h30 == select_47 ? io_inData_48 : _GEN_3055; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3057 = 6'h31 == select_47 ? io_inData_49 : _GEN_3056; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3058 = 6'h32 == select_47 ? io_inData_50 : _GEN_3057; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3059 = 6'h33 == select_47 ? io_inData_51 : _GEN_3058; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3060 = 6'h34 == select_47 ? io_inData_52 : _GEN_3059; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3061 = 6'h35 == select_47 ? io_inData_53 : _GEN_3060; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3062 = 6'h36 == select_47 ? io_inData_54 : _GEN_3061; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3063 = 6'h37 == select_47 ? io_inData_55 : _GEN_3062; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3064 = 6'h38 == select_47 ? io_inData_56 : _GEN_3063; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3065 = 6'h39 == select_47 ? io_inData_57 : _GEN_3064; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3066 = 6'h3a == select_47 ? io_inData_58 : _GEN_3065; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3067 = 6'h3b == select_47 ? io_inData_59 : _GEN_3066; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3068 = 6'h3c == select_47 ? io_inData_60 : _GEN_3067; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3069 = 6'h3d == select_47 ? io_inData_61 : _GEN_3068; // @[Switch.scala 33:19:@15400.4]
  assign _GEN_3070 = 6'h3e == select_47 ? io_inData_62 : _GEN_3069; // @[Switch.scala 33:19:@15400.4]
  assign _T_36074 = {valid_47_7,valid_47_6,valid_47_5,valid_47_4,valid_47_3,valid_47_2,valid_47_1,valid_47_0}; // @[Switch.scala 34:32:@15407.4]
  assign _T_36082 = {valid_47_15,valid_47_14,valid_47_13,valid_47_12,valid_47_11,valid_47_10,valid_47_9,valid_47_8,_T_36074}; // @[Switch.scala 34:32:@15415.4]
  assign _T_36089 = {valid_47_23,valid_47_22,valid_47_21,valid_47_20,valid_47_19,valid_47_18,valid_47_17,valid_47_16}; // @[Switch.scala 34:32:@15422.4]
  assign _T_36098 = {valid_47_31,valid_47_30,valid_47_29,valid_47_28,valid_47_27,valid_47_26,valid_47_25,valid_47_24,_T_36089,_T_36082}; // @[Switch.scala 34:32:@15431.4]
  assign _T_36105 = {valid_47_39,valid_47_38,valid_47_37,valid_47_36,valid_47_35,valid_47_34,valid_47_33,valid_47_32}; // @[Switch.scala 34:32:@15438.4]
  assign _T_36113 = {valid_47_47,valid_47_46,valid_47_45,valid_47_44,valid_47_43,valid_47_42,valid_47_41,valid_47_40,_T_36105}; // @[Switch.scala 34:32:@15446.4]
  assign _T_36120 = {valid_47_55,valid_47_54,valid_47_53,valid_47_52,valid_47_51,valid_47_50,valid_47_49,valid_47_48}; // @[Switch.scala 34:32:@15453.4]
  assign _T_36129 = {valid_47_63,valid_47_62,valid_47_61,valid_47_60,valid_47_59,valid_47_58,valid_47_57,valid_47_56,_T_36120,_T_36113}; // @[Switch.scala 34:32:@15462.4]
  assign _T_36130 = {_T_36129,_T_36098}; // @[Switch.scala 34:32:@15463.4]
  assign _T_36134 = io_inAddr_0 == 6'h30; // @[Switch.scala 30:53:@15466.4]
  assign valid_48_0 = io_inValid_0 & _T_36134; // @[Switch.scala 30:36:@15467.4]
  assign _T_36137 = io_inAddr_1 == 6'h30; // @[Switch.scala 30:53:@15469.4]
  assign valid_48_1 = io_inValid_1 & _T_36137; // @[Switch.scala 30:36:@15470.4]
  assign _T_36140 = io_inAddr_2 == 6'h30; // @[Switch.scala 30:53:@15472.4]
  assign valid_48_2 = io_inValid_2 & _T_36140; // @[Switch.scala 30:36:@15473.4]
  assign _T_36143 = io_inAddr_3 == 6'h30; // @[Switch.scala 30:53:@15475.4]
  assign valid_48_3 = io_inValid_3 & _T_36143; // @[Switch.scala 30:36:@15476.4]
  assign _T_36146 = io_inAddr_4 == 6'h30; // @[Switch.scala 30:53:@15478.4]
  assign valid_48_4 = io_inValid_4 & _T_36146; // @[Switch.scala 30:36:@15479.4]
  assign _T_36149 = io_inAddr_5 == 6'h30; // @[Switch.scala 30:53:@15481.4]
  assign valid_48_5 = io_inValid_5 & _T_36149; // @[Switch.scala 30:36:@15482.4]
  assign _T_36152 = io_inAddr_6 == 6'h30; // @[Switch.scala 30:53:@15484.4]
  assign valid_48_6 = io_inValid_6 & _T_36152; // @[Switch.scala 30:36:@15485.4]
  assign _T_36155 = io_inAddr_7 == 6'h30; // @[Switch.scala 30:53:@15487.4]
  assign valid_48_7 = io_inValid_7 & _T_36155; // @[Switch.scala 30:36:@15488.4]
  assign _T_36158 = io_inAddr_8 == 6'h30; // @[Switch.scala 30:53:@15490.4]
  assign valid_48_8 = io_inValid_8 & _T_36158; // @[Switch.scala 30:36:@15491.4]
  assign _T_36161 = io_inAddr_9 == 6'h30; // @[Switch.scala 30:53:@15493.4]
  assign valid_48_9 = io_inValid_9 & _T_36161; // @[Switch.scala 30:36:@15494.4]
  assign _T_36164 = io_inAddr_10 == 6'h30; // @[Switch.scala 30:53:@15496.4]
  assign valid_48_10 = io_inValid_10 & _T_36164; // @[Switch.scala 30:36:@15497.4]
  assign _T_36167 = io_inAddr_11 == 6'h30; // @[Switch.scala 30:53:@15499.4]
  assign valid_48_11 = io_inValid_11 & _T_36167; // @[Switch.scala 30:36:@15500.4]
  assign _T_36170 = io_inAddr_12 == 6'h30; // @[Switch.scala 30:53:@15502.4]
  assign valid_48_12 = io_inValid_12 & _T_36170; // @[Switch.scala 30:36:@15503.4]
  assign _T_36173 = io_inAddr_13 == 6'h30; // @[Switch.scala 30:53:@15505.4]
  assign valid_48_13 = io_inValid_13 & _T_36173; // @[Switch.scala 30:36:@15506.4]
  assign _T_36176 = io_inAddr_14 == 6'h30; // @[Switch.scala 30:53:@15508.4]
  assign valid_48_14 = io_inValid_14 & _T_36176; // @[Switch.scala 30:36:@15509.4]
  assign _T_36179 = io_inAddr_15 == 6'h30; // @[Switch.scala 30:53:@15511.4]
  assign valid_48_15 = io_inValid_15 & _T_36179; // @[Switch.scala 30:36:@15512.4]
  assign _T_36182 = io_inAddr_16 == 6'h30; // @[Switch.scala 30:53:@15514.4]
  assign valid_48_16 = io_inValid_16 & _T_36182; // @[Switch.scala 30:36:@15515.4]
  assign _T_36185 = io_inAddr_17 == 6'h30; // @[Switch.scala 30:53:@15517.4]
  assign valid_48_17 = io_inValid_17 & _T_36185; // @[Switch.scala 30:36:@15518.4]
  assign _T_36188 = io_inAddr_18 == 6'h30; // @[Switch.scala 30:53:@15520.4]
  assign valid_48_18 = io_inValid_18 & _T_36188; // @[Switch.scala 30:36:@15521.4]
  assign _T_36191 = io_inAddr_19 == 6'h30; // @[Switch.scala 30:53:@15523.4]
  assign valid_48_19 = io_inValid_19 & _T_36191; // @[Switch.scala 30:36:@15524.4]
  assign _T_36194 = io_inAddr_20 == 6'h30; // @[Switch.scala 30:53:@15526.4]
  assign valid_48_20 = io_inValid_20 & _T_36194; // @[Switch.scala 30:36:@15527.4]
  assign _T_36197 = io_inAddr_21 == 6'h30; // @[Switch.scala 30:53:@15529.4]
  assign valid_48_21 = io_inValid_21 & _T_36197; // @[Switch.scala 30:36:@15530.4]
  assign _T_36200 = io_inAddr_22 == 6'h30; // @[Switch.scala 30:53:@15532.4]
  assign valid_48_22 = io_inValid_22 & _T_36200; // @[Switch.scala 30:36:@15533.4]
  assign _T_36203 = io_inAddr_23 == 6'h30; // @[Switch.scala 30:53:@15535.4]
  assign valid_48_23 = io_inValid_23 & _T_36203; // @[Switch.scala 30:36:@15536.4]
  assign _T_36206 = io_inAddr_24 == 6'h30; // @[Switch.scala 30:53:@15538.4]
  assign valid_48_24 = io_inValid_24 & _T_36206; // @[Switch.scala 30:36:@15539.4]
  assign _T_36209 = io_inAddr_25 == 6'h30; // @[Switch.scala 30:53:@15541.4]
  assign valid_48_25 = io_inValid_25 & _T_36209; // @[Switch.scala 30:36:@15542.4]
  assign _T_36212 = io_inAddr_26 == 6'h30; // @[Switch.scala 30:53:@15544.4]
  assign valid_48_26 = io_inValid_26 & _T_36212; // @[Switch.scala 30:36:@15545.4]
  assign _T_36215 = io_inAddr_27 == 6'h30; // @[Switch.scala 30:53:@15547.4]
  assign valid_48_27 = io_inValid_27 & _T_36215; // @[Switch.scala 30:36:@15548.4]
  assign _T_36218 = io_inAddr_28 == 6'h30; // @[Switch.scala 30:53:@15550.4]
  assign valid_48_28 = io_inValid_28 & _T_36218; // @[Switch.scala 30:36:@15551.4]
  assign _T_36221 = io_inAddr_29 == 6'h30; // @[Switch.scala 30:53:@15553.4]
  assign valid_48_29 = io_inValid_29 & _T_36221; // @[Switch.scala 30:36:@15554.4]
  assign _T_36224 = io_inAddr_30 == 6'h30; // @[Switch.scala 30:53:@15556.4]
  assign valid_48_30 = io_inValid_30 & _T_36224; // @[Switch.scala 30:36:@15557.4]
  assign _T_36227 = io_inAddr_31 == 6'h30; // @[Switch.scala 30:53:@15559.4]
  assign valid_48_31 = io_inValid_31 & _T_36227; // @[Switch.scala 30:36:@15560.4]
  assign _T_36230 = io_inAddr_32 == 6'h30; // @[Switch.scala 30:53:@15562.4]
  assign valid_48_32 = io_inValid_32 & _T_36230; // @[Switch.scala 30:36:@15563.4]
  assign _T_36233 = io_inAddr_33 == 6'h30; // @[Switch.scala 30:53:@15565.4]
  assign valid_48_33 = io_inValid_33 & _T_36233; // @[Switch.scala 30:36:@15566.4]
  assign _T_36236 = io_inAddr_34 == 6'h30; // @[Switch.scala 30:53:@15568.4]
  assign valid_48_34 = io_inValid_34 & _T_36236; // @[Switch.scala 30:36:@15569.4]
  assign _T_36239 = io_inAddr_35 == 6'h30; // @[Switch.scala 30:53:@15571.4]
  assign valid_48_35 = io_inValid_35 & _T_36239; // @[Switch.scala 30:36:@15572.4]
  assign _T_36242 = io_inAddr_36 == 6'h30; // @[Switch.scala 30:53:@15574.4]
  assign valid_48_36 = io_inValid_36 & _T_36242; // @[Switch.scala 30:36:@15575.4]
  assign _T_36245 = io_inAddr_37 == 6'h30; // @[Switch.scala 30:53:@15577.4]
  assign valid_48_37 = io_inValid_37 & _T_36245; // @[Switch.scala 30:36:@15578.4]
  assign _T_36248 = io_inAddr_38 == 6'h30; // @[Switch.scala 30:53:@15580.4]
  assign valid_48_38 = io_inValid_38 & _T_36248; // @[Switch.scala 30:36:@15581.4]
  assign _T_36251 = io_inAddr_39 == 6'h30; // @[Switch.scala 30:53:@15583.4]
  assign valid_48_39 = io_inValid_39 & _T_36251; // @[Switch.scala 30:36:@15584.4]
  assign _T_36254 = io_inAddr_40 == 6'h30; // @[Switch.scala 30:53:@15586.4]
  assign valid_48_40 = io_inValid_40 & _T_36254; // @[Switch.scala 30:36:@15587.4]
  assign _T_36257 = io_inAddr_41 == 6'h30; // @[Switch.scala 30:53:@15589.4]
  assign valid_48_41 = io_inValid_41 & _T_36257; // @[Switch.scala 30:36:@15590.4]
  assign _T_36260 = io_inAddr_42 == 6'h30; // @[Switch.scala 30:53:@15592.4]
  assign valid_48_42 = io_inValid_42 & _T_36260; // @[Switch.scala 30:36:@15593.4]
  assign _T_36263 = io_inAddr_43 == 6'h30; // @[Switch.scala 30:53:@15595.4]
  assign valid_48_43 = io_inValid_43 & _T_36263; // @[Switch.scala 30:36:@15596.4]
  assign _T_36266 = io_inAddr_44 == 6'h30; // @[Switch.scala 30:53:@15598.4]
  assign valid_48_44 = io_inValid_44 & _T_36266; // @[Switch.scala 30:36:@15599.4]
  assign _T_36269 = io_inAddr_45 == 6'h30; // @[Switch.scala 30:53:@15601.4]
  assign valid_48_45 = io_inValid_45 & _T_36269; // @[Switch.scala 30:36:@15602.4]
  assign _T_36272 = io_inAddr_46 == 6'h30; // @[Switch.scala 30:53:@15604.4]
  assign valid_48_46 = io_inValid_46 & _T_36272; // @[Switch.scala 30:36:@15605.4]
  assign _T_36275 = io_inAddr_47 == 6'h30; // @[Switch.scala 30:53:@15607.4]
  assign valid_48_47 = io_inValid_47 & _T_36275; // @[Switch.scala 30:36:@15608.4]
  assign _T_36278 = io_inAddr_48 == 6'h30; // @[Switch.scala 30:53:@15610.4]
  assign valid_48_48 = io_inValid_48 & _T_36278; // @[Switch.scala 30:36:@15611.4]
  assign _T_36281 = io_inAddr_49 == 6'h30; // @[Switch.scala 30:53:@15613.4]
  assign valid_48_49 = io_inValid_49 & _T_36281; // @[Switch.scala 30:36:@15614.4]
  assign _T_36284 = io_inAddr_50 == 6'h30; // @[Switch.scala 30:53:@15616.4]
  assign valid_48_50 = io_inValid_50 & _T_36284; // @[Switch.scala 30:36:@15617.4]
  assign _T_36287 = io_inAddr_51 == 6'h30; // @[Switch.scala 30:53:@15619.4]
  assign valid_48_51 = io_inValid_51 & _T_36287; // @[Switch.scala 30:36:@15620.4]
  assign _T_36290 = io_inAddr_52 == 6'h30; // @[Switch.scala 30:53:@15622.4]
  assign valid_48_52 = io_inValid_52 & _T_36290; // @[Switch.scala 30:36:@15623.4]
  assign _T_36293 = io_inAddr_53 == 6'h30; // @[Switch.scala 30:53:@15625.4]
  assign valid_48_53 = io_inValid_53 & _T_36293; // @[Switch.scala 30:36:@15626.4]
  assign _T_36296 = io_inAddr_54 == 6'h30; // @[Switch.scala 30:53:@15628.4]
  assign valid_48_54 = io_inValid_54 & _T_36296; // @[Switch.scala 30:36:@15629.4]
  assign _T_36299 = io_inAddr_55 == 6'h30; // @[Switch.scala 30:53:@15631.4]
  assign valid_48_55 = io_inValid_55 & _T_36299; // @[Switch.scala 30:36:@15632.4]
  assign _T_36302 = io_inAddr_56 == 6'h30; // @[Switch.scala 30:53:@15634.4]
  assign valid_48_56 = io_inValid_56 & _T_36302; // @[Switch.scala 30:36:@15635.4]
  assign _T_36305 = io_inAddr_57 == 6'h30; // @[Switch.scala 30:53:@15637.4]
  assign valid_48_57 = io_inValid_57 & _T_36305; // @[Switch.scala 30:36:@15638.4]
  assign _T_36308 = io_inAddr_58 == 6'h30; // @[Switch.scala 30:53:@15640.4]
  assign valid_48_58 = io_inValid_58 & _T_36308; // @[Switch.scala 30:36:@15641.4]
  assign _T_36311 = io_inAddr_59 == 6'h30; // @[Switch.scala 30:53:@15643.4]
  assign valid_48_59 = io_inValid_59 & _T_36311; // @[Switch.scala 30:36:@15644.4]
  assign _T_36314 = io_inAddr_60 == 6'h30; // @[Switch.scala 30:53:@15646.4]
  assign valid_48_60 = io_inValid_60 & _T_36314; // @[Switch.scala 30:36:@15647.4]
  assign _T_36317 = io_inAddr_61 == 6'h30; // @[Switch.scala 30:53:@15649.4]
  assign valid_48_61 = io_inValid_61 & _T_36317; // @[Switch.scala 30:36:@15650.4]
  assign _T_36320 = io_inAddr_62 == 6'h30; // @[Switch.scala 30:53:@15652.4]
  assign valid_48_62 = io_inValid_62 & _T_36320; // @[Switch.scala 30:36:@15653.4]
  assign _T_36323 = io_inAddr_63 == 6'h30; // @[Switch.scala 30:53:@15655.4]
  assign valid_48_63 = io_inValid_63 & _T_36323; // @[Switch.scala 30:36:@15656.4]
  assign _T_36389 = valid_48_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@15658.4]
  assign _T_36390 = valid_48_61 ? 6'h3d : _T_36389; // @[Mux.scala 31:69:@15659.4]
  assign _T_36391 = valid_48_60 ? 6'h3c : _T_36390; // @[Mux.scala 31:69:@15660.4]
  assign _T_36392 = valid_48_59 ? 6'h3b : _T_36391; // @[Mux.scala 31:69:@15661.4]
  assign _T_36393 = valid_48_58 ? 6'h3a : _T_36392; // @[Mux.scala 31:69:@15662.4]
  assign _T_36394 = valid_48_57 ? 6'h39 : _T_36393; // @[Mux.scala 31:69:@15663.4]
  assign _T_36395 = valid_48_56 ? 6'h38 : _T_36394; // @[Mux.scala 31:69:@15664.4]
  assign _T_36396 = valid_48_55 ? 6'h37 : _T_36395; // @[Mux.scala 31:69:@15665.4]
  assign _T_36397 = valid_48_54 ? 6'h36 : _T_36396; // @[Mux.scala 31:69:@15666.4]
  assign _T_36398 = valid_48_53 ? 6'h35 : _T_36397; // @[Mux.scala 31:69:@15667.4]
  assign _T_36399 = valid_48_52 ? 6'h34 : _T_36398; // @[Mux.scala 31:69:@15668.4]
  assign _T_36400 = valid_48_51 ? 6'h33 : _T_36399; // @[Mux.scala 31:69:@15669.4]
  assign _T_36401 = valid_48_50 ? 6'h32 : _T_36400; // @[Mux.scala 31:69:@15670.4]
  assign _T_36402 = valid_48_49 ? 6'h31 : _T_36401; // @[Mux.scala 31:69:@15671.4]
  assign _T_36403 = valid_48_48 ? 6'h30 : _T_36402; // @[Mux.scala 31:69:@15672.4]
  assign _T_36404 = valid_48_47 ? 6'h2f : _T_36403; // @[Mux.scala 31:69:@15673.4]
  assign _T_36405 = valid_48_46 ? 6'h2e : _T_36404; // @[Mux.scala 31:69:@15674.4]
  assign _T_36406 = valid_48_45 ? 6'h2d : _T_36405; // @[Mux.scala 31:69:@15675.4]
  assign _T_36407 = valid_48_44 ? 6'h2c : _T_36406; // @[Mux.scala 31:69:@15676.4]
  assign _T_36408 = valid_48_43 ? 6'h2b : _T_36407; // @[Mux.scala 31:69:@15677.4]
  assign _T_36409 = valid_48_42 ? 6'h2a : _T_36408; // @[Mux.scala 31:69:@15678.4]
  assign _T_36410 = valid_48_41 ? 6'h29 : _T_36409; // @[Mux.scala 31:69:@15679.4]
  assign _T_36411 = valid_48_40 ? 6'h28 : _T_36410; // @[Mux.scala 31:69:@15680.4]
  assign _T_36412 = valid_48_39 ? 6'h27 : _T_36411; // @[Mux.scala 31:69:@15681.4]
  assign _T_36413 = valid_48_38 ? 6'h26 : _T_36412; // @[Mux.scala 31:69:@15682.4]
  assign _T_36414 = valid_48_37 ? 6'h25 : _T_36413; // @[Mux.scala 31:69:@15683.4]
  assign _T_36415 = valid_48_36 ? 6'h24 : _T_36414; // @[Mux.scala 31:69:@15684.4]
  assign _T_36416 = valid_48_35 ? 6'h23 : _T_36415; // @[Mux.scala 31:69:@15685.4]
  assign _T_36417 = valid_48_34 ? 6'h22 : _T_36416; // @[Mux.scala 31:69:@15686.4]
  assign _T_36418 = valid_48_33 ? 6'h21 : _T_36417; // @[Mux.scala 31:69:@15687.4]
  assign _T_36419 = valid_48_32 ? 6'h20 : _T_36418; // @[Mux.scala 31:69:@15688.4]
  assign _T_36420 = valid_48_31 ? 6'h1f : _T_36419; // @[Mux.scala 31:69:@15689.4]
  assign _T_36421 = valid_48_30 ? 6'h1e : _T_36420; // @[Mux.scala 31:69:@15690.4]
  assign _T_36422 = valid_48_29 ? 6'h1d : _T_36421; // @[Mux.scala 31:69:@15691.4]
  assign _T_36423 = valid_48_28 ? 6'h1c : _T_36422; // @[Mux.scala 31:69:@15692.4]
  assign _T_36424 = valid_48_27 ? 6'h1b : _T_36423; // @[Mux.scala 31:69:@15693.4]
  assign _T_36425 = valid_48_26 ? 6'h1a : _T_36424; // @[Mux.scala 31:69:@15694.4]
  assign _T_36426 = valid_48_25 ? 6'h19 : _T_36425; // @[Mux.scala 31:69:@15695.4]
  assign _T_36427 = valid_48_24 ? 6'h18 : _T_36426; // @[Mux.scala 31:69:@15696.4]
  assign _T_36428 = valid_48_23 ? 6'h17 : _T_36427; // @[Mux.scala 31:69:@15697.4]
  assign _T_36429 = valid_48_22 ? 6'h16 : _T_36428; // @[Mux.scala 31:69:@15698.4]
  assign _T_36430 = valid_48_21 ? 6'h15 : _T_36429; // @[Mux.scala 31:69:@15699.4]
  assign _T_36431 = valid_48_20 ? 6'h14 : _T_36430; // @[Mux.scala 31:69:@15700.4]
  assign _T_36432 = valid_48_19 ? 6'h13 : _T_36431; // @[Mux.scala 31:69:@15701.4]
  assign _T_36433 = valid_48_18 ? 6'h12 : _T_36432; // @[Mux.scala 31:69:@15702.4]
  assign _T_36434 = valid_48_17 ? 6'h11 : _T_36433; // @[Mux.scala 31:69:@15703.4]
  assign _T_36435 = valid_48_16 ? 6'h10 : _T_36434; // @[Mux.scala 31:69:@15704.4]
  assign _T_36436 = valid_48_15 ? 6'hf : _T_36435; // @[Mux.scala 31:69:@15705.4]
  assign _T_36437 = valid_48_14 ? 6'he : _T_36436; // @[Mux.scala 31:69:@15706.4]
  assign _T_36438 = valid_48_13 ? 6'hd : _T_36437; // @[Mux.scala 31:69:@15707.4]
  assign _T_36439 = valid_48_12 ? 6'hc : _T_36438; // @[Mux.scala 31:69:@15708.4]
  assign _T_36440 = valid_48_11 ? 6'hb : _T_36439; // @[Mux.scala 31:69:@15709.4]
  assign _T_36441 = valid_48_10 ? 6'ha : _T_36440; // @[Mux.scala 31:69:@15710.4]
  assign _T_36442 = valid_48_9 ? 6'h9 : _T_36441; // @[Mux.scala 31:69:@15711.4]
  assign _T_36443 = valid_48_8 ? 6'h8 : _T_36442; // @[Mux.scala 31:69:@15712.4]
  assign _T_36444 = valid_48_7 ? 6'h7 : _T_36443; // @[Mux.scala 31:69:@15713.4]
  assign _T_36445 = valid_48_6 ? 6'h6 : _T_36444; // @[Mux.scala 31:69:@15714.4]
  assign _T_36446 = valid_48_5 ? 6'h5 : _T_36445; // @[Mux.scala 31:69:@15715.4]
  assign _T_36447 = valid_48_4 ? 6'h4 : _T_36446; // @[Mux.scala 31:69:@15716.4]
  assign _T_36448 = valid_48_3 ? 6'h3 : _T_36447; // @[Mux.scala 31:69:@15717.4]
  assign _T_36449 = valid_48_2 ? 6'h2 : _T_36448; // @[Mux.scala 31:69:@15718.4]
  assign _T_36450 = valid_48_1 ? 6'h1 : _T_36449; // @[Mux.scala 31:69:@15719.4]
  assign select_48 = valid_48_0 ? 6'h0 : _T_36450; // @[Mux.scala 31:69:@15720.4]
  assign _GEN_3073 = 6'h1 == select_48 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3074 = 6'h2 == select_48 ? io_inData_2 : _GEN_3073; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3075 = 6'h3 == select_48 ? io_inData_3 : _GEN_3074; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3076 = 6'h4 == select_48 ? io_inData_4 : _GEN_3075; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3077 = 6'h5 == select_48 ? io_inData_5 : _GEN_3076; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3078 = 6'h6 == select_48 ? io_inData_6 : _GEN_3077; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3079 = 6'h7 == select_48 ? io_inData_7 : _GEN_3078; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3080 = 6'h8 == select_48 ? io_inData_8 : _GEN_3079; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3081 = 6'h9 == select_48 ? io_inData_9 : _GEN_3080; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3082 = 6'ha == select_48 ? io_inData_10 : _GEN_3081; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3083 = 6'hb == select_48 ? io_inData_11 : _GEN_3082; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3084 = 6'hc == select_48 ? io_inData_12 : _GEN_3083; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3085 = 6'hd == select_48 ? io_inData_13 : _GEN_3084; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3086 = 6'he == select_48 ? io_inData_14 : _GEN_3085; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3087 = 6'hf == select_48 ? io_inData_15 : _GEN_3086; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3088 = 6'h10 == select_48 ? io_inData_16 : _GEN_3087; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3089 = 6'h11 == select_48 ? io_inData_17 : _GEN_3088; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3090 = 6'h12 == select_48 ? io_inData_18 : _GEN_3089; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3091 = 6'h13 == select_48 ? io_inData_19 : _GEN_3090; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3092 = 6'h14 == select_48 ? io_inData_20 : _GEN_3091; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3093 = 6'h15 == select_48 ? io_inData_21 : _GEN_3092; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3094 = 6'h16 == select_48 ? io_inData_22 : _GEN_3093; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3095 = 6'h17 == select_48 ? io_inData_23 : _GEN_3094; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3096 = 6'h18 == select_48 ? io_inData_24 : _GEN_3095; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3097 = 6'h19 == select_48 ? io_inData_25 : _GEN_3096; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3098 = 6'h1a == select_48 ? io_inData_26 : _GEN_3097; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3099 = 6'h1b == select_48 ? io_inData_27 : _GEN_3098; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3100 = 6'h1c == select_48 ? io_inData_28 : _GEN_3099; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3101 = 6'h1d == select_48 ? io_inData_29 : _GEN_3100; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3102 = 6'h1e == select_48 ? io_inData_30 : _GEN_3101; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3103 = 6'h1f == select_48 ? io_inData_31 : _GEN_3102; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3104 = 6'h20 == select_48 ? io_inData_32 : _GEN_3103; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3105 = 6'h21 == select_48 ? io_inData_33 : _GEN_3104; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3106 = 6'h22 == select_48 ? io_inData_34 : _GEN_3105; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3107 = 6'h23 == select_48 ? io_inData_35 : _GEN_3106; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3108 = 6'h24 == select_48 ? io_inData_36 : _GEN_3107; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3109 = 6'h25 == select_48 ? io_inData_37 : _GEN_3108; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3110 = 6'h26 == select_48 ? io_inData_38 : _GEN_3109; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3111 = 6'h27 == select_48 ? io_inData_39 : _GEN_3110; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3112 = 6'h28 == select_48 ? io_inData_40 : _GEN_3111; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3113 = 6'h29 == select_48 ? io_inData_41 : _GEN_3112; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3114 = 6'h2a == select_48 ? io_inData_42 : _GEN_3113; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3115 = 6'h2b == select_48 ? io_inData_43 : _GEN_3114; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3116 = 6'h2c == select_48 ? io_inData_44 : _GEN_3115; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3117 = 6'h2d == select_48 ? io_inData_45 : _GEN_3116; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3118 = 6'h2e == select_48 ? io_inData_46 : _GEN_3117; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3119 = 6'h2f == select_48 ? io_inData_47 : _GEN_3118; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3120 = 6'h30 == select_48 ? io_inData_48 : _GEN_3119; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3121 = 6'h31 == select_48 ? io_inData_49 : _GEN_3120; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3122 = 6'h32 == select_48 ? io_inData_50 : _GEN_3121; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3123 = 6'h33 == select_48 ? io_inData_51 : _GEN_3122; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3124 = 6'h34 == select_48 ? io_inData_52 : _GEN_3123; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3125 = 6'h35 == select_48 ? io_inData_53 : _GEN_3124; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3126 = 6'h36 == select_48 ? io_inData_54 : _GEN_3125; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3127 = 6'h37 == select_48 ? io_inData_55 : _GEN_3126; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3128 = 6'h38 == select_48 ? io_inData_56 : _GEN_3127; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3129 = 6'h39 == select_48 ? io_inData_57 : _GEN_3128; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3130 = 6'h3a == select_48 ? io_inData_58 : _GEN_3129; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3131 = 6'h3b == select_48 ? io_inData_59 : _GEN_3130; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3132 = 6'h3c == select_48 ? io_inData_60 : _GEN_3131; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3133 = 6'h3d == select_48 ? io_inData_61 : _GEN_3132; // @[Switch.scala 33:19:@15722.4]
  assign _GEN_3134 = 6'h3e == select_48 ? io_inData_62 : _GEN_3133; // @[Switch.scala 33:19:@15722.4]
  assign _T_36459 = {valid_48_7,valid_48_6,valid_48_5,valid_48_4,valid_48_3,valid_48_2,valid_48_1,valid_48_0}; // @[Switch.scala 34:32:@15729.4]
  assign _T_36467 = {valid_48_15,valid_48_14,valid_48_13,valid_48_12,valid_48_11,valid_48_10,valid_48_9,valid_48_8,_T_36459}; // @[Switch.scala 34:32:@15737.4]
  assign _T_36474 = {valid_48_23,valid_48_22,valid_48_21,valid_48_20,valid_48_19,valid_48_18,valid_48_17,valid_48_16}; // @[Switch.scala 34:32:@15744.4]
  assign _T_36483 = {valid_48_31,valid_48_30,valid_48_29,valid_48_28,valid_48_27,valid_48_26,valid_48_25,valid_48_24,_T_36474,_T_36467}; // @[Switch.scala 34:32:@15753.4]
  assign _T_36490 = {valid_48_39,valid_48_38,valid_48_37,valid_48_36,valid_48_35,valid_48_34,valid_48_33,valid_48_32}; // @[Switch.scala 34:32:@15760.4]
  assign _T_36498 = {valid_48_47,valid_48_46,valid_48_45,valid_48_44,valid_48_43,valid_48_42,valid_48_41,valid_48_40,_T_36490}; // @[Switch.scala 34:32:@15768.4]
  assign _T_36505 = {valid_48_55,valid_48_54,valid_48_53,valid_48_52,valid_48_51,valid_48_50,valid_48_49,valid_48_48}; // @[Switch.scala 34:32:@15775.4]
  assign _T_36514 = {valid_48_63,valid_48_62,valid_48_61,valid_48_60,valid_48_59,valid_48_58,valid_48_57,valid_48_56,_T_36505,_T_36498}; // @[Switch.scala 34:32:@15784.4]
  assign _T_36515 = {_T_36514,_T_36483}; // @[Switch.scala 34:32:@15785.4]
  assign _T_36519 = io_inAddr_0 == 6'h31; // @[Switch.scala 30:53:@15788.4]
  assign valid_49_0 = io_inValid_0 & _T_36519; // @[Switch.scala 30:36:@15789.4]
  assign _T_36522 = io_inAddr_1 == 6'h31; // @[Switch.scala 30:53:@15791.4]
  assign valid_49_1 = io_inValid_1 & _T_36522; // @[Switch.scala 30:36:@15792.4]
  assign _T_36525 = io_inAddr_2 == 6'h31; // @[Switch.scala 30:53:@15794.4]
  assign valid_49_2 = io_inValid_2 & _T_36525; // @[Switch.scala 30:36:@15795.4]
  assign _T_36528 = io_inAddr_3 == 6'h31; // @[Switch.scala 30:53:@15797.4]
  assign valid_49_3 = io_inValid_3 & _T_36528; // @[Switch.scala 30:36:@15798.4]
  assign _T_36531 = io_inAddr_4 == 6'h31; // @[Switch.scala 30:53:@15800.4]
  assign valid_49_4 = io_inValid_4 & _T_36531; // @[Switch.scala 30:36:@15801.4]
  assign _T_36534 = io_inAddr_5 == 6'h31; // @[Switch.scala 30:53:@15803.4]
  assign valid_49_5 = io_inValid_5 & _T_36534; // @[Switch.scala 30:36:@15804.4]
  assign _T_36537 = io_inAddr_6 == 6'h31; // @[Switch.scala 30:53:@15806.4]
  assign valid_49_6 = io_inValid_6 & _T_36537; // @[Switch.scala 30:36:@15807.4]
  assign _T_36540 = io_inAddr_7 == 6'h31; // @[Switch.scala 30:53:@15809.4]
  assign valid_49_7 = io_inValid_7 & _T_36540; // @[Switch.scala 30:36:@15810.4]
  assign _T_36543 = io_inAddr_8 == 6'h31; // @[Switch.scala 30:53:@15812.4]
  assign valid_49_8 = io_inValid_8 & _T_36543; // @[Switch.scala 30:36:@15813.4]
  assign _T_36546 = io_inAddr_9 == 6'h31; // @[Switch.scala 30:53:@15815.4]
  assign valid_49_9 = io_inValid_9 & _T_36546; // @[Switch.scala 30:36:@15816.4]
  assign _T_36549 = io_inAddr_10 == 6'h31; // @[Switch.scala 30:53:@15818.4]
  assign valid_49_10 = io_inValid_10 & _T_36549; // @[Switch.scala 30:36:@15819.4]
  assign _T_36552 = io_inAddr_11 == 6'h31; // @[Switch.scala 30:53:@15821.4]
  assign valid_49_11 = io_inValid_11 & _T_36552; // @[Switch.scala 30:36:@15822.4]
  assign _T_36555 = io_inAddr_12 == 6'h31; // @[Switch.scala 30:53:@15824.4]
  assign valid_49_12 = io_inValid_12 & _T_36555; // @[Switch.scala 30:36:@15825.4]
  assign _T_36558 = io_inAddr_13 == 6'h31; // @[Switch.scala 30:53:@15827.4]
  assign valid_49_13 = io_inValid_13 & _T_36558; // @[Switch.scala 30:36:@15828.4]
  assign _T_36561 = io_inAddr_14 == 6'h31; // @[Switch.scala 30:53:@15830.4]
  assign valid_49_14 = io_inValid_14 & _T_36561; // @[Switch.scala 30:36:@15831.4]
  assign _T_36564 = io_inAddr_15 == 6'h31; // @[Switch.scala 30:53:@15833.4]
  assign valid_49_15 = io_inValid_15 & _T_36564; // @[Switch.scala 30:36:@15834.4]
  assign _T_36567 = io_inAddr_16 == 6'h31; // @[Switch.scala 30:53:@15836.4]
  assign valid_49_16 = io_inValid_16 & _T_36567; // @[Switch.scala 30:36:@15837.4]
  assign _T_36570 = io_inAddr_17 == 6'h31; // @[Switch.scala 30:53:@15839.4]
  assign valid_49_17 = io_inValid_17 & _T_36570; // @[Switch.scala 30:36:@15840.4]
  assign _T_36573 = io_inAddr_18 == 6'h31; // @[Switch.scala 30:53:@15842.4]
  assign valid_49_18 = io_inValid_18 & _T_36573; // @[Switch.scala 30:36:@15843.4]
  assign _T_36576 = io_inAddr_19 == 6'h31; // @[Switch.scala 30:53:@15845.4]
  assign valid_49_19 = io_inValid_19 & _T_36576; // @[Switch.scala 30:36:@15846.4]
  assign _T_36579 = io_inAddr_20 == 6'h31; // @[Switch.scala 30:53:@15848.4]
  assign valid_49_20 = io_inValid_20 & _T_36579; // @[Switch.scala 30:36:@15849.4]
  assign _T_36582 = io_inAddr_21 == 6'h31; // @[Switch.scala 30:53:@15851.4]
  assign valid_49_21 = io_inValid_21 & _T_36582; // @[Switch.scala 30:36:@15852.4]
  assign _T_36585 = io_inAddr_22 == 6'h31; // @[Switch.scala 30:53:@15854.4]
  assign valid_49_22 = io_inValid_22 & _T_36585; // @[Switch.scala 30:36:@15855.4]
  assign _T_36588 = io_inAddr_23 == 6'h31; // @[Switch.scala 30:53:@15857.4]
  assign valid_49_23 = io_inValid_23 & _T_36588; // @[Switch.scala 30:36:@15858.4]
  assign _T_36591 = io_inAddr_24 == 6'h31; // @[Switch.scala 30:53:@15860.4]
  assign valid_49_24 = io_inValid_24 & _T_36591; // @[Switch.scala 30:36:@15861.4]
  assign _T_36594 = io_inAddr_25 == 6'h31; // @[Switch.scala 30:53:@15863.4]
  assign valid_49_25 = io_inValid_25 & _T_36594; // @[Switch.scala 30:36:@15864.4]
  assign _T_36597 = io_inAddr_26 == 6'h31; // @[Switch.scala 30:53:@15866.4]
  assign valid_49_26 = io_inValid_26 & _T_36597; // @[Switch.scala 30:36:@15867.4]
  assign _T_36600 = io_inAddr_27 == 6'h31; // @[Switch.scala 30:53:@15869.4]
  assign valid_49_27 = io_inValid_27 & _T_36600; // @[Switch.scala 30:36:@15870.4]
  assign _T_36603 = io_inAddr_28 == 6'h31; // @[Switch.scala 30:53:@15872.4]
  assign valid_49_28 = io_inValid_28 & _T_36603; // @[Switch.scala 30:36:@15873.4]
  assign _T_36606 = io_inAddr_29 == 6'h31; // @[Switch.scala 30:53:@15875.4]
  assign valid_49_29 = io_inValid_29 & _T_36606; // @[Switch.scala 30:36:@15876.4]
  assign _T_36609 = io_inAddr_30 == 6'h31; // @[Switch.scala 30:53:@15878.4]
  assign valid_49_30 = io_inValid_30 & _T_36609; // @[Switch.scala 30:36:@15879.4]
  assign _T_36612 = io_inAddr_31 == 6'h31; // @[Switch.scala 30:53:@15881.4]
  assign valid_49_31 = io_inValid_31 & _T_36612; // @[Switch.scala 30:36:@15882.4]
  assign _T_36615 = io_inAddr_32 == 6'h31; // @[Switch.scala 30:53:@15884.4]
  assign valid_49_32 = io_inValid_32 & _T_36615; // @[Switch.scala 30:36:@15885.4]
  assign _T_36618 = io_inAddr_33 == 6'h31; // @[Switch.scala 30:53:@15887.4]
  assign valid_49_33 = io_inValid_33 & _T_36618; // @[Switch.scala 30:36:@15888.4]
  assign _T_36621 = io_inAddr_34 == 6'h31; // @[Switch.scala 30:53:@15890.4]
  assign valid_49_34 = io_inValid_34 & _T_36621; // @[Switch.scala 30:36:@15891.4]
  assign _T_36624 = io_inAddr_35 == 6'h31; // @[Switch.scala 30:53:@15893.4]
  assign valid_49_35 = io_inValid_35 & _T_36624; // @[Switch.scala 30:36:@15894.4]
  assign _T_36627 = io_inAddr_36 == 6'h31; // @[Switch.scala 30:53:@15896.4]
  assign valid_49_36 = io_inValid_36 & _T_36627; // @[Switch.scala 30:36:@15897.4]
  assign _T_36630 = io_inAddr_37 == 6'h31; // @[Switch.scala 30:53:@15899.4]
  assign valid_49_37 = io_inValid_37 & _T_36630; // @[Switch.scala 30:36:@15900.4]
  assign _T_36633 = io_inAddr_38 == 6'h31; // @[Switch.scala 30:53:@15902.4]
  assign valid_49_38 = io_inValid_38 & _T_36633; // @[Switch.scala 30:36:@15903.4]
  assign _T_36636 = io_inAddr_39 == 6'h31; // @[Switch.scala 30:53:@15905.4]
  assign valid_49_39 = io_inValid_39 & _T_36636; // @[Switch.scala 30:36:@15906.4]
  assign _T_36639 = io_inAddr_40 == 6'h31; // @[Switch.scala 30:53:@15908.4]
  assign valid_49_40 = io_inValid_40 & _T_36639; // @[Switch.scala 30:36:@15909.4]
  assign _T_36642 = io_inAddr_41 == 6'h31; // @[Switch.scala 30:53:@15911.4]
  assign valid_49_41 = io_inValid_41 & _T_36642; // @[Switch.scala 30:36:@15912.4]
  assign _T_36645 = io_inAddr_42 == 6'h31; // @[Switch.scala 30:53:@15914.4]
  assign valid_49_42 = io_inValid_42 & _T_36645; // @[Switch.scala 30:36:@15915.4]
  assign _T_36648 = io_inAddr_43 == 6'h31; // @[Switch.scala 30:53:@15917.4]
  assign valid_49_43 = io_inValid_43 & _T_36648; // @[Switch.scala 30:36:@15918.4]
  assign _T_36651 = io_inAddr_44 == 6'h31; // @[Switch.scala 30:53:@15920.4]
  assign valid_49_44 = io_inValid_44 & _T_36651; // @[Switch.scala 30:36:@15921.4]
  assign _T_36654 = io_inAddr_45 == 6'h31; // @[Switch.scala 30:53:@15923.4]
  assign valid_49_45 = io_inValid_45 & _T_36654; // @[Switch.scala 30:36:@15924.4]
  assign _T_36657 = io_inAddr_46 == 6'h31; // @[Switch.scala 30:53:@15926.4]
  assign valid_49_46 = io_inValid_46 & _T_36657; // @[Switch.scala 30:36:@15927.4]
  assign _T_36660 = io_inAddr_47 == 6'h31; // @[Switch.scala 30:53:@15929.4]
  assign valid_49_47 = io_inValid_47 & _T_36660; // @[Switch.scala 30:36:@15930.4]
  assign _T_36663 = io_inAddr_48 == 6'h31; // @[Switch.scala 30:53:@15932.4]
  assign valid_49_48 = io_inValid_48 & _T_36663; // @[Switch.scala 30:36:@15933.4]
  assign _T_36666 = io_inAddr_49 == 6'h31; // @[Switch.scala 30:53:@15935.4]
  assign valid_49_49 = io_inValid_49 & _T_36666; // @[Switch.scala 30:36:@15936.4]
  assign _T_36669 = io_inAddr_50 == 6'h31; // @[Switch.scala 30:53:@15938.4]
  assign valid_49_50 = io_inValid_50 & _T_36669; // @[Switch.scala 30:36:@15939.4]
  assign _T_36672 = io_inAddr_51 == 6'h31; // @[Switch.scala 30:53:@15941.4]
  assign valid_49_51 = io_inValid_51 & _T_36672; // @[Switch.scala 30:36:@15942.4]
  assign _T_36675 = io_inAddr_52 == 6'h31; // @[Switch.scala 30:53:@15944.4]
  assign valid_49_52 = io_inValid_52 & _T_36675; // @[Switch.scala 30:36:@15945.4]
  assign _T_36678 = io_inAddr_53 == 6'h31; // @[Switch.scala 30:53:@15947.4]
  assign valid_49_53 = io_inValid_53 & _T_36678; // @[Switch.scala 30:36:@15948.4]
  assign _T_36681 = io_inAddr_54 == 6'h31; // @[Switch.scala 30:53:@15950.4]
  assign valid_49_54 = io_inValid_54 & _T_36681; // @[Switch.scala 30:36:@15951.4]
  assign _T_36684 = io_inAddr_55 == 6'h31; // @[Switch.scala 30:53:@15953.4]
  assign valid_49_55 = io_inValid_55 & _T_36684; // @[Switch.scala 30:36:@15954.4]
  assign _T_36687 = io_inAddr_56 == 6'h31; // @[Switch.scala 30:53:@15956.4]
  assign valid_49_56 = io_inValid_56 & _T_36687; // @[Switch.scala 30:36:@15957.4]
  assign _T_36690 = io_inAddr_57 == 6'h31; // @[Switch.scala 30:53:@15959.4]
  assign valid_49_57 = io_inValid_57 & _T_36690; // @[Switch.scala 30:36:@15960.4]
  assign _T_36693 = io_inAddr_58 == 6'h31; // @[Switch.scala 30:53:@15962.4]
  assign valid_49_58 = io_inValid_58 & _T_36693; // @[Switch.scala 30:36:@15963.4]
  assign _T_36696 = io_inAddr_59 == 6'h31; // @[Switch.scala 30:53:@15965.4]
  assign valid_49_59 = io_inValid_59 & _T_36696; // @[Switch.scala 30:36:@15966.4]
  assign _T_36699 = io_inAddr_60 == 6'h31; // @[Switch.scala 30:53:@15968.4]
  assign valid_49_60 = io_inValid_60 & _T_36699; // @[Switch.scala 30:36:@15969.4]
  assign _T_36702 = io_inAddr_61 == 6'h31; // @[Switch.scala 30:53:@15971.4]
  assign valid_49_61 = io_inValid_61 & _T_36702; // @[Switch.scala 30:36:@15972.4]
  assign _T_36705 = io_inAddr_62 == 6'h31; // @[Switch.scala 30:53:@15974.4]
  assign valid_49_62 = io_inValid_62 & _T_36705; // @[Switch.scala 30:36:@15975.4]
  assign _T_36708 = io_inAddr_63 == 6'h31; // @[Switch.scala 30:53:@15977.4]
  assign valid_49_63 = io_inValid_63 & _T_36708; // @[Switch.scala 30:36:@15978.4]
  assign _T_36774 = valid_49_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@15980.4]
  assign _T_36775 = valid_49_61 ? 6'h3d : _T_36774; // @[Mux.scala 31:69:@15981.4]
  assign _T_36776 = valid_49_60 ? 6'h3c : _T_36775; // @[Mux.scala 31:69:@15982.4]
  assign _T_36777 = valid_49_59 ? 6'h3b : _T_36776; // @[Mux.scala 31:69:@15983.4]
  assign _T_36778 = valid_49_58 ? 6'h3a : _T_36777; // @[Mux.scala 31:69:@15984.4]
  assign _T_36779 = valid_49_57 ? 6'h39 : _T_36778; // @[Mux.scala 31:69:@15985.4]
  assign _T_36780 = valid_49_56 ? 6'h38 : _T_36779; // @[Mux.scala 31:69:@15986.4]
  assign _T_36781 = valid_49_55 ? 6'h37 : _T_36780; // @[Mux.scala 31:69:@15987.4]
  assign _T_36782 = valid_49_54 ? 6'h36 : _T_36781; // @[Mux.scala 31:69:@15988.4]
  assign _T_36783 = valid_49_53 ? 6'h35 : _T_36782; // @[Mux.scala 31:69:@15989.4]
  assign _T_36784 = valid_49_52 ? 6'h34 : _T_36783; // @[Mux.scala 31:69:@15990.4]
  assign _T_36785 = valid_49_51 ? 6'h33 : _T_36784; // @[Mux.scala 31:69:@15991.4]
  assign _T_36786 = valid_49_50 ? 6'h32 : _T_36785; // @[Mux.scala 31:69:@15992.4]
  assign _T_36787 = valid_49_49 ? 6'h31 : _T_36786; // @[Mux.scala 31:69:@15993.4]
  assign _T_36788 = valid_49_48 ? 6'h30 : _T_36787; // @[Mux.scala 31:69:@15994.4]
  assign _T_36789 = valid_49_47 ? 6'h2f : _T_36788; // @[Mux.scala 31:69:@15995.4]
  assign _T_36790 = valid_49_46 ? 6'h2e : _T_36789; // @[Mux.scala 31:69:@15996.4]
  assign _T_36791 = valid_49_45 ? 6'h2d : _T_36790; // @[Mux.scala 31:69:@15997.4]
  assign _T_36792 = valid_49_44 ? 6'h2c : _T_36791; // @[Mux.scala 31:69:@15998.4]
  assign _T_36793 = valid_49_43 ? 6'h2b : _T_36792; // @[Mux.scala 31:69:@15999.4]
  assign _T_36794 = valid_49_42 ? 6'h2a : _T_36793; // @[Mux.scala 31:69:@16000.4]
  assign _T_36795 = valid_49_41 ? 6'h29 : _T_36794; // @[Mux.scala 31:69:@16001.4]
  assign _T_36796 = valid_49_40 ? 6'h28 : _T_36795; // @[Mux.scala 31:69:@16002.4]
  assign _T_36797 = valid_49_39 ? 6'h27 : _T_36796; // @[Mux.scala 31:69:@16003.4]
  assign _T_36798 = valid_49_38 ? 6'h26 : _T_36797; // @[Mux.scala 31:69:@16004.4]
  assign _T_36799 = valid_49_37 ? 6'h25 : _T_36798; // @[Mux.scala 31:69:@16005.4]
  assign _T_36800 = valid_49_36 ? 6'h24 : _T_36799; // @[Mux.scala 31:69:@16006.4]
  assign _T_36801 = valid_49_35 ? 6'h23 : _T_36800; // @[Mux.scala 31:69:@16007.4]
  assign _T_36802 = valid_49_34 ? 6'h22 : _T_36801; // @[Mux.scala 31:69:@16008.4]
  assign _T_36803 = valid_49_33 ? 6'h21 : _T_36802; // @[Mux.scala 31:69:@16009.4]
  assign _T_36804 = valid_49_32 ? 6'h20 : _T_36803; // @[Mux.scala 31:69:@16010.4]
  assign _T_36805 = valid_49_31 ? 6'h1f : _T_36804; // @[Mux.scala 31:69:@16011.4]
  assign _T_36806 = valid_49_30 ? 6'h1e : _T_36805; // @[Mux.scala 31:69:@16012.4]
  assign _T_36807 = valid_49_29 ? 6'h1d : _T_36806; // @[Mux.scala 31:69:@16013.4]
  assign _T_36808 = valid_49_28 ? 6'h1c : _T_36807; // @[Mux.scala 31:69:@16014.4]
  assign _T_36809 = valid_49_27 ? 6'h1b : _T_36808; // @[Mux.scala 31:69:@16015.4]
  assign _T_36810 = valid_49_26 ? 6'h1a : _T_36809; // @[Mux.scala 31:69:@16016.4]
  assign _T_36811 = valid_49_25 ? 6'h19 : _T_36810; // @[Mux.scala 31:69:@16017.4]
  assign _T_36812 = valid_49_24 ? 6'h18 : _T_36811; // @[Mux.scala 31:69:@16018.4]
  assign _T_36813 = valid_49_23 ? 6'h17 : _T_36812; // @[Mux.scala 31:69:@16019.4]
  assign _T_36814 = valid_49_22 ? 6'h16 : _T_36813; // @[Mux.scala 31:69:@16020.4]
  assign _T_36815 = valid_49_21 ? 6'h15 : _T_36814; // @[Mux.scala 31:69:@16021.4]
  assign _T_36816 = valid_49_20 ? 6'h14 : _T_36815; // @[Mux.scala 31:69:@16022.4]
  assign _T_36817 = valid_49_19 ? 6'h13 : _T_36816; // @[Mux.scala 31:69:@16023.4]
  assign _T_36818 = valid_49_18 ? 6'h12 : _T_36817; // @[Mux.scala 31:69:@16024.4]
  assign _T_36819 = valid_49_17 ? 6'h11 : _T_36818; // @[Mux.scala 31:69:@16025.4]
  assign _T_36820 = valid_49_16 ? 6'h10 : _T_36819; // @[Mux.scala 31:69:@16026.4]
  assign _T_36821 = valid_49_15 ? 6'hf : _T_36820; // @[Mux.scala 31:69:@16027.4]
  assign _T_36822 = valid_49_14 ? 6'he : _T_36821; // @[Mux.scala 31:69:@16028.4]
  assign _T_36823 = valid_49_13 ? 6'hd : _T_36822; // @[Mux.scala 31:69:@16029.4]
  assign _T_36824 = valid_49_12 ? 6'hc : _T_36823; // @[Mux.scala 31:69:@16030.4]
  assign _T_36825 = valid_49_11 ? 6'hb : _T_36824; // @[Mux.scala 31:69:@16031.4]
  assign _T_36826 = valid_49_10 ? 6'ha : _T_36825; // @[Mux.scala 31:69:@16032.4]
  assign _T_36827 = valid_49_9 ? 6'h9 : _T_36826; // @[Mux.scala 31:69:@16033.4]
  assign _T_36828 = valid_49_8 ? 6'h8 : _T_36827; // @[Mux.scala 31:69:@16034.4]
  assign _T_36829 = valid_49_7 ? 6'h7 : _T_36828; // @[Mux.scala 31:69:@16035.4]
  assign _T_36830 = valid_49_6 ? 6'h6 : _T_36829; // @[Mux.scala 31:69:@16036.4]
  assign _T_36831 = valid_49_5 ? 6'h5 : _T_36830; // @[Mux.scala 31:69:@16037.4]
  assign _T_36832 = valid_49_4 ? 6'h4 : _T_36831; // @[Mux.scala 31:69:@16038.4]
  assign _T_36833 = valid_49_3 ? 6'h3 : _T_36832; // @[Mux.scala 31:69:@16039.4]
  assign _T_36834 = valid_49_2 ? 6'h2 : _T_36833; // @[Mux.scala 31:69:@16040.4]
  assign _T_36835 = valid_49_1 ? 6'h1 : _T_36834; // @[Mux.scala 31:69:@16041.4]
  assign select_49 = valid_49_0 ? 6'h0 : _T_36835; // @[Mux.scala 31:69:@16042.4]
  assign _GEN_3137 = 6'h1 == select_49 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3138 = 6'h2 == select_49 ? io_inData_2 : _GEN_3137; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3139 = 6'h3 == select_49 ? io_inData_3 : _GEN_3138; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3140 = 6'h4 == select_49 ? io_inData_4 : _GEN_3139; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3141 = 6'h5 == select_49 ? io_inData_5 : _GEN_3140; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3142 = 6'h6 == select_49 ? io_inData_6 : _GEN_3141; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3143 = 6'h7 == select_49 ? io_inData_7 : _GEN_3142; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3144 = 6'h8 == select_49 ? io_inData_8 : _GEN_3143; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3145 = 6'h9 == select_49 ? io_inData_9 : _GEN_3144; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3146 = 6'ha == select_49 ? io_inData_10 : _GEN_3145; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3147 = 6'hb == select_49 ? io_inData_11 : _GEN_3146; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3148 = 6'hc == select_49 ? io_inData_12 : _GEN_3147; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3149 = 6'hd == select_49 ? io_inData_13 : _GEN_3148; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3150 = 6'he == select_49 ? io_inData_14 : _GEN_3149; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3151 = 6'hf == select_49 ? io_inData_15 : _GEN_3150; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3152 = 6'h10 == select_49 ? io_inData_16 : _GEN_3151; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3153 = 6'h11 == select_49 ? io_inData_17 : _GEN_3152; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3154 = 6'h12 == select_49 ? io_inData_18 : _GEN_3153; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3155 = 6'h13 == select_49 ? io_inData_19 : _GEN_3154; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3156 = 6'h14 == select_49 ? io_inData_20 : _GEN_3155; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3157 = 6'h15 == select_49 ? io_inData_21 : _GEN_3156; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3158 = 6'h16 == select_49 ? io_inData_22 : _GEN_3157; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3159 = 6'h17 == select_49 ? io_inData_23 : _GEN_3158; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3160 = 6'h18 == select_49 ? io_inData_24 : _GEN_3159; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3161 = 6'h19 == select_49 ? io_inData_25 : _GEN_3160; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3162 = 6'h1a == select_49 ? io_inData_26 : _GEN_3161; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3163 = 6'h1b == select_49 ? io_inData_27 : _GEN_3162; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3164 = 6'h1c == select_49 ? io_inData_28 : _GEN_3163; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3165 = 6'h1d == select_49 ? io_inData_29 : _GEN_3164; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3166 = 6'h1e == select_49 ? io_inData_30 : _GEN_3165; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3167 = 6'h1f == select_49 ? io_inData_31 : _GEN_3166; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3168 = 6'h20 == select_49 ? io_inData_32 : _GEN_3167; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3169 = 6'h21 == select_49 ? io_inData_33 : _GEN_3168; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3170 = 6'h22 == select_49 ? io_inData_34 : _GEN_3169; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3171 = 6'h23 == select_49 ? io_inData_35 : _GEN_3170; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3172 = 6'h24 == select_49 ? io_inData_36 : _GEN_3171; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3173 = 6'h25 == select_49 ? io_inData_37 : _GEN_3172; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3174 = 6'h26 == select_49 ? io_inData_38 : _GEN_3173; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3175 = 6'h27 == select_49 ? io_inData_39 : _GEN_3174; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3176 = 6'h28 == select_49 ? io_inData_40 : _GEN_3175; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3177 = 6'h29 == select_49 ? io_inData_41 : _GEN_3176; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3178 = 6'h2a == select_49 ? io_inData_42 : _GEN_3177; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3179 = 6'h2b == select_49 ? io_inData_43 : _GEN_3178; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3180 = 6'h2c == select_49 ? io_inData_44 : _GEN_3179; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3181 = 6'h2d == select_49 ? io_inData_45 : _GEN_3180; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3182 = 6'h2e == select_49 ? io_inData_46 : _GEN_3181; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3183 = 6'h2f == select_49 ? io_inData_47 : _GEN_3182; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3184 = 6'h30 == select_49 ? io_inData_48 : _GEN_3183; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3185 = 6'h31 == select_49 ? io_inData_49 : _GEN_3184; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3186 = 6'h32 == select_49 ? io_inData_50 : _GEN_3185; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3187 = 6'h33 == select_49 ? io_inData_51 : _GEN_3186; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3188 = 6'h34 == select_49 ? io_inData_52 : _GEN_3187; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3189 = 6'h35 == select_49 ? io_inData_53 : _GEN_3188; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3190 = 6'h36 == select_49 ? io_inData_54 : _GEN_3189; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3191 = 6'h37 == select_49 ? io_inData_55 : _GEN_3190; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3192 = 6'h38 == select_49 ? io_inData_56 : _GEN_3191; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3193 = 6'h39 == select_49 ? io_inData_57 : _GEN_3192; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3194 = 6'h3a == select_49 ? io_inData_58 : _GEN_3193; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3195 = 6'h3b == select_49 ? io_inData_59 : _GEN_3194; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3196 = 6'h3c == select_49 ? io_inData_60 : _GEN_3195; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3197 = 6'h3d == select_49 ? io_inData_61 : _GEN_3196; // @[Switch.scala 33:19:@16044.4]
  assign _GEN_3198 = 6'h3e == select_49 ? io_inData_62 : _GEN_3197; // @[Switch.scala 33:19:@16044.4]
  assign _T_36844 = {valid_49_7,valid_49_6,valid_49_5,valid_49_4,valid_49_3,valid_49_2,valid_49_1,valid_49_0}; // @[Switch.scala 34:32:@16051.4]
  assign _T_36852 = {valid_49_15,valid_49_14,valid_49_13,valid_49_12,valid_49_11,valid_49_10,valid_49_9,valid_49_8,_T_36844}; // @[Switch.scala 34:32:@16059.4]
  assign _T_36859 = {valid_49_23,valid_49_22,valid_49_21,valid_49_20,valid_49_19,valid_49_18,valid_49_17,valid_49_16}; // @[Switch.scala 34:32:@16066.4]
  assign _T_36868 = {valid_49_31,valid_49_30,valid_49_29,valid_49_28,valid_49_27,valid_49_26,valid_49_25,valid_49_24,_T_36859,_T_36852}; // @[Switch.scala 34:32:@16075.4]
  assign _T_36875 = {valid_49_39,valid_49_38,valid_49_37,valid_49_36,valid_49_35,valid_49_34,valid_49_33,valid_49_32}; // @[Switch.scala 34:32:@16082.4]
  assign _T_36883 = {valid_49_47,valid_49_46,valid_49_45,valid_49_44,valid_49_43,valid_49_42,valid_49_41,valid_49_40,_T_36875}; // @[Switch.scala 34:32:@16090.4]
  assign _T_36890 = {valid_49_55,valid_49_54,valid_49_53,valid_49_52,valid_49_51,valid_49_50,valid_49_49,valid_49_48}; // @[Switch.scala 34:32:@16097.4]
  assign _T_36899 = {valid_49_63,valid_49_62,valid_49_61,valid_49_60,valid_49_59,valid_49_58,valid_49_57,valid_49_56,_T_36890,_T_36883}; // @[Switch.scala 34:32:@16106.4]
  assign _T_36900 = {_T_36899,_T_36868}; // @[Switch.scala 34:32:@16107.4]
  assign _T_36904 = io_inAddr_0 == 6'h32; // @[Switch.scala 30:53:@16110.4]
  assign valid_50_0 = io_inValid_0 & _T_36904; // @[Switch.scala 30:36:@16111.4]
  assign _T_36907 = io_inAddr_1 == 6'h32; // @[Switch.scala 30:53:@16113.4]
  assign valid_50_1 = io_inValid_1 & _T_36907; // @[Switch.scala 30:36:@16114.4]
  assign _T_36910 = io_inAddr_2 == 6'h32; // @[Switch.scala 30:53:@16116.4]
  assign valid_50_2 = io_inValid_2 & _T_36910; // @[Switch.scala 30:36:@16117.4]
  assign _T_36913 = io_inAddr_3 == 6'h32; // @[Switch.scala 30:53:@16119.4]
  assign valid_50_3 = io_inValid_3 & _T_36913; // @[Switch.scala 30:36:@16120.4]
  assign _T_36916 = io_inAddr_4 == 6'h32; // @[Switch.scala 30:53:@16122.4]
  assign valid_50_4 = io_inValid_4 & _T_36916; // @[Switch.scala 30:36:@16123.4]
  assign _T_36919 = io_inAddr_5 == 6'h32; // @[Switch.scala 30:53:@16125.4]
  assign valid_50_5 = io_inValid_5 & _T_36919; // @[Switch.scala 30:36:@16126.4]
  assign _T_36922 = io_inAddr_6 == 6'h32; // @[Switch.scala 30:53:@16128.4]
  assign valid_50_6 = io_inValid_6 & _T_36922; // @[Switch.scala 30:36:@16129.4]
  assign _T_36925 = io_inAddr_7 == 6'h32; // @[Switch.scala 30:53:@16131.4]
  assign valid_50_7 = io_inValid_7 & _T_36925; // @[Switch.scala 30:36:@16132.4]
  assign _T_36928 = io_inAddr_8 == 6'h32; // @[Switch.scala 30:53:@16134.4]
  assign valid_50_8 = io_inValid_8 & _T_36928; // @[Switch.scala 30:36:@16135.4]
  assign _T_36931 = io_inAddr_9 == 6'h32; // @[Switch.scala 30:53:@16137.4]
  assign valid_50_9 = io_inValid_9 & _T_36931; // @[Switch.scala 30:36:@16138.4]
  assign _T_36934 = io_inAddr_10 == 6'h32; // @[Switch.scala 30:53:@16140.4]
  assign valid_50_10 = io_inValid_10 & _T_36934; // @[Switch.scala 30:36:@16141.4]
  assign _T_36937 = io_inAddr_11 == 6'h32; // @[Switch.scala 30:53:@16143.4]
  assign valid_50_11 = io_inValid_11 & _T_36937; // @[Switch.scala 30:36:@16144.4]
  assign _T_36940 = io_inAddr_12 == 6'h32; // @[Switch.scala 30:53:@16146.4]
  assign valid_50_12 = io_inValid_12 & _T_36940; // @[Switch.scala 30:36:@16147.4]
  assign _T_36943 = io_inAddr_13 == 6'h32; // @[Switch.scala 30:53:@16149.4]
  assign valid_50_13 = io_inValid_13 & _T_36943; // @[Switch.scala 30:36:@16150.4]
  assign _T_36946 = io_inAddr_14 == 6'h32; // @[Switch.scala 30:53:@16152.4]
  assign valid_50_14 = io_inValid_14 & _T_36946; // @[Switch.scala 30:36:@16153.4]
  assign _T_36949 = io_inAddr_15 == 6'h32; // @[Switch.scala 30:53:@16155.4]
  assign valid_50_15 = io_inValid_15 & _T_36949; // @[Switch.scala 30:36:@16156.4]
  assign _T_36952 = io_inAddr_16 == 6'h32; // @[Switch.scala 30:53:@16158.4]
  assign valid_50_16 = io_inValid_16 & _T_36952; // @[Switch.scala 30:36:@16159.4]
  assign _T_36955 = io_inAddr_17 == 6'h32; // @[Switch.scala 30:53:@16161.4]
  assign valid_50_17 = io_inValid_17 & _T_36955; // @[Switch.scala 30:36:@16162.4]
  assign _T_36958 = io_inAddr_18 == 6'h32; // @[Switch.scala 30:53:@16164.4]
  assign valid_50_18 = io_inValid_18 & _T_36958; // @[Switch.scala 30:36:@16165.4]
  assign _T_36961 = io_inAddr_19 == 6'h32; // @[Switch.scala 30:53:@16167.4]
  assign valid_50_19 = io_inValid_19 & _T_36961; // @[Switch.scala 30:36:@16168.4]
  assign _T_36964 = io_inAddr_20 == 6'h32; // @[Switch.scala 30:53:@16170.4]
  assign valid_50_20 = io_inValid_20 & _T_36964; // @[Switch.scala 30:36:@16171.4]
  assign _T_36967 = io_inAddr_21 == 6'h32; // @[Switch.scala 30:53:@16173.4]
  assign valid_50_21 = io_inValid_21 & _T_36967; // @[Switch.scala 30:36:@16174.4]
  assign _T_36970 = io_inAddr_22 == 6'h32; // @[Switch.scala 30:53:@16176.4]
  assign valid_50_22 = io_inValid_22 & _T_36970; // @[Switch.scala 30:36:@16177.4]
  assign _T_36973 = io_inAddr_23 == 6'h32; // @[Switch.scala 30:53:@16179.4]
  assign valid_50_23 = io_inValid_23 & _T_36973; // @[Switch.scala 30:36:@16180.4]
  assign _T_36976 = io_inAddr_24 == 6'h32; // @[Switch.scala 30:53:@16182.4]
  assign valid_50_24 = io_inValid_24 & _T_36976; // @[Switch.scala 30:36:@16183.4]
  assign _T_36979 = io_inAddr_25 == 6'h32; // @[Switch.scala 30:53:@16185.4]
  assign valid_50_25 = io_inValid_25 & _T_36979; // @[Switch.scala 30:36:@16186.4]
  assign _T_36982 = io_inAddr_26 == 6'h32; // @[Switch.scala 30:53:@16188.4]
  assign valid_50_26 = io_inValid_26 & _T_36982; // @[Switch.scala 30:36:@16189.4]
  assign _T_36985 = io_inAddr_27 == 6'h32; // @[Switch.scala 30:53:@16191.4]
  assign valid_50_27 = io_inValid_27 & _T_36985; // @[Switch.scala 30:36:@16192.4]
  assign _T_36988 = io_inAddr_28 == 6'h32; // @[Switch.scala 30:53:@16194.4]
  assign valid_50_28 = io_inValid_28 & _T_36988; // @[Switch.scala 30:36:@16195.4]
  assign _T_36991 = io_inAddr_29 == 6'h32; // @[Switch.scala 30:53:@16197.4]
  assign valid_50_29 = io_inValid_29 & _T_36991; // @[Switch.scala 30:36:@16198.4]
  assign _T_36994 = io_inAddr_30 == 6'h32; // @[Switch.scala 30:53:@16200.4]
  assign valid_50_30 = io_inValid_30 & _T_36994; // @[Switch.scala 30:36:@16201.4]
  assign _T_36997 = io_inAddr_31 == 6'h32; // @[Switch.scala 30:53:@16203.4]
  assign valid_50_31 = io_inValid_31 & _T_36997; // @[Switch.scala 30:36:@16204.4]
  assign _T_37000 = io_inAddr_32 == 6'h32; // @[Switch.scala 30:53:@16206.4]
  assign valid_50_32 = io_inValid_32 & _T_37000; // @[Switch.scala 30:36:@16207.4]
  assign _T_37003 = io_inAddr_33 == 6'h32; // @[Switch.scala 30:53:@16209.4]
  assign valid_50_33 = io_inValid_33 & _T_37003; // @[Switch.scala 30:36:@16210.4]
  assign _T_37006 = io_inAddr_34 == 6'h32; // @[Switch.scala 30:53:@16212.4]
  assign valid_50_34 = io_inValid_34 & _T_37006; // @[Switch.scala 30:36:@16213.4]
  assign _T_37009 = io_inAddr_35 == 6'h32; // @[Switch.scala 30:53:@16215.4]
  assign valid_50_35 = io_inValid_35 & _T_37009; // @[Switch.scala 30:36:@16216.4]
  assign _T_37012 = io_inAddr_36 == 6'h32; // @[Switch.scala 30:53:@16218.4]
  assign valid_50_36 = io_inValid_36 & _T_37012; // @[Switch.scala 30:36:@16219.4]
  assign _T_37015 = io_inAddr_37 == 6'h32; // @[Switch.scala 30:53:@16221.4]
  assign valid_50_37 = io_inValid_37 & _T_37015; // @[Switch.scala 30:36:@16222.4]
  assign _T_37018 = io_inAddr_38 == 6'h32; // @[Switch.scala 30:53:@16224.4]
  assign valid_50_38 = io_inValid_38 & _T_37018; // @[Switch.scala 30:36:@16225.4]
  assign _T_37021 = io_inAddr_39 == 6'h32; // @[Switch.scala 30:53:@16227.4]
  assign valid_50_39 = io_inValid_39 & _T_37021; // @[Switch.scala 30:36:@16228.4]
  assign _T_37024 = io_inAddr_40 == 6'h32; // @[Switch.scala 30:53:@16230.4]
  assign valid_50_40 = io_inValid_40 & _T_37024; // @[Switch.scala 30:36:@16231.4]
  assign _T_37027 = io_inAddr_41 == 6'h32; // @[Switch.scala 30:53:@16233.4]
  assign valid_50_41 = io_inValid_41 & _T_37027; // @[Switch.scala 30:36:@16234.4]
  assign _T_37030 = io_inAddr_42 == 6'h32; // @[Switch.scala 30:53:@16236.4]
  assign valid_50_42 = io_inValid_42 & _T_37030; // @[Switch.scala 30:36:@16237.4]
  assign _T_37033 = io_inAddr_43 == 6'h32; // @[Switch.scala 30:53:@16239.4]
  assign valid_50_43 = io_inValid_43 & _T_37033; // @[Switch.scala 30:36:@16240.4]
  assign _T_37036 = io_inAddr_44 == 6'h32; // @[Switch.scala 30:53:@16242.4]
  assign valid_50_44 = io_inValid_44 & _T_37036; // @[Switch.scala 30:36:@16243.4]
  assign _T_37039 = io_inAddr_45 == 6'h32; // @[Switch.scala 30:53:@16245.4]
  assign valid_50_45 = io_inValid_45 & _T_37039; // @[Switch.scala 30:36:@16246.4]
  assign _T_37042 = io_inAddr_46 == 6'h32; // @[Switch.scala 30:53:@16248.4]
  assign valid_50_46 = io_inValid_46 & _T_37042; // @[Switch.scala 30:36:@16249.4]
  assign _T_37045 = io_inAddr_47 == 6'h32; // @[Switch.scala 30:53:@16251.4]
  assign valid_50_47 = io_inValid_47 & _T_37045; // @[Switch.scala 30:36:@16252.4]
  assign _T_37048 = io_inAddr_48 == 6'h32; // @[Switch.scala 30:53:@16254.4]
  assign valid_50_48 = io_inValid_48 & _T_37048; // @[Switch.scala 30:36:@16255.4]
  assign _T_37051 = io_inAddr_49 == 6'h32; // @[Switch.scala 30:53:@16257.4]
  assign valid_50_49 = io_inValid_49 & _T_37051; // @[Switch.scala 30:36:@16258.4]
  assign _T_37054 = io_inAddr_50 == 6'h32; // @[Switch.scala 30:53:@16260.4]
  assign valid_50_50 = io_inValid_50 & _T_37054; // @[Switch.scala 30:36:@16261.4]
  assign _T_37057 = io_inAddr_51 == 6'h32; // @[Switch.scala 30:53:@16263.4]
  assign valid_50_51 = io_inValid_51 & _T_37057; // @[Switch.scala 30:36:@16264.4]
  assign _T_37060 = io_inAddr_52 == 6'h32; // @[Switch.scala 30:53:@16266.4]
  assign valid_50_52 = io_inValid_52 & _T_37060; // @[Switch.scala 30:36:@16267.4]
  assign _T_37063 = io_inAddr_53 == 6'h32; // @[Switch.scala 30:53:@16269.4]
  assign valid_50_53 = io_inValid_53 & _T_37063; // @[Switch.scala 30:36:@16270.4]
  assign _T_37066 = io_inAddr_54 == 6'h32; // @[Switch.scala 30:53:@16272.4]
  assign valid_50_54 = io_inValid_54 & _T_37066; // @[Switch.scala 30:36:@16273.4]
  assign _T_37069 = io_inAddr_55 == 6'h32; // @[Switch.scala 30:53:@16275.4]
  assign valid_50_55 = io_inValid_55 & _T_37069; // @[Switch.scala 30:36:@16276.4]
  assign _T_37072 = io_inAddr_56 == 6'h32; // @[Switch.scala 30:53:@16278.4]
  assign valid_50_56 = io_inValid_56 & _T_37072; // @[Switch.scala 30:36:@16279.4]
  assign _T_37075 = io_inAddr_57 == 6'h32; // @[Switch.scala 30:53:@16281.4]
  assign valid_50_57 = io_inValid_57 & _T_37075; // @[Switch.scala 30:36:@16282.4]
  assign _T_37078 = io_inAddr_58 == 6'h32; // @[Switch.scala 30:53:@16284.4]
  assign valid_50_58 = io_inValid_58 & _T_37078; // @[Switch.scala 30:36:@16285.4]
  assign _T_37081 = io_inAddr_59 == 6'h32; // @[Switch.scala 30:53:@16287.4]
  assign valid_50_59 = io_inValid_59 & _T_37081; // @[Switch.scala 30:36:@16288.4]
  assign _T_37084 = io_inAddr_60 == 6'h32; // @[Switch.scala 30:53:@16290.4]
  assign valid_50_60 = io_inValid_60 & _T_37084; // @[Switch.scala 30:36:@16291.4]
  assign _T_37087 = io_inAddr_61 == 6'h32; // @[Switch.scala 30:53:@16293.4]
  assign valid_50_61 = io_inValid_61 & _T_37087; // @[Switch.scala 30:36:@16294.4]
  assign _T_37090 = io_inAddr_62 == 6'h32; // @[Switch.scala 30:53:@16296.4]
  assign valid_50_62 = io_inValid_62 & _T_37090; // @[Switch.scala 30:36:@16297.4]
  assign _T_37093 = io_inAddr_63 == 6'h32; // @[Switch.scala 30:53:@16299.4]
  assign valid_50_63 = io_inValid_63 & _T_37093; // @[Switch.scala 30:36:@16300.4]
  assign _T_37159 = valid_50_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@16302.4]
  assign _T_37160 = valid_50_61 ? 6'h3d : _T_37159; // @[Mux.scala 31:69:@16303.4]
  assign _T_37161 = valid_50_60 ? 6'h3c : _T_37160; // @[Mux.scala 31:69:@16304.4]
  assign _T_37162 = valid_50_59 ? 6'h3b : _T_37161; // @[Mux.scala 31:69:@16305.4]
  assign _T_37163 = valid_50_58 ? 6'h3a : _T_37162; // @[Mux.scala 31:69:@16306.4]
  assign _T_37164 = valid_50_57 ? 6'h39 : _T_37163; // @[Mux.scala 31:69:@16307.4]
  assign _T_37165 = valid_50_56 ? 6'h38 : _T_37164; // @[Mux.scala 31:69:@16308.4]
  assign _T_37166 = valid_50_55 ? 6'h37 : _T_37165; // @[Mux.scala 31:69:@16309.4]
  assign _T_37167 = valid_50_54 ? 6'h36 : _T_37166; // @[Mux.scala 31:69:@16310.4]
  assign _T_37168 = valid_50_53 ? 6'h35 : _T_37167; // @[Mux.scala 31:69:@16311.4]
  assign _T_37169 = valid_50_52 ? 6'h34 : _T_37168; // @[Mux.scala 31:69:@16312.4]
  assign _T_37170 = valid_50_51 ? 6'h33 : _T_37169; // @[Mux.scala 31:69:@16313.4]
  assign _T_37171 = valid_50_50 ? 6'h32 : _T_37170; // @[Mux.scala 31:69:@16314.4]
  assign _T_37172 = valid_50_49 ? 6'h31 : _T_37171; // @[Mux.scala 31:69:@16315.4]
  assign _T_37173 = valid_50_48 ? 6'h30 : _T_37172; // @[Mux.scala 31:69:@16316.4]
  assign _T_37174 = valid_50_47 ? 6'h2f : _T_37173; // @[Mux.scala 31:69:@16317.4]
  assign _T_37175 = valid_50_46 ? 6'h2e : _T_37174; // @[Mux.scala 31:69:@16318.4]
  assign _T_37176 = valid_50_45 ? 6'h2d : _T_37175; // @[Mux.scala 31:69:@16319.4]
  assign _T_37177 = valid_50_44 ? 6'h2c : _T_37176; // @[Mux.scala 31:69:@16320.4]
  assign _T_37178 = valid_50_43 ? 6'h2b : _T_37177; // @[Mux.scala 31:69:@16321.4]
  assign _T_37179 = valid_50_42 ? 6'h2a : _T_37178; // @[Mux.scala 31:69:@16322.4]
  assign _T_37180 = valid_50_41 ? 6'h29 : _T_37179; // @[Mux.scala 31:69:@16323.4]
  assign _T_37181 = valid_50_40 ? 6'h28 : _T_37180; // @[Mux.scala 31:69:@16324.4]
  assign _T_37182 = valid_50_39 ? 6'h27 : _T_37181; // @[Mux.scala 31:69:@16325.4]
  assign _T_37183 = valid_50_38 ? 6'h26 : _T_37182; // @[Mux.scala 31:69:@16326.4]
  assign _T_37184 = valid_50_37 ? 6'h25 : _T_37183; // @[Mux.scala 31:69:@16327.4]
  assign _T_37185 = valid_50_36 ? 6'h24 : _T_37184; // @[Mux.scala 31:69:@16328.4]
  assign _T_37186 = valid_50_35 ? 6'h23 : _T_37185; // @[Mux.scala 31:69:@16329.4]
  assign _T_37187 = valid_50_34 ? 6'h22 : _T_37186; // @[Mux.scala 31:69:@16330.4]
  assign _T_37188 = valid_50_33 ? 6'h21 : _T_37187; // @[Mux.scala 31:69:@16331.4]
  assign _T_37189 = valid_50_32 ? 6'h20 : _T_37188; // @[Mux.scala 31:69:@16332.4]
  assign _T_37190 = valid_50_31 ? 6'h1f : _T_37189; // @[Mux.scala 31:69:@16333.4]
  assign _T_37191 = valid_50_30 ? 6'h1e : _T_37190; // @[Mux.scala 31:69:@16334.4]
  assign _T_37192 = valid_50_29 ? 6'h1d : _T_37191; // @[Mux.scala 31:69:@16335.4]
  assign _T_37193 = valid_50_28 ? 6'h1c : _T_37192; // @[Mux.scala 31:69:@16336.4]
  assign _T_37194 = valid_50_27 ? 6'h1b : _T_37193; // @[Mux.scala 31:69:@16337.4]
  assign _T_37195 = valid_50_26 ? 6'h1a : _T_37194; // @[Mux.scala 31:69:@16338.4]
  assign _T_37196 = valid_50_25 ? 6'h19 : _T_37195; // @[Mux.scala 31:69:@16339.4]
  assign _T_37197 = valid_50_24 ? 6'h18 : _T_37196; // @[Mux.scala 31:69:@16340.4]
  assign _T_37198 = valid_50_23 ? 6'h17 : _T_37197; // @[Mux.scala 31:69:@16341.4]
  assign _T_37199 = valid_50_22 ? 6'h16 : _T_37198; // @[Mux.scala 31:69:@16342.4]
  assign _T_37200 = valid_50_21 ? 6'h15 : _T_37199; // @[Mux.scala 31:69:@16343.4]
  assign _T_37201 = valid_50_20 ? 6'h14 : _T_37200; // @[Mux.scala 31:69:@16344.4]
  assign _T_37202 = valid_50_19 ? 6'h13 : _T_37201; // @[Mux.scala 31:69:@16345.4]
  assign _T_37203 = valid_50_18 ? 6'h12 : _T_37202; // @[Mux.scala 31:69:@16346.4]
  assign _T_37204 = valid_50_17 ? 6'h11 : _T_37203; // @[Mux.scala 31:69:@16347.4]
  assign _T_37205 = valid_50_16 ? 6'h10 : _T_37204; // @[Mux.scala 31:69:@16348.4]
  assign _T_37206 = valid_50_15 ? 6'hf : _T_37205; // @[Mux.scala 31:69:@16349.4]
  assign _T_37207 = valid_50_14 ? 6'he : _T_37206; // @[Mux.scala 31:69:@16350.4]
  assign _T_37208 = valid_50_13 ? 6'hd : _T_37207; // @[Mux.scala 31:69:@16351.4]
  assign _T_37209 = valid_50_12 ? 6'hc : _T_37208; // @[Mux.scala 31:69:@16352.4]
  assign _T_37210 = valid_50_11 ? 6'hb : _T_37209; // @[Mux.scala 31:69:@16353.4]
  assign _T_37211 = valid_50_10 ? 6'ha : _T_37210; // @[Mux.scala 31:69:@16354.4]
  assign _T_37212 = valid_50_9 ? 6'h9 : _T_37211; // @[Mux.scala 31:69:@16355.4]
  assign _T_37213 = valid_50_8 ? 6'h8 : _T_37212; // @[Mux.scala 31:69:@16356.4]
  assign _T_37214 = valid_50_7 ? 6'h7 : _T_37213; // @[Mux.scala 31:69:@16357.4]
  assign _T_37215 = valid_50_6 ? 6'h6 : _T_37214; // @[Mux.scala 31:69:@16358.4]
  assign _T_37216 = valid_50_5 ? 6'h5 : _T_37215; // @[Mux.scala 31:69:@16359.4]
  assign _T_37217 = valid_50_4 ? 6'h4 : _T_37216; // @[Mux.scala 31:69:@16360.4]
  assign _T_37218 = valid_50_3 ? 6'h3 : _T_37217; // @[Mux.scala 31:69:@16361.4]
  assign _T_37219 = valid_50_2 ? 6'h2 : _T_37218; // @[Mux.scala 31:69:@16362.4]
  assign _T_37220 = valid_50_1 ? 6'h1 : _T_37219; // @[Mux.scala 31:69:@16363.4]
  assign select_50 = valid_50_0 ? 6'h0 : _T_37220; // @[Mux.scala 31:69:@16364.4]
  assign _GEN_3201 = 6'h1 == select_50 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3202 = 6'h2 == select_50 ? io_inData_2 : _GEN_3201; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3203 = 6'h3 == select_50 ? io_inData_3 : _GEN_3202; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3204 = 6'h4 == select_50 ? io_inData_4 : _GEN_3203; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3205 = 6'h5 == select_50 ? io_inData_5 : _GEN_3204; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3206 = 6'h6 == select_50 ? io_inData_6 : _GEN_3205; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3207 = 6'h7 == select_50 ? io_inData_7 : _GEN_3206; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3208 = 6'h8 == select_50 ? io_inData_8 : _GEN_3207; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3209 = 6'h9 == select_50 ? io_inData_9 : _GEN_3208; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3210 = 6'ha == select_50 ? io_inData_10 : _GEN_3209; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3211 = 6'hb == select_50 ? io_inData_11 : _GEN_3210; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3212 = 6'hc == select_50 ? io_inData_12 : _GEN_3211; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3213 = 6'hd == select_50 ? io_inData_13 : _GEN_3212; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3214 = 6'he == select_50 ? io_inData_14 : _GEN_3213; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3215 = 6'hf == select_50 ? io_inData_15 : _GEN_3214; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3216 = 6'h10 == select_50 ? io_inData_16 : _GEN_3215; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3217 = 6'h11 == select_50 ? io_inData_17 : _GEN_3216; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3218 = 6'h12 == select_50 ? io_inData_18 : _GEN_3217; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3219 = 6'h13 == select_50 ? io_inData_19 : _GEN_3218; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3220 = 6'h14 == select_50 ? io_inData_20 : _GEN_3219; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3221 = 6'h15 == select_50 ? io_inData_21 : _GEN_3220; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3222 = 6'h16 == select_50 ? io_inData_22 : _GEN_3221; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3223 = 6'h17 == select_50 ? io_inData_23 : _GEN_3222; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3224 = 6'h18 == select_50 ? io_inData_24 : _GEN_3223; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3225 = 6'h19 == select_50 ? io_inData_25 : _GEN_3224; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3226 = 6'h1a == select_50 ? io_inData_26 : _GEN_3225; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3227 = 6'h1b == select_50 ? io_inData_27 : _GEN_3226; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3228 = 6'h1c == select_50 ? io_inData_28 : _GEN_3227; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3229 = 6'h1d == select_50 ? io_inData_29 : _GEN_3228; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3230 = 6'h1e == select_50 ? io_inData_30 : _GEN_3229; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3231 = 6'h1f == select_50 ? io_inData_31 : _GEN_3230; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3232 = 6'h20 == select_50 ? io_inData_32 : _GEN_3231; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3233 = 6'h21 == select_50 ? io_inData_33 : _GEN_3232; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3234 = 6'h22 == select_50 ? io_inData_34 : _GEN_3233; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3235 = 6'h23 == select_50 ? io_inData_35 : _GEN_3234; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3236 = 6'h24 == select_50 ? io_inData_36 : _GEN_3235; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3237 = 6'h25 == select_50 ? io_inData_37 : _GEN_3236; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3238 = 6'h26 == select_50 ? io_inData_38 : _GEN_3237; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3239 = 6'h27 == select_50 ? io_inData_39 : _GEN_3238; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3240 = 6'h28 == select_50 ? io_inData_40 : _GEN_3239; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3241 = 6'h29 == select_50 ? io_inData_41 : _GEN_3240; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3242 = 6'h2a == select_50 ? io_inData_42 : _GEN_3241; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3243 = 6'h2b == select_50 ? io_inData_43 : _GEN_3242; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3244 = 6'h2c == select_50 ? io_inData_44 : _GEN_3243; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3245 = 6'h2d == select_50 ? io_inData_45 : _GEN_3244; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3246 = 6'h2e == select_50 ? io_inData_46 : _GEN_3245; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3247 = 6'h2f == select_50 ? io_inData_47 : _GEN_3246; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3248 = 6'h30 == select_50 ? io_inData_48 : _GEN_3247; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3249 = 6'h31 == select_50 ? io_inData_49 : _GEN_3248; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3250 = 6'h32 == select_50 ? io_inData_50 : _GEN_3249; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3251 = 6'h33 == select_50 ? io_inData_51 : _GEN_3250; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3252 = 6'h34 == select_50 ? io_inData_52 : _GEN_3251; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3253 = 6'h35 == select_50 ? io_inData_53 : _GEN_3252; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3254 = 6'h36 == select_50 ? io_inData_54 : _GEN_3253; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3255 = 6'h37 == select_50 ? io_inData_55 : _GEN_3254; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3256 = 6'h38 == select_50 ? io_inData_56 : _GEN_3255; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3257 = 6'h39 == select_50 ? io_inData_57 : _GEN_3256; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3258 = 6'h3a == select_50 ? io_inData_58 : _GEN_3257; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3259 = 6'h3b == select_50 ? io_inData_59 : _GEN_3258; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3260 = 6'h3c == select_50 ? io_inData_60 : _GEN_3259; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3261 = 6'h3d == select_50 ? io_inData_61 : _GEN_3260; // @[Switch.scala 33:19:@16366.4]
  assign _GEN_3262 = 6'h3e == select_50 ? io_inData_62 : _GEN_3261; // @[Switch.scala 33:19:@16366.4]
  assign _T_37229 = {valid_50_7,valid_50_6,valid_50_5,valid_50_4,valid_50_3,valid_50_2,valid_50_1,valid_50_0}; // @[Switch.scala 34:32:@16373.4]
  assign _T_37237 = {valid_50_15,valid_50_14,valid_50_13,valid_50_12,valid_50_11,valid_50_10,valid_50_9,valid_50_8,_T_37229}; // @[Switch.scala 34:32:@16381.4]
  assign _T_37244 = {valid_50_23,valid_50_22,valid_50_21,valid_50_20,valid_50_19,valid_50_18,valid_50_17,valid_50_16}; // @[Switch.scala 34:32:@16388.4]
  assign _T_37253 = {valid_50_31,valid_50_30,valid_50_29,valid_50_28,valid_50_27,valid_50_26,valid_50_25,valid_50_24,_T_37244,_T_37237}; // @[Switch.scala 34:32:@16397.4]
  assign _T_37260 = {valid_50_39,valid_50_38,valid_50_37,valid_50_36,valid_50_35,valid_50_34,valid_50_33,valid_50_32}; // @[Switch.scala 34:32:@16404.4]
  assign _T_37268 = {valid_50_47,valid_50_46,valid_50_45,valid_50_44,valid_50_43,valid_50_42,valid_50_41,valid_50_40,_T_37260}; // @[Switch.scala 34:32:@16412.4]
  assign _T_37275 = {valid_50_55,valid_50_54,valid_50_53,valid_50_52,valid_50_51,valid_50_50,valid_50_49,valid_50_48}; // @[Switch.scala 34:32:@16419.4]
  assign _T_37284 = {valid_50_63,valid_50_62,valid_50_61,valid_50_60,valid_50_59,valid_50_58,valid_50_57,valid_50_56,_T_37275,_T_37268}; // @[Switch.scala 34:32:@16428.4]
  assign _T_37285 = {_T_37284,_T_37253}; // @[Switch.scala 34:32:@16429.4]
  assign _T_37289 = io_inAddr_0 == 6'h33; // @[Switch.scala 30:53:@16432.4]
  assign valid_51_0 = io_inValid_0 & _T_37289; // @[Switch.scala 30:36:@16433.4]
  assign _T_37292 = io_inAddr_1 == 6'h33; // @[Switch.scala 30:53:@16435.4]
  assign valid_51_1 = io_inValid_1 & _T_37292; // @[Switch.scala 30:36:@16436.4]
  assign _T_37295 = io_inAddr_2 == 6'h33; // @[Switch.scala 30:53:@16438.4]
  assign valid_51_2 = io_inValid_2 & _T_37295; // @[Switch.scala 30:36:@16439.4]
  assign _T_37298 = io_inAddr_3 == 6'h33; // @[Switch.scala 30:53:@16441.4]
  assign valid_51_3 = io_inValid_3 & _T_37298; // @[Switch.scala 30:36:@16442.4]
  assign _T_37301 = io_inAddr_4 == 6'h33; // @[Switch.scala 30:53:@16444.4]
  assign valid_51_4 = io_inValid_4 & _T_37301; // @[Switch.scala 30:36:@16445.4]
  assign _T_37304 = io_inAddr_5 == 6'h33; // @[Switch.scala 30:53:@16447.4]
  assign valid_51_5 = io_inValid_5 & _T_37304; // @[Switch.scala 30:36:@16448.4]
  assign _T_37307 = io_inAddr_6 == 6'h33; // @[Switch.scala 30:53:@16450.4]
  assign valid_51_6 = io_inValid_6 & _T_37307; // @[Switch.scala 30:36:@16451.4]
  assign _T_37310 = io_inAddr_7 == 6'h33; // @[Switch.scala 30:53:@16453.4]
  assign valid_51_7 = io_inValid_7 & _T_37310; // @[Switch.scala 30:36:@16454.4]
  assign _T_37313 = io_inAddr_8 == 6'h33; // @[Switch.scala 30:53:@16456.4]
  assign valid_51_8 = io_inValid_8 & _T_37313; // @[Switch.scala 30:36:@16457.4]
  assign _T_37316 = io_inAddr_9 == 6'h33; // @[Switch.scala 30:53:@16459.4]
  assign valid_51_9 = io_inValid_9 & _T_37316; // @[Switch.scala 30:36:@16460.4]
  assign _T_37319 = io_inAddr_10 == 6'h33; // @[Switch.scala 30:53:@16462.4]
  assign valid_51_10 = io_inValid_10 & _T_37319; // @[Switch.scala 30:36:@16463.4]
  assign _T_37322 = io_inAddr_11 == 6'h33; // @[Switch.scala 30:53:@16465.4]
  assign valid_51_11 = io_inValid_11 & _T_37322; // @[Switch.scala 30:36:@16466.4]
  assign _T_37325 = io_inAddr_12 == 6'h33; // @[Switch.scala 30:53:@16468.4]
  assign valid_51_12 = io_inValid_12 & _T_37325; // @[Switch.scala 30:36:@16469.4]
  assign _T_37328 = io_inAddr_13 == 6'h33; // @[Switch.scala 30:53:@16471.4]
  assign valid_51_13 = io_inValid_13 & _T_37328; // @[Switch.scala 30:36:@16472.4]
  assign _T_37331 = io_inAddr_14 == 6'h33; // @[Switch.scala 30:53:@16474.4]
  assign valid_51_14 = io_inValid_14 & _T_37331; // @[Switch.scala 30:36:@16475.4]
  assign _T_37334 = io_inAddr_15 == 6'h33; // @[Switch.scala 30:53:@16477.4]
  assign valid_51_15 = io_inValid_15 & _T_37334; // @[Switch.scala 30:36:@16478.4]
  assign _T_37337 = io_inAddr_16 == 6'h33; // @[Switch.scala 30:53:@16480.4]
  assign valid_51_16 = io_inValid_16 & _T_37337; // @[Switch.scala 30:36:@16481.4]
  assign _T_37340 = io_inAddr_17 == 6'h33; // @[Switch.scala 30:53:@16483.4]
  assign valid_51_17 = io_inValid_17 & _T_37340; // @[Switch.scala 30:36:@16484.4]
  assign _T_37343 = io_inAddr_18 == 6'h33; // @[Switch.scala 30:53:@16486.4]
  assign valid_51_18 = io_inValid_18 & _T_37343; // @[Switch.scala 30:36:@16487.4]
  assign _T_37346 = io_inAddr_19 == 6'h33; // @[Switch.scala 30:53:@16489.4]
  assign valid_51_19 = io_inValid_19 & _T_37346; // @[Switch.scala 30:36:@16490.4]
  assign _T_37349 = io_inAddr_20 == 6'h33; // @[Switch.scala 30:53:@16492.4]
  assign valid_51_20 = io_inValid_20 & _T_37349; // @[Switch.scala 30:36:@16493.4]
  assign _T_37352 = io_inAddr_21 == 6'h33; // @[Switch.scala 30:53:@16495.4]
  assign valid_51_21 = io_inValid_21 & _T_37352; // @[Switch.scala 30:36:@16496.4]
  assign _T_37355 = io_inAddr_22 == 6'h33; // @[Switch.scala 30:53:@16498.4]
  assign valid_51_22 = io_inValid_22 & _T_37355; // @[Switch.scala 30:36:@16499.4]
  assign _T_37358 = io_inAddr_23 == 6'h33; // @[Switch.scala 30:53:@16501.4]
  assign valid_51_23 = io_inValid_23 & _T_37358; // @[Switch.scala 30:36:@16502.4]
  assign _T_37361 = io_inAddr_24 == 6'h33; // @[Switch.scala 30:53:@16504.4]
  assign valid_51_24 = io_inValid_24 & _T_37361; // @[Switch.scala 30:36:@16505.4]
  assign _T_37364 = io_inAddr_25 == 6'h33; // @[Switch.scala 30:53:@16507.4]
  assign valid_51_25 = io_inValid_25 & _T_37364; // @[Switch.scala 30:36:@16508.4]
  assign _T_37367 = io_inAddr_26 == 6'h33; // @[Switch.scala 30:53:@16510.4]
  assign valid_51_26 = io_inValid_26 & _T_37367; // @[Switch.scala 30:36:@16511.4]
  assign _T_37370 = io_inAddr_27 == 6'h33; // @[Switch.scala 30:53:@16513.4]
  assign valid_51_27 = io_inValid_27 & _T_37370; // @[Switch.scala 30:36:@16514.4]
  assign _T_37373 = io_inAddr_28 == 6'h33; // @[Switch.scala 30:53:@16516.4]
  assign valid_51_28 = io_inValid_28 & _T_37373; // @[Switch.scala 30:36:@16517.4]
  assign _T_37376 = io_inAddr_29 == 6'h33; // @[Switch.scala 30:53:@16519.4]
  assign valid_51_29 = io_inValid_29 & _T_37376; // @[Switch.scala 30:36:@16520.4]
  assign _T_37379 = io_inAddr_30 == 6'h33; // @[Switch.scala 30:53:@16522.4]
  assign valid_51_30 = io_inValid_30 & _T_37379; // @[Switch.scala 30:36:@16523.4]
  assign _T_37382 = io_inAddr_31 == 6'h33; // @[Switch.scala 30:53:@16525.4]
  assign valid_51_31 = io_inValid_31 & _T_37382; // @[Switch.scala 30:36:@16526.4]
  assign _T_37385 = io_inAddr_32 == 6'h33; // @[Switch.scala 30:53:@16528.4]
  assign valid_51_32 = io_inValid_32 & _T_37385; // @[Switch.scala 30:36:@16529.4]
  assign _T_37388 = io_inAddr_33 == 6'h33; // @[Switch.scala 30:53:@16531.4]
  assign valid_51_33 = io_inValid_33 & _T_37388; // @[Switch.scala 30:36:@16532.4]
  assign _T_37391 = io_inAddr_34 == 6'h33; // @[Switch.scala 30:53:@16534.4]
  assign valid_51_34 = io_inValid_34 & _T_37391; // @[Switch.scala 30:36:@16535.4]
  assign _T_37394 = io_inAddr_35 == 6'h33; // @[Switch.scala 30:53:@16537.4]
  assign valid_51_35 = io_inValid_35 & _T_37394; // @[Switch.scala 30:36:@16538.4]
  assign _T_37397 = io_inAddr_36 == 6'h33; // @[Switch.scala 30:53:@16540.4]
  assign valid_51_36 = io_inValid_36 & _T_37397; // @[Switch.scala 30:36:@16541.4]
  assign _T_37400 = io_inAddr_37 == 6'h33; // @[Switch.scala 30:53:@16543.4]
  assign valid_51_37 = io_inValid_37 & _T_37400; // @[Switch.scala 30:36:@16544.4]
  assign _T_37403 = io_inAddr_38 == 6'h33; // @[Switch.scala 30:53:@16546.4]
  assign valid_51_38 = io_inValid_38 & _T_37403; // @[Switch.scala 30:36:@16547.4]
  assign _T_37406 = io_inAddr_39 == 6'h33; // @[Switch.scala 30:53:@16549.4]
  assign valid_51_39 = io_inValid_39 & _T_37406; // @[Switch.scala 30:36:@16550.4]
  assign _T_37409 = io_inAddr_40 == 6'h33; // @[Switch.scala 30:53:@16552.4]
  assign valid_51_40 = io_inValid_40 & _T_37409; // @[Switch.scala 30:36:@16553.4]
  assign _T_37412 = io_inAddr_41 == 6'h33; // @[Switch.scala 30:53:@16555.4]
  assign valid_51_41 = io_inValid_41 & _T_37412; // @[Switch.scala 30:36:@16556.4]
  assign _T_37415 = io_inAddr_42 == 6'h33; // @[Switch.scala 30:53:@16558.4]
  assign valid_51_42 = io_inValid_42 & _T_37415; // @[Switch.scala 30:36:@16559.4]
  assign _T_37418 = io_inAddr_43 == 6'h33; // @[Switch.scala 30:53:@16561.4]
  assign valid_51_43 = io_inValid_43 & _T_37418; // @[Switch.scala 30:36:@16562.4]
  assign _T_37421 = io_inAddr_44 == 6'h33; // @[Switch.scala 30:53:@16564.4]
  assign valid_51_44 = io_inValid_44 & _T_37421; // @[Switch.scala 30:36:@16565.4]
  assign _T_37424 = io_inAddr_45 == 6'h33; // @[Switch.scala 30:53:@16567.4]
  assign valid_51_45 = io_inValid_45 & _T_37424; // @[Switch.scala 30:36:@16568.4]
  assign _T_37427 = io_inAddr_46 == 6'h33; // @[Switch.scala 30:53:@16570.4]
  assign valid_51_46 = io_inValid_46 & _T_37427; // @[Switch.scala 30:36:@16571.4]
  assign _T_37430 = io_inAddr_47 == 6'h33; // @[Switch.scala 30:53:@16573.4]
  assign valid_51_47 = io_inValid_47 & _T_37430; // @[Switch.scala 30:36:@16574.4]
  assign _T_37433 = io_inAddr_48 == 6'h33; // @[Switch.scala 30:53:@16576.4]
  assign valid_51_48 = io_inValid_48 & _T_37433; // @[Switch.scala 30:36:@16577.4]
  assign _T_37436 = io_inAddr_49 == 6'h33; // @[Switch.scala 30:53:@16579.4]
  assign valid_51_49 = io_inValid_49 & _T_37436; // @[Switch.scala 30:36:@16580.4]
  assign _T_37439 = io_inAddr_50 == 6'h33; // @[Switch.scala 30:53:@16582.4]
  assign valid_51_50 = io_inValid_50 & _T_37439; // @[Switch.scala 30:36:@16583.4]
  assign _T_37442 = io_inAddr_51 == 6'h33; // @[Switch.scala 30:53:@16585.4]
  assign valid_51_51 = io_inValid_51 & _T_37442; // @[Switch.scala 30:36:@16586.4]
  assign _T_37445 = io_inAddr_52 == 6'h33; // @[Switch.scala 30:53:@16588.4]
  assign valid_51_52 = io_inValid_52 & _T_37445; // @[Switch.scala 30:36:@16589.4]
  assign _T_37448 = io_inAddr_53 == 6'h33; // @[Switch.scala 30:53:@16591.4]
  assign valid_51_53 = io_inValid_53 & _T_37448; // @[Switch.scala 30:36:@16592.4]
  assign _T_37451 = io_inAddr_54 == 6'h33; // @[Switch.scala 30:53:@16594.4]
  assign valid_51_54 = io_inValid_54 & _T_37451; // @[Switch.scala 30:36:@16595.4]
  assign _T_37454 = io_inAddr_55 == 6'h33; // @[Switch.scala 30:53:@16597.4]
  assign valid_51_55 = io_inValid_55 & _T_37454; // @[Switch.scala 30:36:@16598.4]
  assign _T_37457 = io_inAddr_56 == 6'h33; // @[Switch.scala 30:53:@16600.4]
  assign valid_51_56 = io_inValid_56 & _T_37457; // @[Switch.scala 30:36:@16601.4]
  assign _T_37460 = io_inAddr_57 == 6'h33; // @[Switch.scala 30:53:@16603.4]
  assign valid_51_57 = io_inValid_57 & _T_37460; // @[Switch.scala 30:36:@16604.4]
  assign _T_37463 = io_inAddr_58 == 6'h33; // @[Switch.scala 30:53:@16606.4]
  assign valid_51_58 = io_inValid_58 & _T_37463; // @[Switch.scala 30:36:@16607.4]
  assign _T_37466 = io_inAddr_59 == 6'h33; // @[Switch.scala 30:53:@16609.4]
  assign valid_51_59 = io_inValid_59 & _T_37466; // @[Switch.scala 30:36:@16610.4]
  assign _T_37469 = io_inAddr_60 == 6'h33; // @[Switch.scala 30:53:@16612.4]
  assign valid_51_60 = io_inValid_60 & _T_37469; // @[Switch.scala 30:36:@16613.4]
  assign _T_37472 = io_inAddr_61 == 6'h33; // @[Switch.scala 30:53:@16615.4]
  assign valid_51_61 = io_inValid_61 & _T_37472; // @[Switch.scala 30:36:@16616.4]
  assign _T_37475 = io_inAddr_62 == 6'h33; // @[Switch.scala 30:53:@16618.4]
  assign valid_51_62 = io_inValid_62 & _T_37475; // @[Switch.scala 30:36:@16619.4]
  assign _T_37478 = io_inAddr_63 == 6'h33; // @[Switch.scala 30:53:@16621.4]
  assign valid_51_63 = io_inValid_63 & _T_37478; // @[Switch.scala 30:36:@16622.4]
  assign _T_37544 = valid_51_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@16624.4]
  assign _T_37545 = valid_51_61 ? 6'h3d : _T_37544; // @[Mux.scala 31:69:@16625.4]
  assign _T_37546 = valid_51_60 ? 6'h3c : _T_37545; // @[Mux.scala 31:69:@16626.4]
  assign _T_37547 = valid_51_59 ? 6'h3b : _T_37546; // @[Mux.scala 31:69:@16627.4]
  assign _T_37548 = valid_51_58 ? 6'h3a : _T_37547; // @[Mux.scala 31:69:@16628.4]
  assign _T_37549 = valid_51_57 ? 6'h39 : _T_37548; // @[Mux.scala 31:69:@16629.4]
  assign _T_37550 = valid_51_56 ? 6'h38 : _T_37549; // @[Mux.scala 31:69:@16630.4]
  assign _T_37551 = valid_51_55 ? 6'h37 : _T_37550; // @[Mux.scala 31:69:@16631.4]
  assign _T_37552 = valid_51_54 ? 6'h36 : _T_37551; // @[Mux.scala 31:69:@16632.4]
  assign _T_37553 = valid_51_53 ? 6'h35 : _T_37552; // @[Mux.scala 31:69:@16633.4]
  assign _T_37554 = valid_51_52 ? 6'h34 : _T_37553; // @[Mux.scala 31:69:@16634.4]
  assign _T_37555 = valid_51_51 ? 6'h33 : _T_37554; // @[Mux.scala 31:69:@16635.4]
  assign _T_37556 = valid_51_50 ? 6'h32 : _T_37555; // @[Mux.scala 31:69:@16636.4]
  assign _T_37557 = valid_51_49 ? 6'h31 : _T_37556; // @[Mux.scala 31:69:@16637.4]
  assign _T_37558 = valid_51_48 ? 6'h30 : _T_37557; // @[Mux.scala 31:69:@16638.4]
  assign _T_37559 = valid_51_47 ? 6'h2f : _T_37558; // @[Mux.scala 31:69:@16639.4]
  assign _T_37560 = valid_51_46 ? 6'h2e : _T_37559; // @[Mux.scala 31:69:@16640.4]
  assign _T_37561 = valid_51_45 ? 6'h2d : _T_37560; // @[Mux.scala 31:69:@16641.4]
  assign _T_37562 = valid_51_44 ? 6'h2c : _T_37561; // @[Mux.scala 31:69:@16642.4]
  assign _T_37563 = valid_51_43 ? 6'h2b : _T_37562; // @[Mux.scala 31:69:@16643.4]
  assign _T_37564 = valid_51_42 ? 6'h2a : _T_37563; // @[Mux.scala 31:69:@16644.4]
  assign _T_37565 = valid_51_41 ? 6'h29 : _T_37564; // @[Mux.scala 31:69:@16645.4]
  assign _T_37566 = valid_51_40 ? 6'h28 : _T_37565; // @[Mux.scala 31:69:@16646.4]
  assign _T_37567 = valid_51_39 ? 6'h27 : _T_37566; // @[Mux.scala 31:69:@16647.4]
  assign _T_37568 = valid_51_38 ? 6'h26 : _T_37567; // @[Mux.scala 31:69:@16648.4]
  assign _T_37569 = valid_51_37 ? 6'h25 : _T_37568; // @[Mux.scala 31:69:@16649.4]
  assign _T_37570 = valid_51_36 ? 6'h24 : _T_37569; // @[Mux.scala 31:69:@16650.4]
  assign _T_37571 = valid_51_35 ? 6'h23 : _T_37570; // @[Mux.scala 31:69:@16651.4]
  assign _T_37572 = valid_51_34 ? 6'h22 : _T_37571; // @[Mux.scala 31:69:@16652.4]
  assign _T_37573 = valid_51_33 ? 6'h21 : _T_37572; // @[Mux.scala 31:69:@16653.4]
  assign _T_37574 = valid_51_32 ? 6'h20 : _T_37573; // @[Mux.scala 31:69:@16654.4]
  assign _T_37575 = valid_51_31 ? 6'h1f : _T_37574; // @[Mux.scala 31:69:@16655.4]
  assign _T_37576 = valid_51_30 ? 6'h1e : _T_37575; // @[Mux.scala 31:69:@16656.4]
  assign _T_37577 = valid_51_29 ? 6'h1d : _T_37576; // @[Mux.scala 31:69:@16657.4]
  assign _T_37578 = valid_51_28 ? 6'h1c : _T_37577; // @[Mux.scala 31:69:@16658.4]
  assign _T_37579 = valid_51_27 ? 6'h1b : _T_37578; // @[Mux.scala 31:69:@16659.4]
  assign _T_37580 = valid_51_26 ? 6'h1a : _T_37579; // @[Mux.scala 31:69:@16660.4]
  assign _T_37581 = valid_51_25 ? 6'h19 : _T_37580; // @[Mux.scala 31:69:@16661.4]
  assign _T_37582 = valid_51_24 ? 6'h18 : _T_37581; // @[Mux.scala 31:69:@16662.4]
  assign _T_37583 = valid_51_23 ? 6'h17 : _T_37582; // @[Mux.scala 31:69:@16663.4]
  assign _T_37584 = valid_51_22 ? 6'h16 : _T_37583; // @[Mux.scala 31:69:@16664.4]
  assign _T_37585 = valid_51_21 ? 6'h15 : _T_37584; // @[Mux.scala 31:69:@16665.4]
  assign _T_37586 = valid_51_20 ? 6'h14 : _T_37585; // @[Mux.scala 31:69:@16666.4]
  assign _T_37587 = valid_51_19 ? 6'h13 : _T_37586; // @[Mux.scala 31:69:@16667.4]
  assign _T_37588 = valid_51_18 ? 6'h12 : _T_37587; // @[Mux.scala 31:69:@16668.4]
  assign _T_37589 = valid_51_17 ? 6'h11 : _T_37588; // @[Mux.scala 31:69:@16669.4]
  assign _T_37590 = valid_51_16 ? 6'h10 : _T_37589; // @[Mux.scala 31:69:@16670.4]
  assign _T_37591 = valid_51_15 ? 6'hf : _T_37590; // @[Mux.scala 31:69:@16671.4]
  assign _T_37592 = valid_51_14 ? 6'he : _T_37591; // @[Mux.scala 31:69:@16672.4]
  assign _T_37593 = valid_51_13 ? 6'hd : _T_37592; // @[Mux.scala 31:69:@16673.4]
  assign _T_37594 = valid_51_12 ? 6'hc : _T_37593; // @[Mux.scala 31:69:@16674.4]
  assign _T_37595 = valid_51_11 ? 6'hb : _T_37594; // @[Mux.scala 31:69:@16675.4]
  assign _T_37596 = valid_51_10 ? 6'ha : _T_37595; // @[Mux.scala 31:69:@16676.4]
  assign _T_37597 = valid_51_9 ? 6'h9 : _T_37596; // @[Mux.scala 31:69:@16677.4]
  assign _T_37598 = valid_51_8 ? 6'h8 : _T_37597; // @[Mux.scala 31:69:@16678.4]
  assign _T_37599 = valid_51_7 ? 6'h7 : _T_37598; // @[Mux.scala 31:69:@16679.4]
  assign _T_37600 = valid_51_6 ? 6'h6 : _T_37599; // @[Mux.scala 31:69:@16680.4]
  assign _T_37601 = valid_51_5 ? 6'h5 : _T_37600; // @[Mux.scala 31:69:@16681.4]
  assign _T_37602 = valid_51_4 ? 6'h4 : _T_37601; // @[Mux.scala 31:69:@16682.4]
  assign _T_37603 = valid_51_3 ? 6'h3 : _T_37602; // @[Mux.scala 31:69:@16683.4]
  assign _T_37604 = valid_51_2 ? 6'h2 : _T_37603; // @[Mux.scala 31:69:@16684.4]
  assign _T_37605 = valid_51_1 ? 6'h1 : _T_37604; // @[Mux.scala 31:69:@16685.4]
  assign select_51 = valid_51_0 ? 6'h0 : _T_37605; // @[Mux.scala 31:69:@16686.4]
  assign _GEN_3265 = 6'h1 == select_51 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3266 = 6'h2 == select_51 ? io_inData_2 : _GEN_3265; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3267 = 6'h3 == select_51 ? io_inData_3 : _GEN_3266; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3268 = 6'h4 == select_51 ? io_inData_4 : _GEN_3267; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3269 = 6'h5 == select_51 ? io_inData_5 : _GEN_3268; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3270 = 6'h6 == select_51 ? io_inData_6 : _GEN_3269; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3271 = 6'h7 == select_51 ? io_inData_7 : _GEN_3270; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3272 = 6'h8 == select_51 ? io_inData_8 : _GEN_3271; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3273 = 6'h9 == select_51 ? io_inData_9 : _GEN_3272; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3274 = 6'ha == select_51 ? io_inData_10 : _GEN_3273; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3275 = 6'hb == select_51 ? io_inData_11 : _GEN_3274; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3276 = 6'hc == select_51 ? io_inData_12 : _GEN_3275; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3277 = 6'hd == select_51 ? io_inData_13 : _GEN_3276; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3278 = 6'he == select_51 ? io_inData_14 : _GEN_3277; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3279 = 6'hf == select_51 ? io_inData_15 : _GEN_3278; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3280 = 6'h10 == select_51 ? io_inData_16 : _GEN_3279; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3281 = 6'h11 == select_51 ? io_inData_17 : _GEN_3280; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3282 = 6'h12 == select_51 ? io_inData_18 : _GEN_3281; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3283 = 6'h13 == select_51 ? io_inData_19 : _GEN_3282; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3284 = 6'h14 == select_51 ? io_inData_20 : _GEN_3283; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3285 = 6'h15 == select_51 ? io_inData_21 : _GEN_3284; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3286 = 6'h16 == select_51 ? io_inData_22 : _GEN_3285; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3287 = 6'h17 == select_51 ? io_inData_23 : _GEN_3286; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3288 = 6'h18 == select_51 ? io_inData_24 : _GEN_3287; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3289 = 6'h19 == select_51 ? io_inData_25 : _GEN_3288; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3290 = 6'h1a == select_51 ? io_inData_26 : _GEN_3289; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3291 = 6'h1b == select_51 ? io_inData_27 : _GEN_3290; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3292 = 6'h1c == select_51 ? io_inData_28 : _GEN_3291; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3293 = 6'h1d == select_51 ? io_inData_29 : _GEN_3292; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3294 = 6'h1e == select_51 ? io_inData_30 : _GEN_3293; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3295 = 6'h1f == select_51 ? io_inData_31 : _GEN_3294; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3296 = 6'h20 == select_51 ? io_inData_32 : _GEN_3295; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3297 = 6'h21 == select_51 ? io_inData_33 : _GEN_3296; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3298 = 6'h22 == select_51 ? io_inData_34 : _GEN_3297; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3299 = 6'h23 == select_51 ? io_inData_35 : _GEN_3298; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3300 = 6'h24 == select_51 ? io_inData_36 : _GEN_3299; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3301 = 6'h25 == select_51 ? io_inData_37 : _GEN_3300; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3302 = 6'h26 == select_51 ? io_inData_38 : _GEN_3301; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3303 = 6'h27 == select_51 ? io_inData_39 : _GEN_3302; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3304 = 6'h28 == select_51 ? io_inData_40 : _GEN_3303; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3305 = 6'h29 == select_51 ? io_inData_41 : _GEN_3304; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3306 = 6'h2a == select_51 ? io_inData_42 : _GEN_3305; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3307 = 6'h2b == select_51 ? io_inData_43 : _GEN_3306; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3308 = 6'h2c == select_51 ? io_inData_44 : _GEN_3307; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3309 = 6'h2d == select_51 ? io_inData_45 : _GEN_3308; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3310 = 6'h2e == select_51 ? io_inData_46 : _GEN_3309; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3311 = 6'h2f == select_51 ? io_inData_47 : _GEN_3310; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3312 = 6'h30 == select_51 ? io_inData_48 : _GEN_3311; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3313 = 6'h31 == select_51 ? io_inData_49 : _GEN_3312; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3314 = 6'h32 == select_51 ? io_inData_50 : _GEN_3313; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3315 = 6'h33 == select_51 ? io_inData_51 : _GEN_3314; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3316 = 6'h34 == select_51 ? io_inData_52 : _GEN_3315; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3317 = 6'h35 == select_51 ? io_inData_53 : _GEN_3316; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3318 = 6'h36 == select_51 ? io_inData_54 : _GEN_3317; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3319 = 6'h37 == select_51 ? io_inData_55 : _GEN_3318; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3320 = 6'h38 == select_51 ? io_inData_56 : _GEN_3319; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3321 = 6'h39 == select_51 ? io_inData_57 : _GEN_3320; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3322 = 6'h3a == select_51 ? io_inData_58 : _GEN_3321; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3323 = 6'h3b == select_51 ? io_inData_59 : _GEN_3322; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3324 = 6'h3c == select_51 ? io_inData_60 : _GEN_3323; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3325 = 6'h3d == select_51 ? io_inData_61 : _GEN_3324; // @[Switch.scala 33:19:@16688.4]
  assign _GEN_3326 = 6'h3e == select_51 ? io_inData_62 : _GEN_3325; // @[Switch.scala 33:19:@16688.4]
  assign _T_37614 = {valid_51_7,valid_51_6,valid_51_5,valid_51_4,valid_51_3,valid_51_2,valid_51_1,valid_51_0}; // @[Switch.scala 34:32:@16695.4]
  assign _T_37622 = {valid_51_15,valid_51_14,valid_51_13,valid_51_12,valid_51_11,valid_51_10,valid_51_9,valid_51_8,_T_37614}; // @[Switch.scala 34:32:@16703.4]
  assign _T_37629 = {valid_51_23,valid_51_22,valid_51_21,valid_51_20,valid_51_19,valid_51_18,valid_51_17,valid_51_16}; // @[Switch.scala 34:32:@16710.4]
  assign _T_37638 = {valid_51_31,valid_51_30,valid_51_29,valid_51_28,valid_51_27,valid_51_26,valid_51_25,valid_51_24,_T_37629,_T_37622}; // @[Switch.scala 34:32:@16719.4]
  assign _T_37645 = {valid_51_39,valid_51_38,valid_51_37,valid_51_36,valid_51_35,valid_51_34,valid_51_33,valid_51_32}; // @[Switch.scala 34:32:@16726.4]
  assign _T_37653 = {valid_51_47,valid_51_46,valid_51_45,valid_51_44,valid_51_43,valid_51_42,valid_51_41,valid_51_40,_T_37645}; // @[Switch.scala 34:32:@16734.4]
  assign _T_37660 = {valid_51_55,valid_51_54,valid_51_53,valid_51_52,valid_51_51,valid_51_50,valid_51_49,valid_51_48}; // @[Switch.scala 34:32:@16741.4]
  assign _T_37669 = {valid_51_63,valid_51_62,valid_51_61,valid_51_60,valid_51_59,valid_51_58,valid_51_57,valid_51_56,_T_37660,_T_37653}; // @[Switch.scala 34:32:@16750.4]
  assign _T_37670 = {_T_37669,_T_37638}; // @[Switch.scala 34:32:@16751.4]
  assign _T_37674 = io_inAddr_0 == 6'h34; // @[Switch.scala 30:53:@16754.4]
  assign valid_52_0 = io_inValid_0 & _T_37674; // @[Switch.scala 30:36:@16755.4]
  assign _T_37677 = io_inAddr_1 == 6'h34; // @[Switch.scala 30:53:@16757.4]
  assign valid_52_1 = io_inValid_1 & _T_37677; // @[Switch.scala 30:36:@16758.4]
  assign _T_37680 = io_inAddr_2 == 6'h34; // @[Switch.scala 30:53:@16760.4]
  assign valid_52_2 = io_inValid_2 & _T_37680; // @[Switch.scala 30:36:@16761.4]
  assign _T_37683 = io_inAddr_3 == 6'h34; // @[Switch.scala 30:53:@16763.4]
  assign valid_52_3 = io_inValid_3 & _T_37683; // @[Switch.scala 30:36:@16764.4]
  assign _T_37686 = io_inAddr_4 == 6'h34; // @[Switch.scala 30:53:@16766.4]
  assign valid_52_4 = io_inValid_4 & _T_37686; // @[Switch.scala 30:36:@16767.4]
  assign _T_37689 = io_inAddr_5 == 6'h34; // @[Switch.scala 30:53:@16769.4]
  assign valid_52_5 = io_inValid_5 & _T_37689; // @[Switch.scala 30:36:@16770.4]
  assign _T_37692 = io_inAddr_6 == 6'h34; // @[Switch.scala 30:53:@16772.4]
  assign valid_52_6 = io_inValid_6 & _T_37692; // @[Switch.scala 30:36:@16773.4]
  assign _T_37695 = io_inAddr_7 == 6'h34; // @[Switch.scala 30:53:@16775.4]
  assign valid_52_7 = io_inValid_7 & _T_37695; // @[Switch.scala 30:36:@16776.4]
  assign _T_37698 = io_inAddr_8 == 6'h34; // @[Switch.scala 30:53:@16778.4]
  assign valid_52_8 = io_inValid_8 & _T_37698; // @[Switch.scala 30:36:@16779.4]
  assign _T_37701 = io_inAddr_9 == 6'h34; // @[Switch.scala 30:53:@16781.4]
  assign valid_52_9 = io_inValid_9 & _T_37701; // @[Switch.scala 30:36:@16782.4]
  assign _T_37704 = io_inAddr_10 == 6'h34; // @[Switch.scala 30:53:@16784.4]
  assign valid_52_10 = io_inValid_10 & _T_37704; // @[Switch.scala 30:36:@16785.4]
  assign _T_37707 = io_inAddr_11 == 6'h34; // @[Switch.scala 30:53:@16787.4]
  assign valid_52_11 = io_inValid_11 & _T_37707; // @[Switch.scala 30:36:@16788.4]
  assign _T_37710 = io_inAddr_12 == 6'h34; // @[Switch.scala 30:53:@16790.4]
  assign valid_52_12 = io_inValid_12 & _T_37710; // @[Switch.scala 30:36:@16791.4]
  assign _T_37713 = io_inAddr_13 == 6'h34; // @[Switch.scala 30:53:@16793.4]
  assign valid_52_13 = io_inValid_13 & _T_37713; // @[Switch.scala 30:36:@16794.4]
  assign _T_37716 = io_inAddr_14 == 6'h34; // @[Switch.scala 30:53:@16796.4]
  assign valid_52_14 = io_inValid_14 & _T_37716; // @[Switch.scala 30:36:@16797.4]
  assign _T_37719 = io_inAddr_15 == 6'h34; // @[Switch.scala 30:53:@16799.4]
  assign valid_52_15 = io_inValid_15 & _T_37719; // @[Switch.scala 30:36:@16800.4]
  assign _T_37722 = io_inAddr_16 == 6'h34; // @[Switch.scala 30:53:@16802.4]
  assign valid_52_16 = io_inValid_16 & _T_37722; // @[Switch.scala 30:36:@16803.4]
  assign _T_37725 = io_inAddr_17 == 6'h34; // @[Switch.scala 30:53:@16805.4]
  assign valid_52_17 = io_inValid_17 & _T_37725; // @[Switch.scala 30:36:@16806.4]
  assign _T_37728 = io_inAddr_18 == 6'h34; // @[Switch.scala 30:53:@16808.4]
  assign valid_52_18 = io_inValid_18 & _T_37728; // @[Switch.scala 30:36:@16809.4]
  assign _T_37731 = io_inAddr_19 == 6'h34; // @[Switch.scala 30:53:@16811.4]
  assign valid_52_19 = io_inValid_19 & _T_37731; // @[Switch.scala 30:36:@16812.4]
  assign _T_37734 = io_inAddr_20 == 6'h34; // @[Switch.scala 30:53:@16814.4]
  assign valid_52_20 = io_inValid_20 & _T_37734; // @[Switch.scala 30:36:@16815.4]
  assign _T_37737 = io_inAddr_21 == 6'h34; // @[Switch.scala 30:53:@16817.4]
  assign valid_52_21 = io_inValid_21 & _T_37737; // @[Switch.scala 30:36:@16818.4]
  assign _T_37740 = io_inAddr_22 == 6'h34; // @[Switch.scala 30:53:@16820.4]
  assign valid_52_22 = io_inValid_22 & _T_37740; // @[Switch.scala 30:36:@16821.4]
  assign _T_37743 = io_inAddr_23 == 6'h34; // @[Switch.scala 30:53:@16823.4]
  assign valid_52_23 = io_inValid_23 & _T_37743; // @[Switch.scala 30:36:@16824.4]
  assign _T_37746 = io_inAddr_24 == 6'h34; // @[Switch.scala 30:53:@16826.4]
  assign valid_52_24 = io_inValid_24 & _T_37746; // @[Switch.scala 30:36:@16827.4]
  assign _T_37749 = io_inAddr_25 == 6'h34; // @[Switch.scala 30:53:@16829.4]
  assign valid_52_25 = io_inValid_25 & _T_37749; // @[Switch.scala 30:36:@16830.4]
  assign _T_37752 = io_inAddr_26 == 6'h34; // @[Switch.scala 30:53:@16832.4]
  assign valid_52_26 = io_inValid_26 & _T_37752; // @[Switch.scala 30:36:@16833.4]
  assign _T_37755 = io_inAddr_27 == 6'h34; // @[Switch.scala 30:53:@16835.4]
  assign valid_52_27 = io_inValid_27 & _T_37755; // @[Switch.scala 30:36:@16836.4]
  assign _T_37758 = io_inAddr_28 == 6'h34; // @[Switch.scala 30:53:@16838.4]
  assign valid_52_28 = io_inValid_28 & _T_37758; // @[Switch.scala 30:36:@16839.4]
  assign _T_37761 = io_inAddr_29 == 6'h34; // @[Switch.scala 30:53:@16841.4]
  assign valid_52_29 = io_inValid_29 & _T_37761; // @[Switch.scala 30:36:@16842.4]
  assign _T_37764 = io_inAddr_30 == 6'h34; // @[Switch.scala 30:53:@16844.4]
  assign valid_52_30 = io_inValid_30 & _T_37764; // @[Switch.scala 30:36:@16845.4]
  assign _T_37767 = io_inAddr_31 == 6'h34; // @[Switch.scala 30:53:@16847.4]
  assign valid_52_31 = io_inValid_31 & _T_37767; // @[Switch.scala 30:36:@16848.4]
  assign _T_37770 = io_inAddr_32 == 6'h34; // @[Switch.scala 30:53:@16850.4]
  assign valid_52_32 = io_inValid_32 & _T_37770; // @[Switch.scala 30:36:@16851.4]
  assign _T_37773 = io_inAddr_33 == 6'h34; // @[Switch.scala 30:53:@16853.4]
  assign valid_52_33 = io_inValid_33 & _T_37773; // @[Switch.scala 30:36:@16854.4]
  assign _T_37776 = io_inAddr_34 == 6'h34; // @[Switch.scala 30:53:@16856.4]
  assign valid_52_34 = io_inValid_34 & _T_37776; // @[Switch.scala 30:36:@16857.4]
  assign _T_37779 = io_inAddr_35 == 6'h34; // @[Switch.scala 30:53:@16859.4]
  assign valid_52_35 = io_inValid_35 & _T_37779; // @[Switch.scala 30:36:@16860.4]
  assign _T_37782 = io_inAddr_36 == 6'h34; // @[Switch.scala 30:53:@16862.4]
  assign valid_52_36 = io_inValid_36 & _T_37782; // @[Switch.scala 30:36:@16863.4]
  assign _T_37785 = io_inAddr_37 == 6'h34; // @[Switch.scala 30:53:@16865.4]
  assign valid_52_37 = io_inValid_37 & _T_37785; // @[Switch.scala 30:36:@16866.4]
  assign _T_37788 = io_inAddr_38 == 6'h34; // @[Switch.scala 30:53:@16868.4]
  assign valid_52_38 = io_inValid_38 & _T_37788; // @[Switch.scala 30:36:@16869.4]
  assign _T_37791 = io_inAddr_39 == 6'h34; // @[Switch.scala 30:53:@16871.4]
  assign valid_52_39 = io_inValid_39 & _T_37791; // @[Switch.scala 30:36:@16872.4]
  assign _T_37794 = io_inAddr_40 == 6'h34; // @[Switch.scala 30:53:@16874.4]
  assign valid_52_40 = io_inValid_40 & _T_37794; // @[Switch.scala 30:36:@16875.4]
  assign _T_37797 = io_inAddr_41 == 6'h34; // @[Switch.scala 30:53:@16877.4]
  assign valid_52_41 = io_inValid_41 & _T_37797; // @[Switch.scala 30:36:@16878.4]
  assign _T_37800 = io_inAddr_42 == 6'h34; // @[Switch.scala 30:53:@16880.4]
  assign valid_52_42 = io_inValid_42 & _T_37800; // @[Switch.scala 30:36:@16881.4]
  assign _T_37803 = io_inAddr_43 == 6'h34; // @[Switch.scala 30:53:@16883.4]
  assign valid_52_43 = io_inValid_43 & _T_37803; // @[Switch.scala 30:36:@16884.4]
  assign _T_37806 = io_inAddr_44 == 6'h34; // @[Switch.scala 30:53:@16886.4]
  assign valid_52_44 = io_inValid_44 & _T_37806; // @[Switch.scala 30:36:@16887.4]
  assign _T_37809 = io_inAddr_45 == 6'h34; // @[Switch.scala 30:53:@16889.4]
  assign valid_52_45 = io_inValid_45 & _T_37809; // @[Switch.scala 30:36:@16890.4]
  assign _T_37812 = io_inAddr_46 == 6'h34; // @[Switch.scala 30:53:@16892.4]
  assign valid_52_46 = io_inValid_46 & _T_37812; // @[Switch.scala 30:36:@16893.4]
  assign _T_37815 = io_inAddr_47 == 6'h34; // @[Switch.scala 30:53:@16895.4]
  assign valid_52_47 = io_inValid_47 & _T_37815; // @[Switch.scala 30:36:@16896.4]
  assign _T_37818 = io_inAddr_48 == 6'h34; // @[Switch.scala 30:53:@16898.4]
  assign valid_52_48 = io_inValid_48 & _T_37818; // @[Switch.scala 30:36:@16899.4]
  assign _T_37821 = io_inAddr_49 == 6'h34; // @[Switch.scala 30:53:@16901.4]
  assign valid_52_49 = io_inValid_49 & _T_37821; // @[Switch.scala 30:36:@16902.4]
  assign _T_37824 = io_inAddr_50 == 6'h34; // @[Switch.scala 30:53:@16904.4]
  assign valid_52_50 = io_inValid_50 & _T_37824; // @[Switch.scala 30:36:@16905.4]
  assign _T_37827 = io_inAddr_51 == 6'h34; // @[Switch.scala 30:53:@16907.4]
  assign valid_52_51 = io_inValid_51 & _T_37827; // @[Switch.scala 30:36:@16908.4]
  assign _T_37830 = io_inAddr_52 == 6'h34; // @[Switch.scala 30:53:@16910.4]
  assign valid_52_52 = io_inValid_52 & _T_37830; // @[Switch.scala 30:36:@16911.4]
  assign _T_37833 = io_inAddr_53 == 6'h34; // @[Switch.scala 30:53:@16913.4]
  assign valid_52_53 = io_inValid_53 & _T_37833; // @[Switch.scala 30:36:@16914.4]
  assign _T_37836 = io_inAddr_54 == 6'h34; // @[Switch.scala 30:53:@16916.4]
  assign valid_52_54 = io_inValid_54 & _T_37836; // @[Switch.scala 30:36:@16917.4]
  assign _T_37839 = io_inAddr_55 == 6'h34; // @[Switch.scala 30:53:@16919.4]
  assign valid_52_55 = io_inValid_55 & _T_37839; // @[Switch.scala 30:36:@16920.4]
  assign _T_37842 = io_inAddr_56 == 6'h34; // @[Switch.scala 30:53:@16922.4]
  assign valid_52_56 = io_inValid_56 & _T_37842; // @[Switch.scala 30:36:@16923.4]
  assign _T_37845 = io_inAddr_57 == 6'h34; // @[Switch.scala 30:53:@16925.4]
  assign valid_52_57 = io_inValid_57 & _T_37845; // @[Switch.scala 30:36:@16926.4]
  assign _T_37848 = io_inAddr_58 == 6'h34; // @[Switch.scala 30:53:@16928.4]
  assign valid_52_58 = io_inValid_58 & _T_37848; // @[Switch.scala 30:36:@16929.4]
  assign _T_37851 = io_inAddr_59 == 6'h34; // @[Switch.scala 30:53:@16931.4]
  assign valid_52_59 = io_inValid_59 & _T_37851; // @[Switch.scala 30:36:@16932.4]
  assign _T_37854 = io_inAddr_60 == 6'h34; // @[Switch.scala 30:53:@16934.4]
  assign valid_52_60 = io_inValid_60 & _T_37854; // @[Switch.scala 30:36:@16935.4]
  assign _T_37857 = io_inAddr_61 == 6'h34; // @[Switch.scala 30:53:@16937.4]
  assign valid_52_61 = io_inValid_61 & _T_37857; // @[Switch.scala 30:36:@16938.4]
  assign _T_37860 = io_inAddr_62 == 6'h34; // @[Switch.scala 30:53:@16940.4]
  assign valid_52_62 = io_inValid_62 & _T_37860; // @[Switch.scala 30:36:@16941.4]
  assign _T_37863 = io_inAddr_63 == 6'h34; // @[Switch.scala 30:53:@16943.4]
  assign valid_52_63 = io_inValid_63 & _T_37863; // @[Switch.scala 30:36:@16944.4]
  assign _T_37929 = valid_52_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@16946.4]
  assign _T_37930 = valid_52_61 ? 6'h3d : _T_37929; // @[Mux.scala 31:69:@16947.4]
  assign _T_37931 = valid_52_60 ? 6'h3c : _T_37930; // @[Mux.scala 31:69:@16948.4]
  assign _T_37932 = valid_52_59 ? 6'h3b : _T_37931; // @[Mux.scala 31:69:@16949.4]
  assign _T_37933 = valid_52_58 ? 6'h3a : _T_37932; // @[Mux.scala 31:69:@16950.4]
  assign _T_37934 = valid_52_57 ? 6'h39 : _T_37933; // @[Mux.scala 31:69:@16951.4]
  assign _T_37935 = valid_52_56 ? 6'h38 : _T_37934; // @[Mux.scala 31:69:@16952.4]
  assign _T_37936 = valid_52_55 ? 6'h37 : _T_37935; // @[Mux.scala 31:69:@16953.4]
  assign _T_37937 = valid_52_54 ? 6'h36 : _T_37936; // @[Mux.scala 31:69:@16954.4]
  assign _T_37938 = valid_52_53 ? 6'h35 : _T_37937; // @[Mux.scala 31:69:@16955.4]
  assign _T_37939 = valid_52_52 ? 6'h34 : _T_37938; // @[Mux.scala 31:69:@16956.4]
  assign _T_37940 = valid_52_51 ? 6'h33 : _T_37939; // @[Mux.scala 31:69:@16957.4]
  assign _T_37941 = valid_52_50 ? 6'h32 : _T_37940; // @[Mux.scala 31:69:@16958.4]
  assign _T_37942 = valid_52_49 ? 6'h31 : _T_37941; // @[Mux.scala 31:69:@16959.4]
  assign _T_37943 = valid_52_48 ? 6'h30 : _T_37942; // @[Mux.scala 31:69:@16960.4]
  assign _T_37944 = valid_52_47 ? 6'h2f : _T_37943; // @[Mux.scala 31:69:@16961.4]
  assign _T_37945 = valid_52_46 ? 6'h2e : _T_37944; // @[Mux.scala 31:69:@16962.4]
  assign _T_37946 = valid_52_45 ? 6'h2d : _T_37945; // @[Mux.scala 31:69:@16963.4]
  assign _T_37947 = valid_52_44 ? 6'h2c : _T_37946; // @[Mux.scala 31:69:@16964.4]
  assign _T_37948 = valid_52_43 ? 6'h2b : _T_37947; // @[Mux.scala 31:69:@16965.4]
  assign _T_37949 = valid_52_42 ? 6'h2a : _T_37948; // @[Mux.scala 31:69:@16966.4]
  assign _T_37950 = valid_52_41 ? 6'h29 : _T_37949; // @[Mux.scala 31:69:@16967.4]
  assign _T_37951 = valid_52_40 ? 6'h28 : _T_37950; // @[Mux.scala 31:69:@16968.4]
  assign _T_37952 = valid_52_39 ? 6'h27 : _T_37951; // @[Mux.scala 31:69:@16969.4]
  assign _T_37953 = valid_52_38 ? 6'h26 : _T_37952; // @[Mux.scala 31:69:@16970.4]
  assign _T_37954 = valid_52_37 ? 6'h25 : _T_37953; // @[Mux.scala 31:69:@16971.4]
  assign _T_37955 = valid_52_36 ? 6'h24 : _T_37954; // @[Mux.scala 31:69:@16972.4]
  assign _T_37956 = valid_52_35 ? 6'h23 : _T_37955; // @[Mux.scala 31:69:@16973.4]
  assign _T_37957 = valid_52_34 ? 6'h22 : _T_37956; // @[Mux.scala 31:69:@16974.4]
  assign _T_37958 = valid_52_33 ? 6'h21 : _T_37957; // @[Mux.scala 31:69:@16975.4]
  assign _T_37959 = valid_52_32 ? 6'h20 : _T_37958; // @[Mux.scala 31:69:@16976.4]
  assign _T_37960 = valid_52_31 ? 6'h1f : _T_37959; // @[Mux.scala 31:69:@16977.4]
  assign _T_37961 = valid_52_30 ? 6'h1e : _T_37960; // @[Mux.scala 31:69:@16978.4]
  assign _T_37962 = valid_52_29 ? 6'h1d : _T_37961; // @[Mux.scala 31:69:@16979.4]
  assign _T_37963 = valid_52_28 ? 6'h1c : _T_37962; // @[Mux.scala 31:69:@16980.4]
  assign _T_37964 = valid_52_27 ? 6'h1b : _T_37963; // @[Mux.scala 31:69:@16981.4]
  assign _T_37965 = valid_52_26 ? 6'h1a : _T_37964; // @[Mux.scala 31:69:@16982.4]
  assign _T_37966 = valid_52_25 ? 6'h19 : _T_37965; // @[Mux.scala 31:69:@16983.4]
  assign _T_37967 = valid_52_24 ? 6'h18 : _T_37966; // @[Mux.scala 31:69:@16984.4]
  assign _T_37968 = valid_52_23 ? 6'h17 : _T_37967; // @[Mux.scala 31:69:@16985.4]
  assign _T_37969 = valid_52_22 ? 6'h16 : _T_37968; // @[Mux.scala 31:69:@16986.4]
  assign _T_37970 = valid_52_21 ? 6'h15 : _T_37969; // @[Mux.scala 31:69:@16987.4]
  assign _T_37971 = valid_52_20 ? 6'h14 : _T_37970; // @[Mux.scala 31:69:@16988.4]
  assign _T_37972 = valid_52_19 ? 6'h13 : _T_37971; // @[Mux.scala 31:69:@16989.4]
  assign _T_37973 = valid_52_18 ? 6'h12 : _T_37972; // @[Mux.scala 31:69:@16990.4]
  assign _T_37974 = valid_52_17 ? 6'h11 : _T_37973; // @[Mux.scala 31:69:@16991.4]
  assign _T_37975 = valid_52_16 ? 6'h10 : _T_37974; // @[Mux.scala 31:69:@16992.4]
  assign _T_37976 = valid_52_15 ? 6'hf : _T_37975; // @[Mux.scala 31:69:@16993.4]
  assign _T_37977 = valid_52_14 ? 6'he : _T_37976; // @[Mux.scala 31:69:@16994.4]
  assign _T_37978 = valid_52_13 ? 6'hd : _T_37977; // @[Mux.scala 31:69:@16995.4]
  assign _T_37979 = valid_52_12 ? 6'hc : _T_37978; // @[Mux.scala 31:69:@16996.4]
  assign _T_37980 = valid_52_11 ? 6'hb : _T_37979; // @[Mux.scala 31:69:@16997.4]
  assign _T_37981 = valid_52_10 ? 6'ha : _T_37980; // @[Mux.scala 31:69:@16998.4]
  assign _T_37982 = valid_52_9 ? 6'h9 : _T_37981; // @[Mux.scala 31:69:@16999.4]
  assign _T_37983 = valid_52_8 ? 6'h8 : _T_37982; // @[Mux.scala 31:69:@17000.4]
  assign _T_37984 = valid_52_7 ? 6'h7 : _T_37983; // @[Mux.scala 31:69:@17001.4]
  assign _T_37985 = valid_52_6 ? 6'h6 : _T_37984; // @[Mux.scala 31:69:@17002.4]
  assign _T_37986 = valid_52_5 ? 6'h5 : _T_37985; // @[Mux.scala 31:69:@17003.4]
  assign _T_37987 = valid_52_4 ? 6'h4 : _T_37986; // @[Mux.scala 31:69:@17004.4]
  assign _T_37988 = valid_52_3 ? 6'h3 : _T_37987; // @[Mux.scala 31:69:@17005.4]
  assign _T_37989 = valid_52_2 ? 6'h2 : _T_37988; // @[Mux.scala 31:69:@17006.4]
  assign _T_37990 = valid_52_1 ? 6'h1 : _T_37989; // @[Mux.scala 31:69:@17007.4]
  assign select_52 = valid_52_0 ? 6'h0 : _T_37990; // @[Mux.scala 31:69:@17008.4]
  assign _GEN_3329 = 6'h1 == select_52 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3330 = 6'h2 == select_52 ? io_inData_2 : _GEN_3329; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3331 = 6'h3 == select_52 ? io_inData_3 : _GEN_3330; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3332 = 6'h4 == select_52 ? io_inData_4 : _GEN_3331; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3333 = 6'h5 == select_52 ? io_inData_5 : _GEN_3332; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3334 = 6'h6 == select_52 ? io_inData_6 : _GEN_3333; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3335 = 6'h7 == select_52 ? io_inData_7 : _GEN_3334; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3336 = 6'h8 == select_52 ? io_inData_8 : _GEN_3335; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3337 = 6'h9 == select_52 ? io_inData_9 : _GEN_3336; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3338 = 6'ha == select_52 ? io_inData_10 : _GEN_3337; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3339 = 6'hb == select_52 ? io_inData_11 : _GEN_3338; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3340 = 6'hc == select_52 ? io_inData_12 : _GEN_3339; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3341 = 6'hd == select_52 ? io_inData_13 : _GEN_3340; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3342 = 6'he == select_52 ? io_inData_14 : _GEN_3341; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3343 = 6'hf == select_52 ? io_inData_15 : _GEN_3342; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3344 = 6'h10 == select_52 ? io_inData_16 : _GEN_3343; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3345 = 6'h11 == select_52 ? io_inData_17 : _GEN_3344; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3346 = 6'h12 == select_52 ? io_inData_18 : _GEN_3345; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3347 = 6'h13 == select_52 ? io_inData_19 : _GEN_3346; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3348 = 6'h14 == select_52 ? io_inData_20 : _GEN_3347; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3349 = 6'h15 == select_52 ? io_inData_21 : _GEN_3348; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3350 = 6'h16 == select_52 ? io_inData_22 : _GEN_3349; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3351 = 6'h17 == select_52 ? io_inData_23 : _GEN_3350; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3352 = 6'h18 == select_52 ? io_inData_24 : _GEN_3351; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3353 = 6'h19 == select_52 ? io_inData_25 : _GEN_3352; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3354 = 6'h1a == select_52 ? io_inData_26 : _GEN_3353; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3355 = 6'h1b == select_52 ? io_inData_27 : _GEN_3354; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3356 = 6'h1c == select_52 ? io_inData_28 : _GEN_3355; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3357 = 6'h1d == select_52 ? io_inData_29 : _GEN_3356; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3358 = 6'h1e == select_52 ? io_inData_30 : _GEN_3357; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3359 = 6'h1f == select_52 ? io_inData_31 : _GEN_3358; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3360 = 6'h20 == select_52 ? io_inData_32 : _GEN_3359; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3361 = 6'h21 == select_52 ? io_inData_33 : _GEN_3360; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3362 = 6'h22 == select_52 ? io_inData_34 : _GEN_3361; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3363 = 6'h23 == select_52 ? io_inData_35 : _GEN_3362; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3364 = 6'h24 == select_52 ? io_inData_36 : _GEN_3363; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3365 = 6'h25 == select_52 ? io_inData_37 : _GEN_3364; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3366 = 6'h26 == select_52 ? io_inData_38 : _GEN_3365; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3367 = 6'h27 == select_52 ? io_inData_39 : _GEN_3366; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3368 = 6'h28 == select_52 ? io_inData_40 : _GEN_3367; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3369 = 6'h29 == select_52 ? io_inData_41 : _GEN_3368; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3370 = 6'h2a == select_52 ? io_inData_42 : _GEN_3369; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3371 = 6'h2b == select_52 ? io_inData_43 : _GEN_3370; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3372 = 6'h2c == select_52 ? io_inData_44 : _GEN_3371; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3373 = 6'h2d == select_52 ? io_inData_45 : _GEN_3372; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3374 = 6'h2e == select_52 ? io_inData_46 : _GEN_3373; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3375 = 6'h2f == select_52 ? io_inData_47 : _GEN_3374; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3376 = 6'h30 == select_52 ? io_inData_48 : _GEN_3375; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3377 = 6'h31 == select_52 ? io_inData_49 : _GEN_3376; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3378 = 6'h32 == select_52 ? io_inData_50 : _GEN_3377; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3379 = 6'h33 == select_52 ? io_inData_51 : _GEN_3378; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3380 = 6'h34 == select_52 ? io_inData_52 : _GEN_3379; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3381 = 6'h35 == select_52 ? io_inData_53 : _GEN_3380; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3382 = 6'h36 == select_52 ? io_inData_54 : _GEN_3381; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3383 = 6'h37 == select_52 ? io_inData_55 : _GEN_3382; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3384 = 6'h38 == select_52 ? io_inData_56 : _GEN_3383; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3385 = 6'h39 == select_52 ? io_inData_57 : _GEN_3384; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3386 = 6'h3a == select_52 ? io_inData_58 : _GEN_3385; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3387 = 6'h3b == select_52 ? io_inData_59 : _GEN_3386; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3388 = 6'h3c == select_52 ? io_inData_60 : _GEN_3387; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3389 = 6'h3d == select_52 ? io_inData_61 : _GEN_3388; // @[Switch.scala 33:19:@17010.4]
  assign _GEN_3390 = 6'h3e == select_52 ? io_inData_62 : _GEN_3389; // @[Switch.scala 33:19:@17010.4]
  assign _T_37999 = {valid_52_7,valid_52_6,valid_52_5,valid_52_4,valid_52_3,valid_52_2,valid_52_1,valid_52_0}; // @[Switch.scala 34:32:@17017.4]
  assign _T_38007 = {valid_52_15,valid_52_14,valid_52_13,valid_52_12,valid_52_11,valid_52_10,valid_52_9,valid_52_8,_T_37999}; // @[Switch.scala 34:32:@17025.4]
  assign _T_38014 = {valid_52_23,valid_52_22,valid_52_21,valid_52_20,valid_52_19,valid_52_18,valid_52_17,valid_52_16}; // @[Switch.scala 34:32:@17032.4]
  assign _T_38023 = {valid_52_31,valid_52_30,valid_52_29,valid_52_28,valid_52_27,valid_52_26,valid_52_25,valid_52_24,_T_38014,_T_38007}; // @[Switch.scala 34:32:@17041.4]
  assign _T_38030 = {valid_52_39,valid_52_38,valid_52_37,valid_52_36,valid_52_35,valid_52_34,valid_52_33,valid_52_32}; // @[Switch.scala 34:32:@17048.4]
  assign _T_38038 = {valid_52_47,valid_52_46,valid_52_45,valid_52_44,valid_52_43,valid_52_42,valid_52_41,valid_52_40,_T_38030}; // @[Switch.scala 34:32:@17056.4]
  assign _T_38045 = {valid_52_55,valid_52_54,valid_52_53,valid_52_52,valid_52_51,valid_52_50,valid_52_49,valid_52_48}; // @[Switch.scala 34:32:@17063.4]
  assign _T_38054 = {valid_52_63,valid_52_62,valid_52_61,valid_52_60,valid_52_59,valid_52_58,valid_52_57,valid_52_56,_T_38045,_T_38038}; // @[Switch.scala 34:32:@17072.4]
  assign _T_38055 = {_T_38054,_T_38023}; // @[Switch.scala 34:32:@17073.4]
  assign _T_38059 = io_inAddr_0 == 6'h35; // @[Switch.scala 30:53:@17076.4]
  assign valid_53_0 = io_inValid_0 & _T_38059; // @[Switch.scala 30:36:@17077.4]
  assign _T_38062 = io_inAddr_1 == 6'h35; // @[Switch.scala 30:53:@17079.4]
  assign valid_53_1 = io_inValid_1 & _T_38062; // @[Switch.scala 30:36:@17080.4]
  assign _T_38065 = io_inAddr_2 == 6'h35; // @[Switch.scala 30:53:@17082.4]
  assign valid_53_2 = io_inValid_2 & _T_38065; // @[Switch.scala 30:36:@17083.4]
  assign _T_38068 = io_inAddr_3 == 6'h35; // @[Switch.scala 30:53:@17085.4]
  assign valid_53_3 = io_inValid_3 & _T_38068; // @[Switch.scala 30:36:@17086.4]
  assign _T_38071 = io_inAddr_4 == 6'h35; // @[Switch.scala 30:53:@17088.4]
  assign valid_53_4 = io_inValid_4 & _T_38071; // @[Switch.scala 30:36:@17089.4]
  assign _T_38074 = io_inAddr_5 == 6'h35; // @[Switch.scala 30:53:@17091.4]
  assign valid_53_5 = io_inValid_5 & _T_38074; // @[Switch.scala 30:36:@17092.4]
  assign _T_38077 = io_inAddr_6 == 6'h35; // @[Switch.scala 30:53:@17094.4]
  assign valid_53_6 = io_inValid_6 & _T_38077; // @[Switch.scala 30:36:@17095.4]
  assign _T_38080 = io_inAddr_7 == 6'h35; // @[Switch.scala 30:53:@17097.4]
  assign valid_53_7 = io_inValid_7 & _T_38080; // @[Switch.scala 30:36:@17098.4]
  assign _T_38083 = io_inAddr_8 == 6'h35; // @[Switch.scala 30:53:@17100.4]
  assign valid_53_8 = io_inValid_8 & _T_38083; // @[Switch.scala 30:36:@17101.4]
  assign _T_38086 = io_inAddr_9 == 6'h35; // @[Switch.scala 30:53:@17103.4]
  assign valid_53_9 = io_inValid_9 & _T_38086; // @[Switch.scala 30:36:@17104.4]
  assign _T_38089 = io_inAddr_10 == 6'h35; // @[Switch.scala 30:53:@17106.4]
  assign valid_53_10 = io_inValid_10 & _T_38089; // @[Switch.scala 30:36:@17107.4]
  assign _T_38092 = io_inAddr_11 == 6'h35; // @[Switch.scala 30:53:@17109.4]
  assign valid_53_11 = io_inValid_11 & _T_38092; // @[Switch.scala 30:36:@17110.4]
  assign _T_38095 = io_inAddr_12 == 6'h35; // @[Switch.scala 30:53:@17112.4]
  assign valid_53_12 = io_inValid_12 & _T_38095; // @[Switch.scala 30:36:@17113.4]
  assign _T_38098 = io_inAddr_13 == 6'h35; // @[Switch.scala 30:53:@17115.4]
  assign valid_53_13 = io_inValid_13 & _T_38098; // @[Switch.scala 30:36:@17116.4]
  assign _T_38101 = io_inAddr_14 == 6'h35; // @[Switch.scala 30:53:@17118.4]
  assign valid_53_14 = io_inValid_14 & _T_38101; // @[Switch.scala 30:36:@17119.4]
  assign _T_38104 = io_inAddr_15 == 6'h35; // @[Switch.scala 30:53:@17121.4]
  assign valid_53_15 = io_inValid_15 & _T_38104; // @[Switch.scala 30:36:@17122.4]
  assign _T_38107 = io_inAddr_16 == 6'h35; // @[Switch.scala 30:53:@17124.4]
  assign valid_53_16 = io_inValid_16 & _T_38107; // @[Switch.scala 30:36:@17125.4]
  assign _T_38110 = io_inAddr_17 == 6'h35; // @[Switch.scala 30:53:@17127.4]
  assign valid_53_17 = io_inValid_17 & _T_38110; // @[Switch.scala 30:36:@17128.4]
  assign _T_38113 = io_inAddr_18 == 6'h35; // @[Switch.scala 30:53:@17130.4]
  assign valid_53_18 = io_inValid_18 & _T_38113; // @[Switch.scala 30:36:@17131.4]
  assign _T_38116 = io_inAddr_19 == 6'h35; // @[Switch.scala 30:53:@17133.4]
  assign valid_53_19 = io_inValid_19 & _T_38116; // @[Switch.scala 30:36:@17134.4]
  assign _T_38119 = io_inAddr_20 == 6'h35; // @[Switch.scala 30:53:@17136.4]
  assign valid_53_20 = io_inValid_20 & _T_38119; // @[Switch.scala 30:36:@17137.4]
  assign _T_38122 = io_inAddr_21 == 6'h35; // @[Switch.scala 30:53:@17139.4]
  assign valid_53_21 = io_inValid_21 & _T_38122; // @[Switch.scala 30:36:@17140.4]
  assign _T_38125 = io_inAddr_22 == 6'h35; // @[Switch.scala 30:53:@17142.4]
  assign valid_53_22 = io_inValid_22 & _T_38125; // @[Switch.scala 30:36:@17143.4]
  assign _T_38128 = io_inAddr_23 == 6'h35; // @[Switch.scala 30:53:@17145.4]
  assign valid_53_23 = io_inValid_23 & _T_38128; // @[Switch.scala 30:36:@17146.4]
  assign _T_38131 = io_inAddr_24 == 6'h35; // @[Switch.scala 30:53:@17148.4]
  assign valid_53_24 = io_inValid_24 & _T_38131; // @[Switch.scala 30:36:@17149.4]
  assign _T_38134 = io_inAddr_25 == 6'h35; // @[Switch.scala 30:53:@17151.4]
  assign valid_53_25 = io_inValid_25 & _T_38134; // @[Switch.scala 30:36:@17152.4]
  assign _T_38137 = io_inAddr_26 == 6'h35; // @[Switch.scala 30:53:@17154.4]
  assign valid_53_26 = io_inValid_26 & _T_38137; // @[Switch.scala 30:36:@17155.4]
  assign _T_38140 = io_inAddr_27 == 6'h35; // @[Switch.scala 30:53:@17157.4]
  assign valid_53_27 = io_inValid_27 & _T_38140; // @[Switch.scala 30:36:@17158.4]
  assign _T_38143 = io_inAddr_28 == 6'h35; // @[Switch.scala 30:53:@17160.4]
  assign valid_53_28 = io_inValid_28 & _T_38143; // @[Switch.scala 30:36:@17161.4]
  assign _T_38146 = io_inAddr_29 == 6'h35; // @[Switch.scala 30:53:@17163.4]
  assign valid_53_29 = io_inValid_29 & _T_38146; // @[Switch.scala 30:36:@17164.4]
  assign _T_38149 = io_inAddr_30 == 6'h35; // @[Switch.scala 30:53:@17166.4]
  assign valid_53_30 = io_inValid_30 & _T_38149; // @[Switch.scala 30:36:@17167.4]
  assign _T_38152 = io_inAddr_31 == 6'h35; // @[Switch.scala 30:53:@17169.4]
  assign valid_53_31 = io_inValid_31 & _T_38152; // @[Switch.scala 30:36:@17170.4]
  assign _T_38155 = io_inAddr_32 == 6'h35; // @[Switch.scala 30:53:@17172.4]
  assign valid_53_32 = io_inValid_32 & _T_38155; // @[Switch.scala 30:36:@17173.4]
  assign _T_38158 = io_inAddr_33 == 6'h35; // @[Switch.scala 30:53:@17175.4]
  assign valid_53_33 = io_inValid_33 & _T_38158; // @[Switch.scala 30:36:@17176.4]
  assign _T_38161 = io_inAddr_34 == 6'h35; // @[Switch.scala 30:53:@17178.4]
  assign valid_53_34 = io_inValid_34 & _T_38161; // @[Switch.scala 30:36:@17179.4]
  assign _T_38164 = io_inAddr_35 == 6'h35; // @[Switch.scala 30:53:@17181.4]
  assign valid_53_35 = io_inValid_35 & _T_38164; // @[Switch.scala 30:36:@17182.4]
  assign _T_38167 = io_inAddr_36 == 6'h35; // @[Switch.scala 30:53:@17184.4]
  assign valid_53_36 = io_inValid_36 & _T_38167; // @[Switch.scala 30:36:@17185.4]
  assign _T_38170 = io_inAddr_37 == 6'h35; // @[Switch.scala 30:53:@17187.4]
  assign valid_53_37 = io_inValid_37 & _T_38170; // @[Switch.scala 30:36:@17188.4]
  assign _T_38173 = io_inAddr_38 == 6'h35; // @[Switch.scala 30:53:@17190.4]
  assign valid_53_38 = io_inValid_38 & _T_38173; // @[Switch.scala 30:36:@17191.4]
  assign _T_38176 = io_inAddr_39 == 6'h35; // @[Switch.scala 30:53:@17193.4]
  assign valid_53_39 = io_inValid_39 & _T_38176; // @[Switch.scala 30:36:@17194.4]
  assign _T_38179 = io_inAddr_40 == 6'h35; // @[Switch.scala 30:53:@17196.4]
  assign valid_53_40 = io_inValid_40 & _T_38179; // @[Switch.scala 30:36:@17197.4]
  assign _T_38182 = io_inAddr_41 == 6'h35; // @[Switch.scala 30:53:@17199.4]
  assign valid_53_41 = io_inValid_41 & _T_38182; // @[Switch.scala 30:36:@17200.4]
  assign _T_38185 = io_inAddr_42 == 6'h35; // @[Switch.scala 30:53:@17202.4]
  assign valid_53_42 = io_inValid_42 & _T_38185; // @[Switch.scala 30:36:@17203.4]
  assign _T_38188 = io_inAddr_43 == 6'h35; // @[Switch.scala 30:53:@17205.4]
  assign valid_53_43 = io_inValid_43 & _T_38188; // @[Switch.scala 30:36:@17206.4]
  assign _T_38191 = io_inAddr_44 == 6'h35; // @[Switch.scala 30:53:@17208.4]
  assign valid_53_44 = io_inValid_44 & _T_38191; // @[Switch.scala 30:36:@17209.4]
  assign _T_38194 = io_inAddr_45 == 6'h35; // @[Switch.scala 30:53:@17211.4]
  assign valid_53_45 = io_inValid_45 & _T_38194; // @[Switch.scala 30:36:@17212.4]
  assign _T_38197 = io_inAddr_46 == 6'h35; // @[Switch.scala 30:53:@17214.4]
  assign valid_53_46 = io_inValid_46 & _T_38197; // @[Switch.scala 30:36:@17215.4]
  assign _T_38200 = io_inAddr_47 == 6'h35; // @[Switch.scala 30:53:@17217.4]
  assign valid_53_47 = io_inValid_47 & _T_38200; // @[Switch.scala 30:36:@17218.4]
  assign _T_38203 = io_inAddr_48 == 6'h35; // @[Switch.scala 30:53:@17220.4]
  assign valid_53_48 = io_inValid_48 & _T_38203; // @[Switch.scala 30:36:@17221.4]
  assign _T_38206 = io_inAddr_49 == 6'h35; // @[Switch.scala 30:53:@17223.4]
  assign valid_53_49 = io_inValid_49 & _T_38206; // @[Switch.scala 30:36:@17224.4]
  assign _T_38209 = io_inAddr_50 == 6'h35; // @[Switch.scala 30:53:@17226.4]
  assign valid_53_50 = io_inValid_50 & _T_38209; // @[Switch.scala 30:36:@17227.4]
  assign _T_38212 = io_inAddr_51 == 6'h35; // @[Switch.scala 30:53:@17229.4]
  assign valid_53_51 = io_inValid_51 & _T_38212; // @[Switch.scala 30:36:@17230.4]
  assign _T_38215 = io_inAddr_52 == 6'h35; // @[Switch.scala 30:53:@17232.4]
  assign valid_53_52 = io_inValid_52 & _T_38215; // @[Switch.scala 30:36:@17233.4]
  assign _T_38218 = io_inAddr_53 == 6'h35; // @[Switch.scala 30:53:@17235.4]
  assign valid_53_53 = io_inValid_53 & _T_38218; // @[Switch.scala 30:36:@17236.4]
  assign _T_38221 = io_inAddr_54 == 6'h35; // @[Switch.scala 30:53:@17238.4]
  assign valid_53_54 = io_inValid_54 & _T_38221; // @[Switch.scala 30:36:@17239.4]
  assign _T_38224 = io_inAddr_55 == 6'h35; // @[Switch.scala 30:53:@17241.4]
  assign valid_53_55 = io_inValid_55 & _T_38224; // @[Switch.scala 30:36:@17242.4]
  assign _T_38227 = io_inAddr_56 == 6'h35; // @[Switch.scala 30:53:@17244.4]
  assign valid_53_56 = io_inValid_56 & _T_38227; // @[Switch.scala 30:36:@17245.4]
  assign _T_38230 = io_inAddr_57 == 6'h35; // @[Switch.scala 30:53:@17247.4]
  assign valid_53_57 = io_inValid_57 & _T_38230; // @[Switch.scala 30:36:@17248.4]
  assign _T_38233 = io_inAddr_58 == 6'h35; // @[Switch.scala 30:53:@17250.4]
  assign valid_53_58 = io_inValid_58 & _T_38233; // @[Switch.scala 30:36:@17251.4]
  assign _T_38236 = io_inAddr_59 == 6'h35; // @[Switch.scala 30:53:@17253.4]
  assign valid_53_59 = io_inValid_59 & _T_38236; // @[Switch.scala 30:36:@17254.4]
  assign _T_38239 = io_inAddr_60 == 6'h35; // @[Switch.scala 30:53:@17256.4]
  assign valid_53_60 = io_inValid_60 & _T_38239; // @[Switch.scala 30:36:@17257.4]
  assign _T_38242 = io_inAddr_61 == 6'h35; // @[Switch.scala 30:53:@17259.4]
  assign valid_53_61 = io_inValid_61 & _T_38242; // @[Switch.scala 30:36:@17260.4]
  assign _T_38245 = io_inAddr_62 == 6'h35; // @[Switch.scala 30:53:@17262.4]
  assign valid_53_62 = io_inValid_62 & _T_38245; // @[Switch.scala 30:36:@17263.4]
  assign _T_38248 = io_inAddr_63 == 6'h35; // @[Switch.scala 30:53:@17265.4]
  assign valid_53_63 = io_inValid_63 & _T_38248; // @[Switch.scala 30:36:@17266.4]
  assign _T_38314 = valid_53_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@17268.4]
  assign _T_38315 = valid_53_61 ? 6'h3d : _T_38314; // @[Mux.scala 31:69:@17269.4]
  assign _T_38316 = valid_53_60 ? 6'h3c : _T_38315; // @[Mux.scala 31:69:@17270.4]
  assign _T_38317 = valid_53_59 ? 6'h3b : _T_38316; // @[Mux.scala 31:69:@17271.4]
  assign _T_38318 = valid_53_58 ? 6'h3a : _T_38317; // @[Mux.scala 31:69:@17272.4]
  assign _T_38319 = valid_53_57 ? 6'h39 : _T_38318; // @[Mux.scala 31:69:@17273.4]
  assign _T_38320 = valid_53_56 ? 6'h38 : _T_38319; // @[Mux.scala 31:69:@17274.4]
  assign _T_38321 = valid_53_55 ? 6'h37 : _T_38320; // @[Mux.scala 31:69:@17275.4]
  assign _T_38322 = valid_53_54 ? 6'h36 : _T_38321; // @[Mux.scala 31:69:@17276.4]
  assign _T_38323 = valid_53_53 ? 6'h35 : _T_38322; // @[Mux.scala 31:69:@17277.4]
  assign _T_38324 = valid_53_52 ? 6'h34 : _T_38323; // @[Mux.scala 31:69:@17278.4]
  assign _T_38325 = valid_53_51 ? 6'h33 : _T_38324; // @[Mux.scala 31:69:@17279.4]
  assign _T_38326 = valid_53_50 ? 6'h32 : _T_38325; // @[Mux.scala 31:69:@17280.4]
  assign _T_38327 = valid_53_49 ? 6'h31 : _T_38326; // @[Mux.scala 31:69:@17281.4]
  assign _T_38328 = valid_53_48 ? 6'h30 : _T_38327; // @[Mux.scala 31:69:@17282.4]
  assign _T_38329 = valid_53_47 ? 6'h2f : _T_38328; // @[Mux.scala 31:69:@17283.4]
  assign _T_38330 = valid_53_46 ? 6'h2e : _T_38329; // @[Mux.scala 31:69:@17284.4]
  assign _T_38331 = valid_53_45 ? 6'h2d : _T_38330; // @[Mux.scala 31:69:@17285.4]
  assign _T_38332 = valid_53_44 ? 6'h2c : _T_38331; // @[Mux.scala 31:69:@17286.4]
  assign _T_38333 = valid_53_43 ? 6'h2b : _T_38332; // @[Mux.scala 31:69:@17287.4]
  assign _T_38334 = valid_53_42 ? 6'h2a : _T_38333; // @[Mux.scala 31:69:@17288.4]
  assign _T_38335 = valid_53_41 ? 6'h29 : _T_38334; // @[Mux.scala 31:69:@17289.4]
  assign _T_38336 = valid_53_40 ? 6'h28 : _T_38335; // @[Mux.scala 31:69:@17290.4]
  assign _T_38337 = valid_53_39 ? 6'h27 : _T_38336; // @[Mux.scala 31:69:@17291.4]
  assign _T_38338 = valid_53_38 ? 6'h26 : _T_38337; // @[Mux.scala 31:69:@17292.4]
  assign _T_38339 = valid_53_37 ? 6'h25 : _T_38338; // @[Mux.scala 31:69:@17293.4]
  assign _T_38340 = valid_53_36 ? 6'h24 : _T_38339; // @[Mux.scala 31:69:@17294.4]
  assign _T_38341 = valid_53_35 ? 6'h23 : _T_38340; // @[Mux.scala 31:69:@17295.4]
  assign _T_38342 = valid_53_34 ? 6'h22 : _T_38341; // @[Mux.scala 31:69:@17296.4]
  assign _T_38343 = valid_53_33 ? 6'h21 : _T_38342; // @[Mux.scala 31:69:@17297.4]
  assign _T_38344 = valid_53_32 ? 6'h20 : _T_38343; // @[Mux.scala 31:69:@17298.4]
  assign _T_38345 = valid_53_31 ? 6'h1f : _T_38344; // @[Mux.scala 31:69:@17299.4]
  assign _T_38346 = valid_53_30 ? 6'h1e : _T_38345; // @[Mux.scala 31:69:@17300.4]
  assign _T_38347 = valid_53_29 ? 6'h1d : _T_38346; // @[Mux.scala 31:69:@17301.4]
  assign _T_38348 = valid_53_28 ? 6'h1c : _T_38347; // @[Mux.scala 31:69:@17302.4]
  assign _T_38349 = valid_53_27 ? 6'h1b : _T_38348; // @[Mux.scala 31:69:@17303.4]
  assign _T_38350 = valid_53_26 ? 6'h1a : _T_38349; // @[Mux.scala 31:69:@17304.4]
  assign _T_38351 = valid_53_25 ? 6'h19 : _T_38350; // @[Mux.scala 31:69:@17305.4]
  assign _T_38352 = valid_53_24 ? 6'h18 : _T_38351; // @[Mux.scala 31:69:@17306.4]
  assign _T_38353 = valid_53_23 ? 6'h17 : _T_38352; // @[Mux.scala 31:69:@17307.4]
  assign _T_38354 = valid_53_22 ? 6'h16 : _T_38353; // @[Mux.scala 31:69:@17308.4]
  assign _T_38355 = valid_53_21 ? 6'h15 : _T_38354; // @[Mux.scala 31:69:@17309.4]
  assign _T_38356 = valid_53_20 ? 6'h14 : _T_38355; // @[Mux.scala 31:69:@17310.4]
  assign _T_38357 = valid_53_19 ? 6'h13 : _T_38356; // @[Mux.scala 31:69:@17311.4]
  assign _T_38358 = valid_53_18 ? 6'h12 : _T_38357; // @[Mux.scala 31:69:@17312.4]
  assign _T_38359 = valid_53_17 ? 6'h11 : _T_38358; // @[Mux.scala 31:69:@17313.4]
  assign _T_38360 = valid_53_16 ? 6'h10 : _T_38359; // @[Mux.scala 31:69:@17314.4]
  assign _T_38361 = valid_53_15 ? 6'hf : _T_38360; // @[Mux.scala 31:69:@17315.4]
  assign _T_38362 = valid_53_14 ? 6'he : _T_38361; // @[Mux.scala 31:69:@17316.4]
  assign _T_38363 = valid_53_13 ? 6'hd : _T_38362; // @[Mux.scala 31:69:@17317.4]
  assign _T_38364 = valid_53_12 ? 6'hc : _T_38363; // @[Mux.scala 31:69:@17318.4]
  assign _T_38365 = valid_53_11 ? 6'hb : _T_38364; // @[Mux.scala 31:69:@17319.4]
  assign _T_38366 = valid_53_10 ? 6'ha : _T_38365; // @[Mux.scala 31:69:@17320.4]
  assign _T_38367 = valid_53_9 ? 6'h9 : _T_38366; // @[Mux.scala 31:69:@17321.4]
  assign _T_38368 = valid_53_8 ? 6'h8 : _T_38367; // @[Mux.scala 31:69:@17322.4]
  assign _T_38369 = valid_53_7 ? 6'h7 : _T_38368; // @[Mux.scala 31:69:@17323.4]
  assign _T_38370 = valid_53_6 ? 6'h6 : _T_38369; // @[Mux.scala 31:69:@17324.4]
  assign _T_38371 = valid_53_5 ? 6'h5 : _T_38370; // @[Mux.scala 31:69:@17325.4]
  assign _T_38372 = valid_53_4 ? 6'h4 : _T_38371; // @[Mux.scala 31:69:@17326.4]
  assign _T_38373 = valid_53_3 ? 6'h3 : _T_38372; // @[Mux.scala 31:69:@17327.4]
  assign _T_38374 = valid_53_2 ? 6'h2 : _T_38373; // @[Mux.scala 31:69:@17328.4]
  assign _T_38375 = valid_53_1 ? 6'h1 : _T_38374; // @[Mux.scala 31:69:@17329.4]
  assign select_53 = valid_53_0 ? 6'h0 : _T_38375; // @[Mux.scala 31:69:@17330.4]
  assign _GEN_3393 = 6'h1 == select_53 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3394 = 6'h2 == select_53 ? io_inData_2 : _GEN_3393; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3395 = 6'h3 == select_53 ? io_inData_3 : _GEN_3394; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3396 = 6'h4 == select_53 ? io_inData_4 : _GEN_3395; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3397 = 6'h5 == select_53 ? io_inData_5 : _GEN_3396; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3398 = 6'h6 == select_53 ? io_inData_6 : _GEN_3397; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3399 = 6'h7 == select_53 ? io_inData_7 : _GEN_3398; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3400 = 6'h8 == select_53 ? io_inData_8 : _GEN_3399; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3401 = 6'h9 == select_53 ? io_inData_9 : _GEN_3400; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3402 = 6'ha == select_53 ? io_inData_10 : _GEN_3401; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3403 = 6'hb == select_53 ? io_inData_11 : _GEN_3402; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3404 = 6'hc == select_53 ? io_inData_12 : _GEN_3403; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3405 = 6'hd == select_53 ? io_inData_13 : _GEN_3404; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3406 = 6'he == select_53 ? io_inData_14 : _GEN_3405; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3407 = 6'hf == select_53 ? io_inData_15 : _GEN_3406; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3408 = 6'h10 == select_53 ? io_inData_16 : _GEN_3407; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3409 = 6'h11 == select_53 ? io_inData_17 : _GEN_3408; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3410 = 6'h12 == select_53 ? io_inData_18 : _GEN_3409; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3411 = 6'h13 == select_53 ? io_inData_19 : _GEN_3410; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3412 = 6'h14 == select_53 ? io_inData_20 : _GEN_3411; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3413 = 6'h15 == select_53 ? io_inData_21 : _GEN_3412; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3414 = 6'h16 == select_53 ? io_inData_22 : _GEN_3413; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3415 = 6'h17 == select_53 ? io_inData_23 : _GEN_3414; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3416 = 6'h18 == select_53 ? io_inData_24 : _GEN_3415; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3417 = 6'h19 == select_53 ? io_inData_25 : _GEN_3416; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3418 = 6'h1a == select_53 ? io_inData_26 : _GEN_3417; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3419 = 6'h1b == select_53 ? io_inData_27 : _GEN_3418; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3420 = 6'h1c == select_53 ? io_inData_28 : _GEN_3419; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3421 = 6'h1d == select_53 ? io_inData_29 : _GEN_3420; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3422 = 6'h1e == select_53 ? io_inData_30 : _GEN_3421; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3423 = 6'h1f == select_53 ? io_inData_31 : _GEN_3422; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3424 = 6'h20 == select_53 ? io_inData_32 : _GEN_3423; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3425 = 6'h21 == select_53 ? io_inData_33 : _GEN_3424; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3426 = 6'h22 == select_53 ? io_inData_34 : _GEN_3425; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3427 = 6'h23 == select_53 ? io_inData_35 : _GEN_3426; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3428 = 6'h24 == select_53 ? io_inData_36 : _GEN_3427; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3429 = 6'h25 == select_53 ? io_inData_37 : _GEN_3428; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3430 = 6'h26 == select_53 ? io_inData_38 : _GEN_3429; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3431 = 6'h27 == select_53 ? io_inData_39 : _GEN_3430; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3432 = 6'h28 == select_53 ? io_inData_40 : _GEN_3431; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3433 = 6'h29 == select_53 ? io_inData_41 : _GEN_3432; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3434 = 6'h2a == select_53 ? io_inData_42 : _GEN_3433; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3435 = 6'h2b == select_53 ? io_inData_43 : _GEN_3434; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3436 = 6'h2c == select_53 ? io_inData_44 : _GEN_3435; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3437 = 6'h2d == select_53 ? io_inData_45 : _GEN_3436; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3438 = 6'h2e == select_53 ? io_inData_46 : _GEN_3437; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3439 = 6'h2f == select_53 ? io_inData_47 : _GEN_3438; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3440 = 6'h30 == select_53 ? io_inData_48 : _GEN_3439; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3441 = 6'h31 == select_53 ? io_inData_49 : _GEN_3440; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3442 = 6'h32 == select_53 ? io_inData_50 : _GEN_3441; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3443 = 6'h33 == select_53 ? io_inData_51 : _GEN_3442; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3444 = 6'h34 == select_53 ? io_inData_52 : _GEN_3443; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3445 = 6'h35 == select_53 ? io_inData_53 : _GEN_3444; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3446 = 6'h36 == select_53 ? io_inData_54 : _GEN_3445; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3447 = 6'h37 == select_53 ? io_inData_55 : _GEN_3446; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3448 = 6'h38 == select_53 ? io_inData_56 : _GEN_3447; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3449 = 6'h39 == select_53 ? io_inData_57 : _GEN_3448; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3450 = 6'h3a == select_53 ? io_inData_58 : _GEN_3449; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3451 = 6'h3b == select_53 ? io_inData_59 : _GEN_3450; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3452 = 6'h3c == select_53 ? io_inData_60 : _GEN_3451; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3453 = 6'h3d == select_53 ? io_inData_61 : _GEN_3452; // @[Switch.scala 33:19:@17332.4]
  assign _GEN_3454 = 6'h3e == select_53 ? io_inData_62 : _GEN_3453; // @[Switch.scala 33:19:@17332.4]
  assign _T_38384 = {valid_53_7,valid_53_6,valid_53_5,valid_53_4,valid_53_3,valid_53_2,valid_53_1,valid_53_0}; // @[Switch.scala 34:32:@17339.4]
  assign _T_38392 = {valid_53_15,valid_53_14,valid_53_13,valid_53_12,valid_53_11,valid_53_10,valid_53_9,valid_53_8,_T_38384}; // @[Switch.scala 34:32:@17347.4]
  assign _T_38399 = {valid_53_23,valid_53_22,valid_53_21,valid_53_20,valid_53_19,valid_53_18,valid_53_17,valid_53_16}; // @[Switch.scala 34:32:@17354.4]
  assign _T_38408 = {valid_53_31,valid_53_30,valid_53_29,valid_53_28,valid_53_27,valid_53_26,valid_53_25,valid_53_24,_T_38399,_T_38392}; // @[Switch.scala 34:32:@17363.4]
  assign _T_38415 = {valid_53_39,valid_53_38,valid_53_37,valid_53_36,valid_53_35,valid_53_34,valid_53_33,valid_53_32}; // @[Switch.scala 34:32:@17370.4]
  assign _T_38423 = {valid_53_47,valid_53_46,valid_53_45,valid_53_44,valid_53_43,valid_53_42,valid_53_41,valid_53_40,_T_38415}; // @[Switch.scala 34:32:@17378.4]
  assign _T_38430 = {valid_53_55,valid_53_54,valid_53_53,valid_53_52,valid_53_51,valid_53_50,valid_53_49,valid_53_48}; // @[Switch.scala 34:32:@17385.4]
  assign _T_38439 = {valid_53_63,valid_53_62,valid_53_61,valid_53_60,valid_53_59,valid_53_58,valid_53_57,valid_53_56,_T_38430,_T_38423}; // @[Switch.scala 34:32:@17394.4]
  assign _T_38440 = {_T_38439,_T_38408}; // @[Switch.scala 34:32:@17395.4]
  assign _T_38444 = io_inAddr_0 == 6'h36; // @[Switch.scala 30:53:@17398.4]
  assign valid_54_0 = io_inValid_0 & _T_38444; // @[Switch.scala 30:36:@17399.4]
  assign _T_38447 = io_inAddr_1 == 6'h36; // @[Switch.scala 30:53:@17401.4]
  assign valid_54_1 = io_inValid_1 & _T_38447; // @[Switch.scala 30:36:@17402.4]
  assign _T_38450 = io_inAddr_2 == 6'h36; // @[Switch.scala 30:53:@17404.4]
  assign valid_54_2 = io_inValid_2 & _T_38450; // @[Switch.scala 30:36:@17405.4]
  assign _T_38453 = io_inAddr_3 == 6'h36; // @[Switch.scala 30:53:@17407.4]
  assign valid_54_3 = io_inValid_3 & _T_38453; // @[Switch.scala 30:36:@17408.4]
  assign _T_38456 = io_inAddr_4 == 6'h36; // @[Switch.scala 30:53:@17410.4]
  assign valid_54_4 = io_inValid_4 & _T_38456; // @[Switch.scala 30:36:@17411.4]
  assign _T_38459 = io_inAddr_5 == 6'h36; // @[Switch.scala 30:53:@17413.4]
  assign valid_54_5 = io_inValid_5 & _T_38459; // @[Switch.scala 30:36:@17414.4]
  assign _T_38462 = io_inAddr_6 == 6'h36; // @[Switch.scala 30:53:@17416.4]
  assign valid_54_6 = io_inValid_6 & _T_38462; // @[Switch.scala 30:36:@17417.4]
  assign _T_38465 = io_inAddr_7 == 6'h36; // @[Switch.scala 30:53:@17419.4]
  assign valid_54_7 = io_inValid_7 & _T_38465; // @[Switch.scala 30:36:@17420.4]
  assign _T_38468 = io_inAddr_8 == 6'h36; // @[Switch.scala 30:53:@17422.4]
  assign valid_54_8 = io_inValid_8 & _T_38468; // @[Switch.scala 30:36:@17423.4]
  assign _T_38471 = io_inAddr_9 == 6'h36; // @[Switch.scala 30:53:@17425.4]
  assign valid_54_9 = io_inValid_9 & _T_38471; // @[Switch.scala 30:36:@17426.4]
  assign _T_38474 = io_inAddr_10 == 6'h36; // @[Switch.scala 30:53:@17428.4]
  assign valid_54_10 = io_inValid_10 & _T_38474; // @[Switch.scala 30:36:@17429.4]
  assign _T_38477 = io_inAddr_11 == 6'h36; // @[Switch.scala 30:53:@17431.4]
  assign valid_54_11 = io_inValid_11 & _T_38477; // @[Switch.scala 30:36:@17432.4]
  assign _T_38480 = io_inAddr_12 == 6'h36; // @[Switch.scala 30:53:@17434.4]
  assign valid_54_12 = io_inValid_12 & _T_38480; // @[Switch.scala 30:36:@17435.4]
  assign _T_38483 = io_inAddr_13 == 6'h36; // @[Switch.scala 30:53:@17437.4]
  assign valid_54_13 = io_inValid_13 & _T_38483; // @[Switch.scala 30:36:@17438.4]
  assign _T_38486 = io_inAddr_14 == 6'h36; // @[Switch.scala 30:53:@17440.4]
  assign valid_54_14 = io_inValid_14 & _T_38486; // @[Switch.scala 30:36:@17441.4]
  assign _T_38489 = io_inAddr_15 == 6'h36; // @[Switch.scala 30:53:@17443.4]
  assign valid_54_15 = io_inValid_15 & _T_38489; // @[Switch.scala 30:36:@17444.4]
  assign _T_38492 = io_inAddr_16 == 6'h36; // @[Switch.scala 30:53:@17446.4]
  assign valid_54_16 = io_inValid_16 & _T_38492; // @[Switch.scala 30:36:@17447.4]
  assign _T_38495 = io_inAddr_17 == 6'h36; // @[Switch.scala 30:53:@17449.4]
  assign valid_54_17 = io_inValid_17 & _T_38495; // @[Switch.scala 30:36:@17450.4]
  assign _T_38498 = io_inAddr_18 == 6'h36; // @[Switch.scala 30:53:@17452.4]
  assign valid_54_18 = io_inValid_18 & _T_38498; // @[Switch.scala 30:36:@17453.4]
  assign _T_38501 = io_inAddr_19 == 6'h36; // @[Switch.scala 30:53:@17455.4]
  assign valid_54_19 = io_inValid_19 & _T_38501; // @[Switch.scala 30:36:@17456.4]
  assign _T_38504 = io_inAddr_20 == 6'h36; // @[Switch.scala 30:53:@17458.4]
  assign valid_54_20 = io_inValid_20 & _T_38504; // @[Switch.scala 30:36:@17459.4]
  assign _T_38507 = io_inAddr_21 == 6'h36; // @[Switch.scala 30:53:@17461.4]
  assign valid_54_21 = io_inValid_21 & _T_38507; // @[Switch.scala 30:36:@17462.4]
  assign _T_38510 = io_inAddr_22 == 6'h36; // @[Switch.scala 30:53:@17464.4]
  assign valid_54_22 = io_inValid_22 & _T_38510; // @[Switch.scala 30:36:@17465.4]
  assign _T_38513 = io_inAddr_23 == 6'h36; // @[Switch.scala 30:53:@17467.4]
  assign valid_54_23 = io_inValid_23 & _T_38513; // @[Switch.scala 30:36:@17468.4]
  assign _T_38516 = io_inAddr_24 == 6'h36; // @[Switch.scala 30:53:@17470.4]
  assign valid_54_24 = io_inValid_24 & _T_38516; // @[Switch.scala 30:36:@17471.4]
  assign _T_38519 = io_inAddr_25 == 6'h36; // @[Switch.scala 30:53:@17473.4]
  assign valid_54_25 = io_inValid_25 & _T_38519; // @[Switch.scala 30:36:@17474.4]
  assign _T_38522 = io_inAddr_26 == 6'h36; // @[Switch.scala 30:53:@17476.4]
  assign valid_54_26 = io_inValid_26 & _T_38522; // @[Switch.scala 30:36:@17477.4]
  assign _T_38525 = io_inAddr_27 == 6'h36; // @[Switch.scala 30:53:@17479.4]
  assign valid_54_27 = io_inValid_27 & _T_38525; // @[Switch.scala 30:36:@17480.4]
  assign _T_38528 = io_inAddr_28 == 6'h36; // @[Switch.scala 30:53:@17482.4]
  assign valid_54_28 = io_inValid_28 & _T_38528; // @[Switch.scala 30:36:@17483.4]
  assign _T_38531 = io_inAddr_29 == 6'h36; // @[Switch.scala 30:53:@17485.4]
  assign valid_54_29 = io_inValid_29 & _T_38531; // @[Switch.scala 30:36:@17486.4]
  assign _T_38534 = io_inAddr_30 == 6'h36; // @[Switch.scala 30:53:@17488.4]
  assign valid_54_30 = io_inValid_30 & _T_38534; // @[Switch.scala 30:36:@17489.4]
  assign _T_38537 = io_inAddr_31 == 6'h36; // @[Switch.scala 30:53:@17491.4]
  assign valid_54_31 = io_inValid_31 & _T_38537; // @[Switch.scala 30:36:@17492.4]
  assign _T_38540 = io_inAddr_32 == 6'h36; // @[Switch.scala 30:53:@17494.4]
  assign valid_54_32 = io_inValid_32 & _T_38540; // @[Switch.scala 30:36:@17495.4]
  assign _T_38543 = io_inAddr_33 == 6'h36; // @[Switch.scala 30:53:@17497.4]
  assign valid_54_33 = io_inValid_33 & _T_38543; // @[Switch.scala 30:36:@17498.4]
  assign _T_38546 = io_inAddr_34 == 6'h36; // @[Switch.scala 30:53:@17500.4]
  assign valid_54_34 = io_inValid_34 & _T_38546; // @[Switch.scala 30:36:@17501.4]
  assign _T_38549 = io_inAddr_35 == 6'h36; // @[Switch.scala 30:53:@17503.4]
  assign valid_54_35 = io_inValid_35 & _T_38549; // @[Switch.scala 30:36:@17504.4]
  assign _T_38552 = io_inAddr_36 == 6'h36; // @[Switch.scala 30:53:@17506.4]
  assign valid_54_36 = io_inValid_36 & _T_38552; // @[Switch.scala 30:36:@17507.4]
  assign _T_38555 = io_inAddr_37 == 6'h36; // @[Switch.scala 30:53:@17509.4]
  assign valid_54_37 = io_inValid_37 & _T_38555; // @[Switch.scala 30:36:@17510.4]
  assign _T_38558 = io_inAddr_38 == 6'h36; // @[Switch.scala 30:53:@17512.4]
  assign valid_54_38 = io_inValid_38 & _T_38558; // @[Switch.scala 30:36:@17513.4]
  assign _T_38561 = io_inAddr_39 == 6'h36; // @[Switch.scala 30:53:@17515.4]
  assign valid_54_39 = io_inValid_39 & _T_38561; // @[Switch.scala 30:36:@17516.4]
  assign _T_38564 = io_inAddr_40 == 6'h36; // @[Switch.scala 30:53:@17518.4]
  assign valid_54_40 = io_inValid_40 & _T_38564; // @[Switch.scala 30:36:@17519.4]
  assign _T_38567 = io_inAddr_41 == 6'h36; // @[Switch.scala 30:53:@17521.4]
  assign valid_54_41 = io_inValid_41 & _T_38567; // @[Switch.scala 30:36:@17522.4]
  assign _T_38570 = io_inAddr_42 == 6'h36; // @[Switch.scala 30:53:@17524.4]
  assign valid_54_42 = io_inValid_42 & _T_38570; // @[Switch.scala 30:36:@17525.4]
  assign _T_38573 = io_inAddr_43 == 6'h36; // @[Switch.scala 30:53:@17527.4]
  assign valid_54_43 = io_inValid_43 & _T_38573; // @[Switch.scala 30:36:@17528.4]
  assign _T_38576 = io_inAddr_44 == 6'h36; // @[Switch.scala 30:53:@17530.4]
  assign valid_54_44 = io_inValid_44 & _T_38576; // @[Switch.scala 30:36:@17531.4]
  assign _T_38579 = io_inAddr_45 == 6'h36; // @[Switch.scala 30:53:@17533.4]
  assign valid_54_45 = io_inValid_45 & _T_38579; // @[Switch.scala 30:36:@17534.4]
  assign _T_38582 = io_inAddr_46 == 6'h36; // @[Switch.scala 30:53:@17536.4]
  assign valid_54_46 = io_inValid_46 & _T_38582; // @[Switch.scala 30:36:@17537.4]
  assign _T_38585 = io_inAddr_47 == 6'h36; // @[Switch.scala 30:53:@17539.4]
  assign valid_54_47 = io_inValid_47 & _T_38585; // @[Switch.scala 30:36:@17540.4]
  assign _T_38588 = io_inAddr_48 == 6'h36; // @[Switch.scala 30:53:@17542.4]
  assign valid_54_48 = io_inValid_48 & _T_38588; // @[Switch.scala 30:36:@17543.4]
  assign _T_38591 = io_inAddr_49 == 6'h36; // @[Switch.scala 30:53:@17545.4]
  assign valid_54_49 = io_inValid_49 & _T_38591; // @[Switch.scala 30:36:@17546.4]
  assign _T_38594 = io_inAddr_50 == 6'h36; // @[Switch.scala 30:53:@17548.4]
  assign valid_54_50 = io_inValid_50 & _T_38594; // @[Switch.scala 30:36:@17549.4]
  assign _T_38597 = io_inAddr_51 == 6'h36; // @[Switch.scala 30:53:@17551.4]
  assign valid_54_51 = io_inValid_51 & _T_38597; // @[Switch.scala 30:36:@17552.4]
  assign _T_38600 = io_inAddr_52 == 6'h36; // @[Switch.scala 30:53:@17554.4]
  assign valid_54_52 = io_inValid_52 & _T_38600; // @[Switch.scala 30:36:@17555.4]
  assign _T_38603 = io_inAddr_53 == 6'h36; // @[Switch.scala 30:53:@17557.4]
  assign valid_54_53 = io_inValid_53 & _T_38603; // @[Switch.scala 30:36:@17558.4]
  assign _T_38606 = io_inAddr_54 == 6'h36; // @[Switch.scala 30:53:@17560.4]
  assign valid_54_54 = io_inValid_54 & _T_38606; // @[Switch.scala 30:36:@17561.4]
  assign _T_38609 = io_inAddr_55 == 6'h36; // @[Switch.scala 30:53:@17563.4]
  assign valid_54_55 = io_inValid_55 & _T_38609; // @[Switch.scala 30:36:@17564.4]
  assign _T_38612 = io_inAddr_56 == 6'h36; // @[Switch.scala 30:53:@17566.4]
  assign valid_54_56 = io_inValid_56 & _T_38612; // @[Switch.scala 30:36:@17567.4]
  assign _T_38615 = io_inAddr_57 == 6'h36; // @[Switch.scala 30:53:@17569.4]
  assign valid_54_57 = io_inValid_57 & _T_38615; // @[Switch.scala 30:36:@17570.4]
  assign _T_38618 = io_inAddr_58 == 6'h36; // @[Switch.scala 30:53:@17572.4]
  assign valid_54_58 = io_inValid_58 & _T_38618; // @[Switch.scala 30:36:@17573.4]
  assign _T_38621 = io_inAddr_59 == 6'h36; // @[Switch.scala 30:53:@17575.4]
  assign valid_54_59 = io_inValid_59 & _T_38621; // @[Switch.scala 30:36:@17576.4]
  assign _T_38624 = io_inAddr_60 == 6'h36; // @[Switch.scala 30:53:@17578.4]
  assign valid_54_60 = io_inValid_60 & _T_38624; // @[Switch.scala 30:36:@17579.4]
  assign _T_38627 = io_inAddr_61 == 6'h36; // @[Switch.scala 30:53:@17581.4]
  assign valid_54_61 = io_inValid_61 & _T_38627; // @[Switch.scala 30:36:@17582.4]
  assign _T_38630 = io_inAddr_62 == 6'h36; // @[Switch.scala 30:53:@17584.4]
  assign valid_54_62 = io_inValid_62 & _T_38630; // @[Switch.scala 30:36:@17585.4]
  assign _T_38633 = io_inAddr_63 == 6'h36; // @[Switch.scala 30:53:@17587.4]
  assign valid_54_63 = io_inValid_63 & _T_38633; // @[Switch.scala 30:36:@17588.4]
  assign _T_38699 = valid_54_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@17590.4]
  assign _T_38700 = valid_54_61 ? 6'h3d : _T_38699; // @[Mux.scala 31:69:@17591.4]
  assign _T_38701 = valid_54_60 ? 6'h3c : _T_38700; // @[Mux.scala 31:69:@17592.4]
  assign _T_38702 = valid_54_59 ? 6'h3b : _T_38701; // @[Mux.scala 31:69:@17593.4]
  assign _T_38703 = valid_54_58 ? 6'h3a : _T_38702; // @[Mux.scala 31:69:@17594.4]
  assign _T_38704 = valid_54_57 ? 6'h39 : _T_38703; // @[Mux.scala 31:69:@17595.4]
  assign _T_38705 = valid_54_56 ? 6'h38 : _T_38704; // @[Mux.scala 31:69:@17596.4]
  assign _T_38706 = valid_54_55 ? 6'h37 : _T_38705; // @[Mux.scala 31:69:@17597.4]
  assign _T_38707 = valid_54_54 ? 6'h36 : _T_38706; // @[Mux.scala 31:69:@17598.4]
  assign _T_38708 = valid_54_53 ? 6'h35 : _T_38707; // @[Mux.scala 31:69:@17599.4]
  assign _T_38709 = valid_54_52 ? 6'h34 : _T_38708; // @[Mux.scala 31:69:@17600.4]
  assign _T_38710 = valid_54_51 ? 6'h33 : _T_38709; // @[Mux.scala 31:69:@17601.4]
  assign _T_38711 = valid_54_50 ? 6'h32 : _T_38710; // @[Mux.scala 31:69:@17602.4]
  assign _T_38712 = valid_54_49 ? 6'h31 : _T_38711; // @[Mux.scala 31:69:@17603.4]
  assign _T_38713 = valid_54_48 ? 6'h30 : _T_38712; // @[Mux.scala 31:69:@17604.4]
  assign _T_38714 = valid_54_47 ? 6'h2f : _T_38713; // @[Mux.scala 31:69:@17605.4]
  assign _T_38715 = valid_54_46 ? 6'h2e : _T_38714; // @[Mux.scala 31:69:@17606.4]
  assign _T_38716 = valid_54_45 ? 6'h2d : _T_38715; // @[Mux.scala 31:69:@17607.4]
  assign _T_38717 = valid_54_44 ? 6'h2c : _T_38716; // @[Mux.scala 31:69:@17608.4]
  assign _T_38718 = valid_54_43 ? 6'h2b : _T_38717; // @[Mux.scala 31:69:@17609.4]
  assign _T_38719 = valid_54_42 ? 6'h2a : _T_38718; // @[Mux.scala 31:69:@17610.4]
  assign _T_38720 = valid_54_41 ? 6'h29 : _T_38719; // @[Mux.scala 31:69:@17611.4]
  assign _T_38721 = valid_54_40 ? 6'h28 : _T_38720; // @[Mux.scala 31:69:@17612.4]
  assign _T_38722 = valid_54_39 ? 6'h27 : _T_38721; // @[Mux.scala 31:69:@17613.4]
  assign _T_38723 = valid_54_38 ? 6'h26 : _T_38722; // @[Mux.scala 31:69:@17614.4]
  assign _T_38724 = valid_54_37 ? 6'h25 : _T_38723; // @[Mux.scala 31:69:@17615.4]
  assign _T_38725 = valid_54_36 ? 6'h24 : _T_38724; // @[Mux.scala 31:69:@17616.4]
  assign _T_38726 = valid_54_35 ? 6'h23 : _T_38725; // @[Mux.scala 31:69:@17617.4]
  assign _T_38727 = valid_54_34 ? 6'h22 : _T_38726; // @[Mux.scala 31:69:@17618.4]
  assign _T_38728 = valid_54_33 ? 6'h21 : _T_38727; // @[Mux.scala 31:69:@17619.4]
  assign _T_38729 = valid_54_32 ? 6'h20 : _T_38728; // @[Mux.scala 31:69:@17620.4]
  assign _T_38730 = valid_54_31 ? 6'h1f : _T_38729; // @[Mux.scala 31:69:@17621.4]
  assign _T_38731 = valid_54_30 ? 6'h1e : _T_38730; // @[Mux.scala 31:69:@17622.4]
  assign _T_38732 = valid_54_29 ? 6'h1d : _T_38731; // @[Mux.scala 31:69:@17623.4]
  assign _T_38733 = valid_54_28 ? 6'h1c : _T_38732; // @[Mux.scala 31:69:@17624.4]
  assign _T_38734 = valid_54_27 ? 6'h1b : _T_38733; // @[Mux.scala 31:69:@17625.4]
  assign _T_38735 = valid_54_26 ? 6'h1a : _T_38734; // @[Mux.scala 31:69:@17626.4]
  assign _T_38736 = valid_54_25 ? 6'h19 : _T_38735; // @[Mux.scala 31:69:@17627.4]
  assign _T_38737 = valid_54_24 ? 6'h18 : _T_38736; // @[Mux.scala 31:69:@17628.4]
  assign _T_38738 = valid_54_23 ? 6'h17 : _T_38737; // @[Mux.scala 31:69:@17629.4]
  assign _T_38739 = valid_54_22 ? 6'h16 : _T_38738; // @[Mux.scala 31:69:@17630.4]
  assign _T_38740 = valid_54_21 ? 6'h15 : _T_38739; // @[Mux.scala 31:69:@17631.4]
  assign _T_38741 = valid_54_20 ? 6'h14 : _T_38740; // @[Mux.scala 31:69:@17632.4]
  assign _T_38742 = valid_54_19 ? 6'h13 : _T_38741; // @[Mux.scala 31:69:@17633.4]
  assign _T_38743 = valid_54_18 ? 6'h12 : _T_38742; // @[Mux.scala 31:69:@17634.4]
  assign _T_38744 = valid_54_17 ? 6'h11 : _T_38743; // @[Mux.scala 31:69:@17635.4]
  assign _T_38745 = valid_54_16 ? 6'h10 : _T_38744; // @[Mux.scala 31:69:@17636.4]
  assign _T_38746 = valid_54_15 ? 6'hf : _T_38745; // @[Mux.scala 31:69:@17637.4]
  assign _T_38747 = valid_54_14 ? 6'he : _T_38746; // @[Mux.scala 31:69:@17638.4]
  assign _T_38748 = valid_54_13 ? 6'hd : _T_38747; // @[Mux.scala 31:69:@17639.4]
  assign _T_38749 = valid_54_12 ? 6'hc : _T_38748; // @[Mux.scala 31:69:@17640.4]
  assign _T_38750 = valid_54_11 ? 6'hb : _T_38749; // @[Mux.scala 31:69:@17641.4]
  assign _T_38751 = valid_54_10 ? 6'ha : _T_38750; // @[Mux.scala 31:69:@17642.4]
  assign _T_38752 = valid_54_9 ? 6'h9 : _T_38751; // @[Mux.scala 31:69:@17643.4]
  assign _T_38753 = valid_54_8 ? 6'h8 : _T_38752; // @[Mux.scala 31:69:@17644.4]
  assign _T_38754 = valid_54_7 ? 6'h7 : _T_38753; // @[Mux.scala 31:69:@17645.4]
  assign _T_38755 = valid_54_6 ? 6'h6 : _T_38754; // @[Mux.scala 31:69:@17646.4]
  assign _T_38756 = valid_54_5 ? 6'h5 : _T_38755; // @[Mux.scala 31:69:@17647.4]
  assign _T_38757 = valid_54_4 ? 6'h4 : _T_38756; // @[Mux.scala 31:69:@17648.4]
  assign _T_38758 = valid_54_3 ? 6'h3 : _T_38757; // @[Mux.scala 31:69:@17649.4]
  assign _T_38759 = valid_54_2 ? 6'h2 : _T_38758; // @[Mux.scala 31:69:@17650.4]
  assign _T_38760 = valid_54_1 ? 6'h1 : _T_38759; // @[Mux.scala 31:69:@17651.4]
  assign select_54 = valid_54_0 ? 6'h0 : _T_38760; // @[Mux.scala 31:69:@17652.4]
  assign _GEN_3457 = 6'h1 == select_54 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3458 = 6'h2 == select_54 ? io_inData_2 : _GEN_3457; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3459 = 6'h3 == select_54 ? io_inData_3 : _GEN_3458; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3460 = 6'h4 == select_54 ? io_inData_4 : _GEN_3459; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3461 = 6'h5 == select_54 ? io_inData_5 : _GEN_3460; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3462 = 6'h6 == select_54 ? io_inData_6 : _GEN_3461; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3463 = 6'h7 == select_54 ? io_inData_7 : _GEN_3462; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3464 = 6'h8 == select_54 ? io_inData_8 : _GEN_3463; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3465 = 6'h9 == select_54 ? io_inData_9 : _GEN_3464; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3466 = 6'ha == select_54 ? io_inData_10 : _GEN_3465; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3467 = 6'hb == select_54 ? io_inData_11 : _GEN_3466; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3468 = 6'hc == select_54 ? io_inData_12 : _GEN_3467; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3469 = 6'hd == select_54 ? io_inData_13 : _GEN_3468; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3470 = 6'he == select_54 ? io_inData_14 : _GEN_3469; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3471 = 6'hf == select_54 ? io_inData_15 : _GEN_3470; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3472 = 6'h10 == select_54 ? io_inData_16 : _GEN_3471; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3473 = 6'h11 == select_54 ? io_inData_17 : _GEN_3472; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3474 = 6'h12 == select_54 ? io_inData_18 : _GEN_3473; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3475 = 6'h13 == select_54 ? io_inData_19 : _GEN_3474; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3476 = 6'h14 == select_54 ? io_inData_20 : _GEN_3475; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3477 = 6'h15 == select_54 ? io_inData_21 : _GEN_3476; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3478 = 6'h16 == select_54 ? io_inData_22 : _GEN_3477; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3479 = 6'h17 == select_54 ? io_inData_23 : _GEN_3478; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3480 = 6'h18 == select_54 ? io_inData_24 : _GEN_3479; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3481 = 6'h19 == select_54 ? io_inData_25 : _GEN_3480; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3482 = 6'h1a == select_54 ? io_inData_26 : _GEN_3481; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3483 = 6'h1b == select_54 ? io_inData_27 : _GEN_3482; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3484 = 6'h1c == select_54 ? io_inData_28 : _GEN_3483; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3485 = 6'h1d == select_54 ? io_inData_29 : _GEN_3484; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3486 = 6'h1e == select_54 ? io_inData_30 : _GEN_3485; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3487 = 6'h1f == select_54 ? io_inData_31 : _GEN_3486; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3488 = 6'h20 == select_54 ? io_inData_32 : _GEN_3487; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3489 = 6'h21 == select_54 ? io_inData_33 : _GEN_3488; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3490 = 6'h22 == select_54 ? io_inData_34 : _GEN_3489; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3491 = 6'h23 == select_54 ? io_inData_35 : _GEN_3490; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3492 = 6'h24 == select_54 ? io_inData_36 : _GEN_3491; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3493 = 6'h25 == select_54 ? io_inData_37 : _GEN_3492; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3494 = 6'h26 == select_54 ? io_inData_38 : _GEN_3493; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3495 = 6'h27 == select_54 ? io_inData_39 : _GEN_3494; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3496 = 6'h28 == select_54 ? io_inData_40 : _GEN_3495; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3497 = 6'h29 == select_54 ? io_inData_41 : _GEN_3496; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3498 = 6'h2a == select_54 ? io_inData_42 : _GEN_3497; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3499 = 6'h2b == select_54 ? io_inData_43 : _GEN_3498; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3500 = 6'h2c == select_54 ? io_inData_44 : _GEN_3499; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3501 = 6'h2d == select_54 ? io_inData_45 : _GEN_3500; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3502 = 6'h2e == select_54 ? io_inData_46 : _GEN_3501; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3503 = 6'h2f == select_54 ? io_inData_47 : _GEN_3502; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3504 = 6'h30 == select_54 ? io_inData_48 : _GEN_3503; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3505 = 6'h31 == select_54 ? io_inData_49 : _GEN_3504; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3506 = 6'h32 == select_54 ? io_inData_50 : _GEN_3505; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3507 = 6'h33 == select_54 ? io_inData_51 : _GEN_3506; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3508 = 6'h34 == select_54 ? io_inData_52 : _GEN_3507; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3509 = 6'h35 == select_54 ? io_inData_53 : _GEN_3508; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3510 = 6'h36 == select_54 ? io_inData_54 : _GEN_3509; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3511 = 6'h37 == select_54 ? io_inData_55 : _GEN_3510; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3512 = 6'h38 == select_54 ? io_inData_56 : _GEN_3511; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3513 = 6'h39 == select_54 ? io_inData_57 : _GEN_3512; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3514 = 6'h3a == select_54 ? io_inData_58 : _GEN_3513; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3515 = 6'h3b == select_54 ? io_inData_59 : _GEN_3514; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3516 = 6'h3c == select_54 ? io_inData_60 : _GEN_3515; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3517 = 6'h3d == select_54 ? io_inData_61 : _GEN_3516; // @[Switch.scala 33:19:@17654.4]
  assign _GEN_3518 = 6'h3e == select_54 ? io_inData_62 : _GEN_3517; // @[Switch.scala 33:19:@17654.4]
  assign _T_38769 = {valid_54_7,valid_54_6,valid_54_5,valid_54_4,valid_54_3,valid_54_2,valid_54_1,valid_54_0}; // @[Switch.scala 34:32:@17661.4]
  assign _T_38777 = {valid_54_15,valid_54_14,valid_54_13,valid_54_12,valid_54_11,valid_54_10,valid_54_9,valid_54_8,_T_38769}; // @[Switch.scala 34:32:@17669.4]
  assign _T_38784 = {valid_54_23,valid_54_22,valid_54_21,valid_54_20,valid_54_19,valid_54_18,valid_54_17,valid_54_16}; // @[Switch.scala 34:32:@17676.4]
  assign _T_38793 = {valid_54_31,valid_54_30,valid_54_29,valid_54_28,valid_54_27,valid_54_26,valid_54_25,valid_54_24,_T_38784,_T_38777}; // @[Switch.scala 34:32:@17685.4]
  assign _T_38800 = {valid_54_39,valid_54_38,valid_54_37,valid_54_36,valid_54_35,valid_54_34,valid_54_33,valid_54_32}; // @[Switch.scala 34:32:@17692.4]
  assign _T_38808 = {valid_54_47,valid_54_46,valid_54_45,valid_54_44,valid_54_43,valid_54_42,valid_54_41,valid_54_40,_T_38800}; // @[Switch.scala 34:32:@17700.4]
  assign _T_38815 = {valid_54_55,valid_54_54,valid_54_53,valid_54_52,valid_54_51,valid_54_50,valid_54_49,valid_54_48}; // @[Switch.scala 34:32:@17707.4]
  assign _T_38824 = {valid_54_63,valid_54_62,valid_54_61,valid_54_60,valid_54_59,valid_54_58,valid_54_57,valid_54_56,_T_38815,_T_38808}; // @[Switch.scala 34:32:@17716.4]
  assign _T_38825 = {_T_38824,_T_38793}; // @[Switch.scala 34:32:@17717.4]
  assign _T_38829 = io_inAddr_0 == 6'h37; // @[Switch.scala 30:53:@17720.4]
  assign valid_55_0 = io_inValid_0 & _T_38829; // @[Switch.scala 30:36:@17721.4]
  assign _T_38832 = io_inAddr_1 == 6'h37; // @[Switch.scala 30:53:@17723.4]
  assign valid_55_1 = io_inValid_1 & _T_38832; // @[Switch.scala 30:36:@17724.4]
  assign _T_38835 = io_inAddr_2 == 6'h37; // @[Switch.scala 30:53:@17726.4]
  assign valid_55_2 = io_inValid_2 & _T_38835; // @[Switch.scala 30:36:@17727.4]
  assign _T_38838 = io_inAddr_3 == 6'h37; // @[Switch.scala 30:53:@17729.4]
  assign valid_55_3 = io_inValid_3 & _T_38838; // @[Switch.scala 30:36:@17730.4]
  assign _T_38841 = io_inAddr_4 == 6'h37; // @[Switch.scala 30:53:@17732.4]
  assign valid_55_4 = io_inValid_4 & _T_38841; // @[Switch.scala 30:36:@17733.4]
  assign _T_38844 = io_inAddr_5 == 6'h37; // @[Switch.scala 30:53:@17735.4]
  assign valid_55_5 = io_inValid_5 & _T_38844; // @[Switch.scala 30:36:@17736.4]
  assign _T_38847 = io_inAddr_6 == 6'h37; // @[Switch.scala 30:53:@17738.4]
  assign valid_55_6 = io_inValid_6 & _T_38847; // @[Switch.scala 30:36:@17739.4]
  assign _T_38850 = io_inAddr_7 == 6'h37; // @[Switch.scala 30:53:@17741.4]
  assign valid_55_7 = io_inValid_7 & _T_38850; // @[Switch.scala 30:36:@17742.4]
  assign _T_38853 = io_inAddr_8 == 6'h37; // @[Switch.scala 30:53:@17744.4]
  assign valid_55_8 = io_inValid_8 & _T_38853; // @[Switch.scala 30:36:@17745.4]
  assign _T_38856 = io_inAddr_9 == 6'h37; // @[Switch.scala 30:53:@17747.4]
  assign valid_55_9 = io_inValid_9 & _T_38856; // @[Switch.scala 30:36:@17748.4]
  assign _T_38859 = io_inAddr_10 == 6'h37; // @[Switch.scala 30:53:@17750.4]
  assign valid_55_10 = io_inValid_10 & _T_38859; // @[Switch.scala 30:36:@17751.4]
  assign _T_38862 = io_inAddr_11 == 6'h37; // @[Switch.scala 30:53:@17753.4]
  assign valid_55_11 = io_inValid_11 & _T_38862; // @[Switch.scala 30:36:@17754.4]
  assign _T_38865 = io_inAddr_12 == 6'h37; // @[Switch.scala 30:53:@17756.4]
  assign valid_55_12 = io_inValid_12 & _T_38865; // @[Switch.scala 30:36:@17757.4]
  assign _T_38868 = io_inAddr_13 == 6'h37; // @[Switch.scala 30:53:@17759.4]
  assign valid_55_13 = io_inValid_13 & _T_38868; // @[Switch.scala 30:36:@17760.4]
  assign _T_38871 = io_inAddr_14 == 6'h37; // @[Switch.scala 30:53:@17762.4]
  assign valid_55_14 = io_inValid_14 & _T_38871; // @[Switch.scala 30:36:@17763.4]
  assign _T_38874 = io_inAddr_15 == 6'h37; // @[Switch.scala 30:53:@17765.4]
  assign valid_55_15 = io_inValid_15 & _T_38874; // @[Switch.scala 30:36:@17766.4]
  assign _T_38877 = io_inAddr_16 == 6'h37; // @[Switch.scala 30:53:@17768.4]
  assign valid_55_16 = io_inValid_16 & _T_38877; // @[Switch.scala 30:36:@17769.4]
  assign _T_38880 = io_inAddr_17 == 6'h37; // @[Switch.scala 30:53:@17771.4]
  assign valid_55_17 = io_inValid_17 & _T_38880; // @[Switch.scala 30:36:@17772.4]
  assign _T_38883 = io_inAddr_18 == 6'h37; // @[Switch.scala 30:53:@17774.4]
  assign valid_55_18 = io_inValid_18 & _T_38883; // @[Switch.scala 30:36:@17775.4]
  assign _T_38886 = io_inAddr_19 == 6'h37; // @[Switch.scala 30:53:@17777.4]
  assign valid_55_19 = io_inValid_19 & _T_38886; // @[Switch.scala 30:36:@17778.4]
  assign _T_38889 = io_inAddr_20 == 6'h37; // @[Switch.scala 30:53:@17780.4]
  assign valid_55_20 = io_inValid_20 & _T_38889; // @[Switch.scala 30:36:@17781.4]
  assign _T_38892 = io_inAddr_21 == 6'h37; // @[Switch.scala 30:53:@17783.4]
  assign valid_55_21 = io_inValid_21 & _T_38892; // @[Switch.scala 30:36:@17784.4]
  assign _T_38895 = io_inAddr_22 == 6'h37; // @[Switch.scala 30:53:@17786.4]
  assign valid_55_22 = io_inValid_22 & _T_38895; // @[Switch.scala 30:36:@17787.4]
  assign _T_38898 = io_inAddr_23 == 6'h37; // @[Switch.scala 30:53:@17789.4]
  assign valid_55_23 = io_inValid_23 & _T_38898; // @[Switch.scala 30:36:@17790.4]
  assign _T_38901 = io_inAddr_24 == 6'h37; // @[Switch.scala 30:53:@17792.4]
  assign valid_55_24 = io_inValid_24 & _T_38901; // @[Switch.scala 30:36:@17793.4]
  assign _T_38904 = io_inAddr_25 == 6'h37; // @[Switch.scala 30:53:@17795.4]
  assign valid_55_25 = io_inValid_25 & _T_38904; // @[Switch.scala 30:36:@17796.4]
  assign _T_38907 = io_inAddr_26 == 6'h37; // @[Switch.scala 30:53:@17798.4]
  assign valid_55_26 = io_inValid_26 & _T_38907; // @[Switch.scala 30:36:@17799.4]
  assign _T_38910 = io_inAddr_27 == 6'h37; // @[Switch.scala 30:53:@17801.4]
  assign valid_55_27 = io_inValid_27 & _T_38910; // @[Switch.scala 30:36:@17802.4]
  assign _T_38913 = io_inAddr_28 == 6'h37; // @[Switch.scala 30:53:@17804.4]
  assign valid_55_28 = io_inValid_28 & _T_38913; // @[Switch.scala 30:36:@17805.4]
  assign _T_38916 = io_inAddr_29 == 6'h37; // @[Switch.scala 30:53:@17807.4]
  assign valid_55_29 = io_inValid_29 & _T_38916; // @[Switch.scala 30:36:@17808.4]
  assign _T_38919 = io_inAddr_30 == 6'h37; // @[Switch.scala 30:53:@17810.4]
  assign valid_55_30 = io_inValid_30 & _T_38919; // @[Switch.scala 30:36:@17811.4]
  assign _T_38922 = io_inAddr_31 == 6'h37; // @[Switch.scala 30:53:@17813.4]
  assign valid_55_31 = io_inValid_31 & _T_38922; // @[Switch.scala 30:36:@17814.4]
  assign _T_38925 = io_inAddr_32 == 6'h37; // @[Switch.scala 30:53:@17816.4]
  assign valid_55_32 = io_inValid_32 & _T_38925; // @[Switch.scala 30:36:@17817.4]
  assign _T_38928 = io_inAddr_33 == 6'h37; // @[Switch.scala 30:53:@17819.4]
  assign valid_55_33 = io_inValid_33 & _T_38928; // @[Switch.scala 30:36:@17820.4]
  assign _T_38931 = io_inAddr_34 == 6'h37; // @[Switch.scala 30:53:@17822.4]
  assign valid_55_34 = io_inValid_34 & _T_38931; // @[Switch.scala 30:36:@17823.4]
  assign _T_38934 = io_inAddr_35 == 6'h37; // @[Switch.scala 30:53:@17825.4]
  assign valid_55_35 = io_inValid_35 & _T_38934; // @[Switch.scala 30:36:@17826.4]
  assign _T_38937 = io_inAddr_36 == 6'h37; // @[Switch.scala 30:53:@17828.4]
  assign valid_55_36 = io_inValid_36 & _T_38937; // @[Switch.scala 30:36:@17829.4]
  assign _T_38940 = io_inAddr_37 == 6'h37; // @[Switch.scala 30:53:@17831.4]
  assign valid_55_37 = io_inValid_37 & _T_38940; // @[Switch.scala 30:36:@17832.4]
  assign _T_38943 = io_inAddr_38 == 6'h37; // @[Switch.scala 30:53:@17834.4]
  assign valid_55_38 = io_inValid_38 & _T_38943; // @[Switch.scala 30:36:@17835.4]
  assign _T_38946 = io_inAddr_39 == 6'h37; // @[Switch.scala 30:53:@17837.4]
  assign valid_55_39 = io_inValid_39 & _T_38946; // @[Switch.scala 30:36:@17838.4]
  assign _T_38949 = io_inAddr_40 == 6'h37; // @[Switch.scala 30:53:@17840.4]
  assign valid_55_40 = io_inValid_40 & _T_38949; // @[Switch.scala 30:36:@17841.4]
  assign _T_38952 = io_inAddr_41 == 6'h37; // @[Switch.scala 30:53:@17843.4]
  assign valid_55_41 = io_inValid_41 & _T_38952; // @[Switch.scala 30:36:@17844.4]
  assign _T_38955 = io_inAddr_42 == 6'h37; // @[Switch.scala 30:53:@17846.4]
  assign valid_55_42 = io_inValid_42 & _T_38955; // @[Switch.scala 30:36:@17847.4]
  assign _T_38958 = io_inAddr_43 == 6'h37; // @[Switch.scala 30:53:@17849.4]
  assign valid_55_43 = io_inValid_43 & _T_38958; // @[Switch.scala 30:36:@17850.4]
  assign _T_38961 = io_inAddr_44 == 6'h37; // @[Switch.scala 30:53:@17852.4]
  assign valid_55_44 = io_inValid_44 & _T_38961; // @[Switch.scala 30:36:@17853.4]
  assign _T_38964 = io_inAddr_45 == 6'h37; // @[Switch.scala 30:53:@17855.4]
  assign valid_55_45 = io_inValid_45 & _T_38964; // @[Switch.scala 30:36:@17856.4]
  assign _T_38967 = io_inAddr_46 == 6'h37; // @[Switch.scala 30:53:@17858.4]
  assign valid_55_46 = io_inValid_46 & _T_38967; // @[Switch.scala 30:36:@17859.4]
  assign _T_38970 = io_inAddr_47 == 6'h37; // @[Switch.scala 30:53:@17861.4]
  assign valid_55_47 = io_inValid_47 & _T_38970; // @[Switch.scala 30:36:@17862.4]
  assign _T_38973 = io_inAddr_48 == 6'h37; // @[Switch.scala 30:53:@17864.4]
  assign valid_55_48 = io_inValid_48 & _T_38973; // @[Switch.scala 30:36:@17865.4]
  assign _T_38976 = io_inAddr_49 == 6'h37; // @[Switch.scala 30:53:@17867.4]
  assign valid_55_49 = io_inValid_49 & _T_38976; // @[Switch.scala 30:36:@17868.4]
  assign _T_38979 = io_inAddr_50 == 6'h37; // @[Switch.scala 30:53:@17870.4]
  assign valid_55_50 = io_inValid_50 & _T_38979; // @[Switch.scala 30:36:@17871.4]
  assign _T_38982 = io_inAddr_51 == 6'h37; // @[Switch.scala 30:53:@17873.4]
  assign valid_55_51 = io_inValid_51 & _T_38982; // @[Switch.scala 30:36:@17874.4]
  assign _T_38985 = io_inAddr_52 == 6'h37; // @[Switch.scala 30:53:@17876.4]
  assign valid_55_52 = io_inValid_52 & _T_38985; // @[Switch.scala 30:36:@17877.4]
  assign _T_38988 = io_inAddr_53 == 6'h37; // @[Switch.scala 30:53:@17879.4]
  assign valid_55_53 = io_inValid_53 & _T_38988; // @[Switch.scala 30:36:@17880.4]
  assign _T_38991 = io_inAddr_54 == 6'h37; // @[Switch.scala 30:53:@17882.4]
  assign valid_55_54 = io_inValid_54 & _T_38991; // @[Switch.scala 30:36:@17883.4]
  assign _T_38994 = io_inAddr_55 == 6'h37; // @[Switch.scala 30:53:@17885.4]
  assign valid_55_55 = io_inValid_55 & _T_38994; // @[Switch.scala 30:36:@17886.4]
  assign _T_38997 = io_inAddr_56 == 6'h37; // @[Switch.scala 30:53:@17888.4]
  assign valid_55_56 = io_inValid_56 & _T_38997; // @[Switch.scala 30:36:@17889.4]
  assign _T_39000 = io_inAddr_57 == 6'h37; // @[Switch.scala 30:53:@17891.4]
  assign valid_55_57 = io_inValid_57 & _T_39000; // @[Switch.scala 30:36:@17892.4]
  assign _T_39003 = io_inAddr_58 == 6'h37; // @[Switch.scala 30:53:@17894.4]
  assign valid_55_58 = io_inValid_58 & _T_39003; // @[Switch.scala 30:36:@17895.4]
  assign _T_39006 = io_inAddr_59 == 6'h37; // @[Switch.scala 30:53:@17897.4]
  assign valid_55_59 = io_inValid_59 & _T_39006; // @[Switch.scala 30:36:@17898.4]
  assign _T_39009 = io_inAddr_60 == 6'h37; // @[Switch.scala 30:53:@17900.4]
  assign valid_55_60 = io_inValid_60 & _T_39009; // @[Switch.scala 30:36:@17901.4]
  assign _T_39012 = io_inAddr_61 == 6'h37; // @[Switch.scala 30:53:@17903.4]
  assign valid_55_61 = io_inValid_61 & _T_39012; // @[Switch.scala 30:36:@17904.4]
  assign _T_39015 = io_inAddr_62 == 6'h37; // @[Switch.scala 30:53:@17906.4]
  assign valid_55_62 = io_inValid_62 & _T_39015; // @[Switch.scala 30:36:@17907.4]
  assign _T_39018 = io_inAddr_63 == 6'h37; // @[Switch.scala 30:53:@17909.4]
  assign valid_55_63 = io_inValid_63 & _T_39018; // @[Switch.scala 30:36:@17910.4]
  assign _T_39084 = valid_55_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@17912.4]
  assign _T_39085 = valid_55_61 ? 6'h3d : _T_39084; // @[Mux.scala 31:69:@17913.4]
  assign _T_39086 = valid_55_60 ? 6'h3c : _T_39085; // @[Mux.scala 31:69:@17914.4]
  assign _T_39087 = valid_55_59 ? 6'h3b : _T_39086; // @[Mux.scala 31:69:@17915.4]
  assign _T_39088 = valid_55_58 ? 6'h3a : _T_39087; // @[Mux.scala 31:69:@17916.4]
  assign _T_39089 = valid_55_57 ? 6'h39 : _T_39088; // @[Mux.scala 31:69:@17917.4]
  assign _T_39090 = valid_55_56 ? 6'h38 : _T_39089; // @[Mux.scala 31:69:@17918.4]
  assign _T_39091 = valid_55_55 ? 6'h37 : _T_39090; // @[Mux.scala 31:69:@17919.4]
  assign _T_39092 = valid_55_54 ? 6'h36 : _T_39091; // @[Mux.scala 31:69:@17920.4]
  assign _T_39093 = valid_55_53 ? 6'h35 : _T_39092; // @[Mux.scala 31:69:@17921.4]
  assign _T_39094 = valid_55_52 ? 6'h34 : _T_39093; // @[Mux.scala 31:69:@17922.4]
  assign _T_39095 = valid_55_51 ? 6'h33 : _T_39094; // @[Mux.scala 31:69:@17923.4]
  assign _T_39096 = valid_55_50 ? 6'h32 : _T_39095; // @[Mux.scala 31:69:@17924.4]
  assign _T_39097 = valid_55_49 ? 6'h31 : _T_39096; // @[Mux.scala 31:69:@17925.4]
  assign _T_39098 = valid_55_48 ? 6'h30 : _T_39097; // @[Mux.scala 31:69:@17926.4]
  assign _T_39099 = valid_55_47 ? 6'h2f : _T_39098; // @[Mux.scala 31:69:@17927.4]
  assign _T_39100 = valid_55_46 ? 6'h2e : _T_39099; // @[Mux.scala 31:69:@17928.4]
  assign _T_39101 = valid_55_45 ? 6'h2d : _T_39100; // @[Mux.scala 31:69:@17929.4]
  assign _T_39102 = valid_55_44 ? 6'h2c : _T_39101; // @[Mux.scala 31:69:@17930.4]
  assign _T_39103 = valid_55_43 ? 6'h2b : _T_39102; // @[Mux.scala 31:69:@17931.4]
  assign _T_39104 = valid_55_42 ? 6'h2a : _T_39103; // @[Mux.scala 31:69:@17932.4]
  assign _T_39105 = valid_55_41 ? 6'h29 : _T_39104; // @[Mux.scala 31:69:@17933.4]
  assign _T_39106 = valid_55_40 ? 6'h28 : _T_39105; // @[Mux.scala 31:69:@17934.4]
  assign _T_39107 = valid_55_39 ? 6'h27 : _T_39106; // @[Mux.scala 31:69:@17935.4]
  assign _T_39108 = valid_55_38 ? 6'h26 : _T_39107; // @[Mux.scala 31:69:@17936.4]
  assign _T_39109 = valid_55_37 ? 6'h25 : _T_39108; // @[Mux.scala 31:69:@17937.4]
  assign _T_39110 = valid_55_36 ? 6'h24 : _T_39109; // @[Mux.scala 31:69:@17938.4]
  assign _T_39111 = valid_55_35 ? 6'h23 : _T_39110; // @[Mux.scala 31:69:@17939.4]
  assign _T_39112 = valid_55_34 ? 6'h22 : _T_39111; // @[Mux.scala 31:69:@17940.4]
  assign _T_39113 = valid_55_33 ? 6'h21 : _T_39112; // @[Mux.scala 31:69:@17941.4]
  assign _T_39114 = valid_55_32 ? 6'h20 : _T_39113; // @[Mux.scala 31:69:@17942.4]
  assign _T_39115 = valid_55_31 ? 6'h1f : _T_39114; // @[Mux.scala 31:69:@17943.4]
  assign _T_39116 = valid_55_30 ? 6'h1e : _T_39115; // @[Mux.scala 31:69:@17944.4]
  assign _T_39117 = valid_55_29 ? 6'h1d : _T_39116; // @[Mux.scala 31:69:@17945.4]
  assign _T_39118 = valid_55_28 ? 6'h1c : _T_39117; // @[Mux.scala 31:69:@17946.4]
  assign _T_39119 = valid_55_27 ? 6'h1b : _T_39118; // @[Mux.scala 31:69:@17947.4]
  assign _T_39120 = valid_55_26 ? 6'h1a : _T_39119; // @[Mux.scala 31:69:@17948.4]
  assign _T_39121 = valid_55_25 ? 6'h19 : _T_39120; // @[Mux.scala 31:69:@17949.4]
  assign _T_39122 = valid_55_24 ? 6'h18 : _T_39121; // @[Mux.scala 31:69:@17950.4]
  assign _T_39123 = valid_55_23 ? 6'h17 : _T_39122; // @[Mux.scala 31:69:@17951.4]
  assign _T_39124 = valid_55_22 ? 6'h16 : _T_39123; // @[Mux.scala 31:69:@17952.4]
  assign _T_39125 = valid_55_21 ? 6'h15 : _T_39124; // @[Mux.scala 31:69:@17953.4]
  assign _T_39126 = valid_55_20 ? 6'h14 : _T_39125; // @[Mux.scala 31:69:@17954.4]
  assign _T_39127 = valid_55_19 ? 6'h13 : _T_39126; // @[Mux.scala 31:69:@17955.4]
  assign _T_39128 = valid_55_18 ? 6'h12 : _T_39127; // @[Mux.scala 31:69:@17956.4]
  assign _T_39129 = valid_55_17 ? 6'h11 : _T_39128; // @[Mux.scala 31:69:@17957.4]
  assign _T_39130 = valid_55_16 ? 6'h10 : _T_39129; // @[Mux.scala 31:69:@17958.4]
  assign _T_39131 = valid_55_15 ? 6'hf : _T_39130; // @[Mux.scala 31:69:@17959.4]
  assign _T_39132 = valid_55_14 ? 6'he : _T_39131; // @[Mux.scala 31:69:@17960.4]
  assign _T_39133 = valid_55_13 ? 6'hd : _T_39132; // @[Mux.scala 31:69:@17961.4]
  assign _T_39134 = valid_55_12 ? 6'hc : _T_39133; // @[Mux.scala 31:69:@17962.4]
  assign _T_39135 = valid_55_11 ? 6'hb : _T_39134; // @[Mux.scala 31:69:@17963.4]
  assign _T_39136 = valid_55_10 ? 6'ha : _T_39135; // @[Mux.scala 31:69:@17964.4]
  assign _T_39137 = valid_55_9 ? 6'h9 : _T_39136; // @[Mux.scala 31:69:@17965.4]
  assign _T_39138 = valid_55_8 ? 6'h8 : _T_39137; // @[Mux.scala 31:69:@17966.4]
  assign _T_39139 = valid_55_7 ? 6'h7 : _T_39138; // @[Mux.scala 31:69:@17967.4]
  assign _T_39140 = valid_55_6 ? 6'h6 : _T_39139; // @[Mux.scala 31:69:@17968.4]
  assign _T_39141 = valid_55_5 ? 6'h5 : _T_39140; // @[Mux.scala 31:69:@17969.4]
  assign _T_39142 = valid_55_4 ? 6'h4 : _T_39141; // @[Mux.scala 31:69:@17970.4]
  assign _T_39143 = valid_55_3 ? 6'h3 : _T_39142; // @[Mux.scala 31:69:@17971.4]
  assign _T_39144 = valid_55_2 ? 6'h2 : _T_39143; // @[Mux.scala 31:69:@17972.4]
  assign _T_39145 = valid_55_1 ? 6'h1 : _T_39144; // @[Mux.scala 31:69:@17973.4]
  assign select_55 = valid_55_0 ? 6'h0 : _T_39145; // @[Mux.scala 31:69:@17974.4]
  assign _GEN_3521 = 6'h1 == select_55 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3522 = 6'h2 == select_55 ? io_inData_2 : _GEN_3521; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3523 = 6'h3 == select_55 ? io_inData_3 : _GEN_3522; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3524 = 6'h4 == select_55 ? io_inData_4 : _GEN_3523; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3525 = 6'h5 == select_55 ? io_inData_5 : _GEN_3524; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3526 = 6'h6 == select_55 ? io_inData_6 : _GEN_3525; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3527 = 6'h7 == select_55 ? io_inData_7 : _GEN_3526; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3528 = 6'h8 == select_55 ? io_inData_8 : _GEN_3527; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3529 = 6'h9 == select_55 ? io_inData_9 : _GEN_3528; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3530 = 6'ha == select_55 ? io_inData_10 : _GEN_3529; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3531 = 6'hb == select_55 ? io_inData_11 : _GEN_3530; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3532 = 6'hc == select_55 ? io_inData_12 : _GEN_3531; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3533 = 6'hd == select_55 ? io_inData_13 : _GEN_3532; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3534 = 6'he == select_55 ? io_inData_14 : _GEN_3533; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3535 = 6'hf == select_55 ? io_inData_15 : _GEN_3534; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3536 = 6'h10 == select_55 ? io_inData_16 : _GEN_3535; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3537 = 6'h11 == select_55 ? io_inData_17 : _GEN_3536; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3538 = 6'h12 == select_55 ? io_inData_18 : _GEN_3537; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3539 = 6'h13 == select_55 ? io_inData_19 : _GEN_3538; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3540 = 6'h14 == select_55 ? io_inData_20 : _GEN_3539; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3541 = 6'h15 == select_55 ? io_inData_21 : _GEN_3540; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3542 = 6'h16 == select_55 ? io_inData_22 : _GEN_3541; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3543 = 6'h17 == select_55 ? io_inData_23 : _GEN_3542; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3544 = 6'h18 == select_55 ? io_inData_24 : _GEN_3543; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3545 = 6'h19 == select_55 ? io_inData_25 : _GEN_3544; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3546 = 6'h1a == select_55 ? io_inData_26 : _GEN_3545; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3547 = 6'h1b == select_55 ? io_inData_27 : _GEN_3546; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3548 = 6'h1c == select_55 ? io_inData_28 : _GEN_3547; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3549 = 6'h1d == select_55 ? io_inData_29 : _GEN_3548; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3550 = 6'h1e == select_55 ? io_inData_30 : _GEN_3549; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3551 = 6'h1f == select_55 ? io_inData_31 : _GEN_3550; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3552 = 6'h20 == select_55 ? io_inData_32 : _GEN_3551; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3553 = 6'h21 == select_55 ? io_inData_33 : _GEN_3552; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3554 = 6'h22 == select_55 ? io_inData_34 : _GEN_3553; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3555 = 6'h23 == select_55 ? io_inData_35 : _GEN_3554; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3556 = 6'h24 == select_55 ? io_inData_36 : _GEN_3555; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3557 = 6'h25 == select_55 ? io_inData_37 : _GEN_3556; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3558 = 6'h26 == select_55 ? io_inData_38 : _GEN_3557; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3559 = 6'h27 == select_55 ? io_inData_39 : _GEN_3558; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3560 = 6'h28 == select_55 ? io_inData_40 : _GEN_3559; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3561 = 6'h29 == select_55 ? io_inData_41 : _GEN_3560; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3562 = 6'h2a == select_55 ? io_inData_42 : _GEN_3561; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3563 = 6'h2b == select_55 ? io_inData_43 : _GEN_3562; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3564 = 6'h2c == select_55 ? io_inData_44 : _GEN_3563; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3565 = 6'h2d == select_55 ? io_inData_45 : _GEN_3564; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3566 = 6'h2e == select_55 ? io_inData_46 : _GEN_3565; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3567 = 6'h2f == select_55 ? io_inData_47 : _GEN_3566; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3568 = 6'h30 == select_55 ? io_inData_48 : _GEN_3567; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3569 = 6'h31 == select_55 ? io_inData_49 : _GEN_3568; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3570 = 6'h32 == select_55 ? io_inData_50 : _GEN_3569; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3571 = 6'h33 == select_55 ? io_inData_51 : _GEN_3570; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3572 = 6'h34 == select_55 ? io_inData_52 : _GEN_3571; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3573 = 6'h35 == select_55 ? io_inData_53 : _GEN_3572; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3574 = 6'h36 == select_55 ? io_inData_54 : _GEN_3573; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3575 = 6'h37 == select_55 ? io_inData_55 : _GEN_3574; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3576 = 6'h38 == select_55 ? io_inData_56 : _GEN_3575; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3577 = 6'h39 == select_55 ? io_inData_57 : _GEN_3576; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3578 = 6'h3a == select_55 ? io_inData_58 : _GEN_3577; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3579 = 6'h3b == select_55 ? io_inData_59 : _GEN_3578; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3580 = 6'h3c == select_55 ? io_inData_60 : _GEN_3579; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3581 = 6'h3d == select_55 ? io_inData_61 : _GEN_3580; // @[Switch.scala 33:19:@17976.4]
  assign _GEN_3582 = 6'h3e == select_55 ? io_inData_62 : _GEN_3581; // @[Switch.scala 33:19:@17976.4]
  assign _T_39154 = {valid_55_7,valid_55_6,valid_55_5,valid_55_4,valid_55_3,valid_55_2,valid_55_1,valid_55_0}; // @[Switch.scala 34:32:@17983.4]
  assign _T_39162 = {valid_55_15,valid_55_14,valid_55_13,valid_55_12,valid_55_11,valid_55_10,valid_55_9,valid_55_8,_T_39154}; // @[Switch.scala 34:32:@17991.4]
  assign _T_39169 = {valid_55_23,valid_55_22,valid_55_21,valid_55_20,valid_55_19,valid_55_18,valid_55_17,valid_55_16}; // @[Switch.scala 34:32:@17998.4]
  assign _T_39178 = {valid_55_31,valid_55_30,valid_55_29,valid_55_28,valid_55_27,valid_55_26,valid_55_25,valid_55_24,_T_39169,_T_39162}; // @[Switch.scala 34:32:@18007.4]
  assign _T_39185 = {valid_55_39,valid_55_38,valid_55_37,valid_55_36,valid_55_35,valid_55_34,valid_55_33,valid_55_32}; // @[Switch.scala 34:32:@18014.4]
  assign _T_39193 = {valid_55_47,valid_55_46,valid_55_45,valid_55_44,valid_55_43,valid_55_42,valid_55_41,valid_55_40,_T_39185}; // @[Switch.scala 34:32:@18022.4]
  assign _T_39200 = {valid_55_55,valid_55_54,valid_55_53,valid_55_52,valid_55_51,valid_55_50,valid_55_49,valid_55_48}; // @[Switch.scala 34:32:@18029.4]
  assign _T_39209 = {valid_55_63,valid_55_62,valid_55_61,valid_55_60,valid_55_59,valid_55_58,valid_55_57,valid_55_56,_T_39200,_T_39193}; // @[Switch.scala 34:32:@18038.4]
  assign _T_39210 = {_T_39209,_T_39178}; // @[Switch.scala 34:32:@18039.4]
  assign _T_39214 = io_inAddr_0 == 6'h38; // @[Switch.scala 30:53:@18042.4]
  assign valid_56_0 = io_inValid_0 & _T_39214; // @[Switch.scala 30:36:@18043.4]
  assign _T_39217 = io_inAddr_1 == 6'h38; // @[Switch.scala 30:53:@18045.4]
  assign valid_56_1 = io_inValid_1 & _T_39217; // @[Switch.scala 30:36:@18046.4]
  assign _T_39220 = io_inAddr_2 == 6'h38; // @[Switch.scala 30:53:@18048.4]
  assign valid_56_2 = io_inValid_2 & _T_39220; // @[Switch.scala 30:36:@18049.4]
  assign _T_39223 = io_inAddr_3 == 6'h38; // @[Switch.scala 30:53:@18051.4]
  assign valid_56_3 = io_inValid_3 & _T_39223; // @[Switch.scala 30:36:@18052.4]
  assign _T_39226 = io_inAddr_4 == 6'h38; // @[Switch.scala 30:53:@18054.4]
  assign valid_56_4 = io_inValid_4 & _T_39226; // @[Switch.scala 30:36:@18055.4]
  assign _T_39229 = io_inAddr_5 == 6'h38; // @[Switch.scala 30:53:@18057.4]
  assign valid_56_5 = io_inValid_5 & _T_39229; // @[Switch.scala 30:36:@18058.4]
  assign _T_39232 = io_inAddr_6 == 6'h38; // @[Switch.scala 30:53:@18060.4]
  assign valid_56_6 = io_inValid_6 & _T_39232; // @[Switch.scala 30:36:@18061.4]
  assign _T_39235 = io_inAddr_7 == 6'h38; // @[Switch.scala 30:53:@18063.4]
  assign valid_56_7 = io_inValid_7 & _T_39235; // @[Switch.scala 30:36:@18064.4]
  assign _T_39238 = io_inAddr_8 == 6'h38; // @[Switch.scala 30:53:@18066.4]
  assign valid_56_8 = io_inValid_8 & _T_39238; // @[Switch.scala 30:36:@18067.4]
  assign _T_39241 = io_inAddr_9 == 6'h38; // @[Switch.scala 30:53:@18069.4]
  assign valid_56_9 = io_inValid_9 & _T_39241; // @[Switch.scala 30:36:@18070.4]
  assign _T_39244 = io_inAddr_10 == 6'h38; // @[Switch.scala 30:53:@18072.4]
  assign valid_56_10 = io_inValid_10 & _T_39244; // @[Switch.scala 30:36:@18073.4]
  assign _T_39247 = io_inAddr_11 == 6'h38; // @[Switch.scala 30:53:@18075.4]
  assign valid_56_11 = io_inValid_11 & _T_39247; // @[Switch.scala 30:36:@18076.4]
  assign _T_39250 = io_inAddr_12 == 6'h38; // @[Switch.scala 30:53:@18078.4]
  assign valid_56_12 = io_inValid_12 & _T_39250; // @[Switch.scala 30:36:@18079.4]
  assign _T_39253 = io_inAddr_13 == 6'h38; // @[Switch.scala 30:53:@18081.4]
  assign valid_56_13 = io_inValid_13 & _T_39253; // @[Switch.scala 30:36:@18082.4]
  assign _T_39256 = io_inAddr_14 == 6'h38; // @[Switch.scala 30:53:@18084.4]
  assign valid_56_14 = io_inValid_14 & _T_39256; // @[Switch.scala 30:36:@18085.4]
  assign _T_39259 = io_inAddr_15 == 6'h38; // @[Switch.scala 30:53:@18087.4]
  assign valid_56_15 = io_inValid_15 & _T_39259; // @[Switch.scala 30:36:@18088.4]
  assign _T_39262 = io_inAddr_16 == 6'h38; // @[Switch.scala 30:53:@18090.4]
  assign valid_56_16 = io_inValid_16 & _T_39262; // @[Switch.scala 30:36:@18091.4]
  assign _T_39265 = io_inAddr_17 == 6'h38; // @[Switch.scala 30:53:@18093.4]
  assign valid_56_17 = io_inValid_17 & _T_39265; // @[Switch.scala 30:36:@18094.4]
  assign _T_39268 = io_inAddr_18 == 6'h38; // @[Switch.scala 30:53:@18096.4]
  assign valid_56_18 = io_inValid_18 & _T_39268; // @[Switch.scala 30:36:@18097.4]
  assign _T_39271 = io_inAddr_19 == 6'h38; // @[Switch.scala 30:53:@18099.4]
  assign valid_56_19 = io_inValid_19 & _T_39271; // @[Switch.scala 30:36:@18100.4]
  assign _T_39274 = io_inAddr_20 == 6'h38; // @[Switch.scala 30:53:@18102.4]
  assign valid_56_20 = io_inValid_20 & _T_39274; // @[Switch.scala 30:36:@18103.4]
  assign _T_39277 = io_inAddr_21 == 6'h38; // @[Switch.scala 30:53:@18105.4]
  assign valid_56_21 = io_inValid_21 & _T_39277; // @[Switch.scala 30:36:@18106.4]
  assign _T_39280 = io_inAddr_22 == 6'h38; // @[Switch.scala 30:53:@18108.4]
  assign valid_56_22 = io_inValid_22 & _T_39280; // @[Switch.scala 30:36:@18109.4]
  assign _T_39283 = io_inAddr_23 == 6'h38; // @[Switch.scala 30:53:@18111.4]
  assign valid_56_23 = io_inValid_23 & _T_39283; // @[Switch.scala 30:36:@18112.4]
  assign _T_39286 = io_inAddr_24 == 6'h38; // @[Switch.scala 30:53:@18114.4]
  assign valid_56_24 = io_inValid_24 & _T_39286; // @[Switch.scala 30:36:@18115.4]
  assign _T_39289 = io_inAddr_25 == 6'h38; // @[Switch.scala 30:53:@18117.4]
  assign valid_56_25 = io_inValid_25 & _T_39289; // @[Switch.scala 30:36:@18118.4]
  assign _T_39292 = io_inAddr_26 == 6'h38; // @[Switch.scala 30:53:@18120.4]
  assign valid_56_26 = io_inValid_26 & _T_39292; // @[Switch.scala 30:36:@18121.4]
  assign _T_39295 = io_inAddr_27 == 6'h38; // @[Switch.scala 30:53:@18123.4]
  assign valid_56_27 = io_inValid_27 & _T_39295; // @[Switch.scala 30:36:@18124.4]
  assign _T_39298 = io_inAddr_28 == 6'h38; // @[Switch.scala 30:53:@18126.4]
  assign valid_56_28 = io_inValid_28 & _T_39298; // @[Switch.scala 30:36:@18127.4]
  assign _T_39301 = io_inAddr_29 == 6'h38; // @[Switch.scala 30:53:@18129.4]
  assign valid_56_29 = io_inValid_29 & _T_39301; // @[Switch.scala 30:36:@18130.4]
  assign _T_39304 = io_inAddr_30 == 6'h38; // @[Switch.scala 30:53:@18132.4]
  assign valid_56_30 = io_inValid_30 & _T_39304; // @[Switch.scala 30:36:@18133.4]
  assign _T_39307 = io_inAddr_31 == 6'h38; // @[Switch.scala 30:53:@18135.4]
  assign valid_56_31 = io_inValid_31 & _T_39307; // @[Switch.scala 30:36:@18136.4]
  assign _T_39310 = io_inAddr_32 == 6'h38; // @[Switch.scala 30:53:@18138.4]
  assign valid_56_32 = io_inValid_32 & _T_39310; // @[Switch.scala 30:36:@18139.4]
  assign _T_39313 = io_inAddr_33 == 6'h38; // @[Switch.scala 30:53:@18141.4]
  assign valid_56_33 = io_inValid_33 & _T_39313; // @[Switch.scala 30:36:@18142.4]
  assign _T_39316 = io_inAddr_34 == 6'h38; // @[Switch.scala 30:53:@18144.4]
  assign valid_56_34 = io_inValid_34 & _T_39316; // @[Switch.scala 30:36:@18145.4]
  assign _T_39319 = io_inAddr_35 == 6'h38; // @[Switch.scala 30:53:@18147.4]
  assign valid_56_35 = io_inValid_35 & _T_39319; // @[Switch.scala 30:36:@18148.4]
  assign _T_39322 = io_inAddr_36 == 6'h38; // @[Switch.scala 30:53:@18150.4]
  assign valid_56_36 = io_inValid_36 & _T_39322; // @[Switch.scala 30:36:@18151.4]
  assign _T_39325 = io_inAddr_37 == 6'h38; // @[Switch.scala 30:53:@18153.4]
  assign valid_56_37 = io_inValid_37 & _T_39325; // @[Switch.scala 30:36:@18154.4]
  assign _T_39328 = io_inAddr_38 == 6'h38; // @[Switch.scala 30:53:@18156.4]
  assign valid_56_38 = io_inValid_38 & _T_39328; // @[Switch.scala 30:36:@18157.4]
  assign _T_39331 = io_inAddr_39 == 6'h38; // @[Switch.scala 30:53:@18159.4]
  assign valid_56_39 = io_inValid_39 & _T_39331; // @[Switch.scala 30:36:@18160.4]
  assign _T_39334 = io_inAddr_40 == 6'h38; // @[Switch.scala 30:53:@18162.4]
  assign valid_56_40 = io_inValid_40 & _T_39334; // @[Switch.scala 30:36:@18163.4]
  assign _T_39337 = io_inAddr_41 == 6'h38; // @[Switch.scala 30:53:@18165.4]
  assign valid_56_41 = io_inValid_41 & _T_39337; // @[Switch.scala 30:36:@18166.4]
  assign _T_39340 = io_inAddr_42 == 6'h38; // @[Switch.scala 30:53:@18168.4]
  assign valid_56_42 = io_inValid_42 & _T_39340; // @[Switch.scala 30:36:@18169.4]
  assign _T_39343 = io_inAddr_43 == 6'h38; // @[Switch.scala 30:53:@18171.4]
  assign valid_56_43 = io_inValid_43 & _T_39343; // @[Switch.scala 30:36:@18172.4]
  assign _T_39346 = io_inAddr_44 == 6'h38; // @[Switch.scala 30:53:@18174.4]
  assign valid_56_44 = io_inValid_44 & _T_39346; // @[Switch.scala 30:36:@18175.4]
  assign _T_39349 = io_inAddr_45 == 6'h38; // @[Switch.scala 30:53:@18177.4]
  assign valid_56_45 = io_inValid_45 & _T_39349; // @[Switch.scala 30:36:@18178.4]
  assign _T_39352 = io_inAddr_46 == 6'h38; // @[Switch.scala 30:53:@18180.4]
  assign valid_56_46 = io_inValid_46 & _T_39352; // @[Switch.scala 30:36:@18181.4]
  assign _T_39355 = io_inAddr_47 == 6'h38; // @[Switch.scala 30:53:@18183.4]
  assign valid_56_47 = io_inValid_47 & _T_39355; // @[Switch.scala 30:36:@18184.4]
  assign _T_39358 = io_inAddr_48 == 6'h38; // @[Switch.scala 30:53:@18186.4]
  assign valid_56_48 = io_inValid_48 & _T_39358; // @[Switch.scala 30:36:@18187.4]
  assign _T_39361 = io_inAddr_49 == 6'h38; // @[Switch.scala 30:53:@18189.4]
  assign valid_56_49 = io_inValid_49 & _T_39361; // @[Switch.scala 30:36:@18190.4]
  assign _T_39364 = io_inAddr_50 == 6'h38; // @[Switch.scala 30:53:@18192.4]
  assign valid_56_50 = io_inValid_50 & _T_39364; // @[Switch.scala 30:36:@18193.4]
  assign _T_39367 = io_inAddr_51 == 6'h38; // @[Switch.scala 30:53:@18195.4]
  assign valid_56_51 = io_inValid_51 & _T_39367; // @[Switch.scala 30:36:@18196.4]
  assign _T_39370 = io_inAddr_52 == 6'h38; // @[Switch.scala 30:53:@18198.4]
  assign valid_56_52 = io_inValid_52 & _T_39370; // @[Switch.scala 30:36:@18199.4]
  assign _T_39373 = io_inAddr_53 == 6'h38; // @[Switch.scala 30:53:@18201.4]
  assign valid_56_53 = io_inValid_53 & _T_39373; // @[Switch.scala 30:36:@18202.4]
  assign _T_39376 = io_inAddr_54 == 6'h38; // @[Switch.scala 30:53:@18204.4]
  assign valid_56_54 = io_inValid_54 & _T_39376; // @[Switch.scala 30:36:@18205.4]
  assign _T_39379 = io_inAddr_55 == 6'h38; // @[Switch.scala 30:53:@18207.4]
  assign valid_56_55 = io_inValid_55 & _T_39379; // @[Switch.scala 30:36:@18208.4]
  assign _T_39382 = io_inAddr_56 == 6'h38; // @[Switch.scala 30:53:@18210.4]
  assign valid_56_56 = io_inValid_56 & _T_39382; // @[Switch.scala 30:36:@18211.4]
  assign _T_39385 = io_inAddr_57 == 6'h38; // @[Switch.scala 30:53:@18213.4]
  assign valid_56_57 = io_inValid_57 & _T_39385; // @[Switch.scala 30:36:@18214.4]
  assign _T_39388 = io_inAddr_58 == 6'h38; // @[Switch.scala 30:53:@18216.4]
  assign valid_56_58 = io_inValid_58 & _T_39388; // @[Switch.scala 30:36:@18217.4]
  assign _T_39391 = io_inAddr_59 == 6'h38; // @[Switch.scala 30:53:@18219.4]
  assign valid_56_59 = io_inValid_59 & _T_39391; // @[Switch.scala 30:36:@18220.4]
  assign _T_39394 = io_inAddr_60 == 6'h38; // @[Switch.scala 30:53:@18222.4]
  assign valid_56_60 = io_inValid_60 & _T_39394; // @[Switch.scala 30:36:@18223.4]
  assign _T_39397 = io_inAddr_61 == 6'h38; // @[Switch.scala 30:53:@18225.4]
  assign valid_56_61 = io_inValid_61 & _T_39397; // @[Switch.scala 30:36:@18226.4]
  assign _T_39400 = io_inAddr_62 == 6'h38; // @[Switch.scala 30:53:@18228.4]
  assign valid_56_62 = io_inValid_62 & _T_39400; // @[Switch.scala 30:36:@18229.4]
  assign _T_39403 = io_inAddr_63 == 6'h38; // @[Switch.scala 30:53:@18231.4]
  assign valid_56_63 = io_inValid_63 & _T_39403; // @[Switch.scala 30:36:@18232.4]
  assign _T_39469 = valid_56_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@18234.4]
  assign _T_39470 = valid_56_61 ? 6'h3d : _T_39469; // @[Mux.scala 31:69:@18235.4]
  assign _T_39471 = valid_56_60 ? 6'h3c : _T_39470; // @[Mux.scala 31:69:@18236.4]
  assign _T_39472 = valid_56_59 ? 6'h3b : _T_39471; // @[Mux.scala 31:69:@18237.4]
  assign _T_39473 = valid_56_58 ? 6'h3a : _T_39472; // @[Mux.scala 31:69:@18238.4]
  assign _T_39474 = valid_56_57 ? 6'h39 : _T_39473; // @[Mux.scala 31:69:@18239.4]
  assign _T_39475 = valid_56_56 ? 6'h38 : _T_39474; // @[Mux.scala 31:69:@18240.4]
  assign _T_39476 = valid_56_55 ? 6'h37 : _T_39475; // @[Mux.scala 31:69:@18241.4]
  assign _T_39477 = valid_56_54 ? 6'h36 : _T_39476; // @[Mux.scala 31:69:@18242.4]
  assign _T_39478 = valid_56_53 ? 6'h35 : _T_39477; // @[Mux.scala 31:69:@18243.4]
  assign _T_39479 = valid_56_52 ? 6'h34 : _T_39478; // @[Mux.scala 31:69:@18244.4]
  assign _T_39480 = valid_56_51 ? 6'h33 : _T_39479; // @[Mux.scala 31:69:@18245.4]
  assign _T_39481 = valid_56_50 ? 6'h32 : _T_39480; // @[Mux.scala 31:69:@18246.4]
  assign _T_39482 = valid_56_49 ? 6'h31 : _T_39481; // @[Mux.scala 31:69:@18247.4]
  assign _T_39483 = valid_56_48 ? 6'h30 : _T_39482; // @[Mux.scala 31:69:@18248.4]
  assign _T_39484 = valid_56_47 ? 6'h2f : _T_39483; // @[Mux.scala 31:69:@18249.4]
  assign _T_39485 = valid_56_46 ? 6'h2e : _T_39484; // @[Mux.scala 31:69:@18250.4]
  assign _T_39486 = valid_56_45 ? 6'h2d : _T_39485; // @[Mux.scala 31:69:@18251.4]
  assign _T_39487 = valid_56_44 ? 6'h2c : _T_39486; // @[Mux.scala 31:69:@18252.4]
  assign _T_39488 = valid_56_43 ? 6'h2b : _T_39487; // @[Mux.scala 31:69:@18253.4]
  assign _T_39489 = valid_56_42 ? 6'h2a : _T_39488; // @[Mux.scala 31:69:@18254.4]
  assign _T_39490 = valid_56_41 ? 6'h29 : _T_39489; // @[Mux.scala 31:69:@18255.4]
  assign _T_39491 = valid_56_40 ? 6'h28 : _T_39490; // @[Mux.scala 31:69:@18256.4]
  assign _T_39492 = valid_56_39 ? 6'h27 : _T_39491; // @[Mux.scala 31:69:@18257.4]
  assign _T_39493 = valid_56_38 ? 6'h26 : _T_39492; // @[Mux.scala 31:69:@18258.4]
  assign _T_39494 = valid_56_37 ? 6'h25 : _T_39493; // @[Mux.scala 31:69:@18259.4]
  assign _T_39495 = valid_56_36 ? 6'h24 : _T_39494; // @[Mux.scala 31:69:@18260.4]
  assign _T_39496 = valid_56_35 ? 6'h23 : _T_39495; // @[Mux.scala 31:69:@18261.4]
  assign _T_39497 = valid_56_34 ? 6'h22 : _T_39496; // @[Mux.scala 31:69:@18262.4]
  assign _T_39498 = valid_56_33 ? 6'h21 : _T_39497; // @[Mux.scala 31:69:@18263.4]
  assign _T_39499 = valid_56_32 ? 6'h20 : _T_39498; // @[Mux.scala 31:69:@18264.4]
  assign _T_39500 = valid_56_31 ? 6'h1f : _T_39499; // @[Mux.scala 31:69:@18265.4]
  assign _T_39501 = valid_56_30 ? 6'h1e : _T_39500; // @[Mux.scala 31:69:@18266.4]
  assign _T_39502 = valid_56_29 ? 6'h1d : _T_39501; // @[Mux.scala 31:69:@18267.4]
  assign _T_39503 = valid_56_28 ? 6'h1c : _T_39502; // @[Mux.scala 31:69:@18268.4]
  assign _T_39504 = valid_56_27 ? 6'h1b : _T_39503; // @[Mux.scala 31:69:@18269.4]
  assign _T_39505 = valid_56_26 ? 6'h1a : _T_39504; // @[Mux.scala 31:69:@18270.4]
  assign _T_39506 = valid_56_25 ? 6'h19 : _T_39505; // @[Mux.scala 31:69:@18271.4]
  assign _T_39507 = valid_56_24 ? 6'h18 : _T_39506; // @[Mux.scala 31:69:@18272.4]
  assign _T_39508 = valid_56_23 ? 6'h17 : _T_39507; // @[Mux.scala 31:69:@18273.4]
  assign _T_39509 = valid_56_22 ? 6'h16 : _T_39508; // @[Mux.scala 31:69:@18274.4]
  assign _T_39510 = valid_56_21 ? 6'h15 : _T_39509; // @[Mux.scala 31:69:@18275.4]
  assign _T_39511 = valid_56_20 ? 6'h14 : _T_39510; // @[Mux.scala 31:69:@18276.4]
  assign _T_39512 = valid_56_19 ? 6'h13 : _T_39511; // @[Mux.scala 31:69:@18277.4]
  assign _T_39513 = valid_56_18 ? 6'h12 : _T_39512; // @[Mux.scala 31:69:@18278.4]
  assign _T_39514 = valid_56_17 ? 6'h11 : _T_39513; // @[Mux.scala 31:69:@18279.4]
  assign _T_39515 = valid_56_16 ? 6'h10 : _T_39514; // @[Mux.scala 31:69:@18280.4]
  assign _T_39516 = valid_56_15 ? 6'hf : _T_39515; // @[Mux.scala 31:69:@18281.4]
  assign _T_39517 = valid_56_14 ? 6'he : _T_39516; // @[Mux.scala 31:69:@18282.4]
  assign _T_39518 = valid_56_13 ? 6'hd : _T_39517; // @[Mux.scala 31:69:@18283.4]
  assign _T_39519 = valid_56_12 ? 6'hc : _T_39518; // @[Mux.scala 31:69:@18284.4]
  assign _T_39520 = valid_56_11 ? 6'hb : _T_39519; // @[Mux.scala 31:69:@18285.4]
  assign _T_39521 = valid_56_10 ? 6'ha : _T_39520; // @[Mux.scala 31:69:@18286.4]
  assign _T_39522 = valid_56_9 ? 6'h9 : _T_39521; // @[Mux.scala 31:69:@18287.4]
  assign _T_39523 = valid_56_8 ? 6'h8 : _T_39522; // @[Mux.scala 31:69:@18288.4]
  assign _T_39524 = valid_56_7 ? 6'h7 : _T_39523; // @[Mux.scala 31:69:@18289.4]
  assign _T_39525 = valid_56_6 ? 6'h6 : _T_39524; // @[Mux.scala 31:69:@18290.4]
  assign _T_39526 = valid_56_5 ? 6'h5 : _T_39525; // @[Mux.scala 31:69:@18291.4]
  assign _T_39527 = valid_56_4 ? 6'h4 : _T_39526; // @[Mux.scala 31:69:@18292.4]
  assign _T_39528 = valid_56_3 ? 6'h3 : _T_39527; // @[Mux.scala 31:69:@18293.4]
  assign _T_39529 = valid_56_2 ? 6'h2 : _T_39528; // @[Mux.scala 31:69:@18294.4]
  assign _T_39530 = valid_56_1 ? 6'h1 : _T_39529; // @[Mux.scala 31:69:@18295.4]
  assign select_56 = valid_56_0 ? 6'h0 : _T_39530; // @[Mux.scala 31:69:@18296.4]
  assign _GEN_3585 = 6'h1 == select_56 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3586 = 6'h2 == select_56 ? io_inData_2 : _GEN_3585; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3587 = 6'h3 == select_56 ? io_inData_3 : _GEN_3586; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3588 = 6'h4 == select_56 ? io_inData_4 : _GEN_3587; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3589 = 6'h5 == select_56 ? io_inData_5 : _GEN_3588; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3590 = 6'h6 == select_56 ? io_inData_6 : _GEN_3589; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3591 = 6'h7 == select_56 ? io_inData_7 : _GEN_3590; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3592 = 6'h8 == select_56 ? io_inData_8 : _GEN_3591; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3593 = 6'h9 == select_56 ? io_inData_9 : _GEN_3592; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3594 = 6'ha == select_56 ? io_inData_10 : _GEN_3593; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3595 = 6'hb == select_56 ? io_inData_11 : _GEN_3594; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3596 = 6'hc == select_56 ? io_inData_12 : _GEN_3595; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3597 = 6'hd == select_56 ? io_inData_13 : _GEN_3596; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3598 = 6'he == select_56 ? io_inData_14 : _GEN_3597; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3599 = 6'hf == select_56 ? io_inData_15 : _GEN_3598; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3600 = 6'h10 == select_56 ? io_inData_16 : _GEN_3599; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3601 = 6'h11 == select_56 ? io_inData_17 : _GEN_3600; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3602 = 6'h12 == select_56 ? io_inData_18 : _GEN_3601; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3603 = 6'h13 == select_56 ? io_inData_19 : _GEN_3602; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3604 = 6'h14 == select_56 ? io_inData_20 : _GEN_3603; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3605 = 6'h15 == select_56 ? io_inData_21 : _GEN_3604; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3606 = 6'h16 == select_56 ? io_inData_22 : _GEN_3605; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3607 = 6'h17 == select_56 ? io_inData_23 : _GEN_3606; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3608 = 6'h18 == select_56 ? io_inData_24 : _GEN_3607; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3609 = 6'h19 == select_56 ? io_inData_25 : _GEN_3608; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3610 = 6'h1a == select_56 ? io_inData_26 : _GEN_3609; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3611 = 6'h1b == select_56 ? io_inData_27 : _GEN_3610; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3612 = 6'h1c == select_56 ? io_inData_28 : _GEN_3611; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3613 = 6'h1d == select_56 ? io_inData_29 : _GEN_3612; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3614 = 6'h1e == select_56 ? io_inData_30 : _GEN_3613; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3615 = 6'h1f == select_56 ? io_inData_31 : _GEN_3614; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3616 = 6'h20 == select_56 ? io_inData_32 : _GEN_3615; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3617 = 6'h21 == select_56 ? io_inData_33 : _GEN_3616; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3618 = 6'h22 == select_56 ? io_inData_34 : _GEN_3617; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3619 = 6'h23 == select_56 ? io_inData_35 : _GEN_3618; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3620 = 6'h24 == select_56 ? io_inData_36 : _GEN_3619; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3621 = 6'h25 == select_56 ? io_inData_37 : _GEN_3620; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3622 = 6'h26 == select_56 ? io_inData_38 : _GEN_3621; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3623 = 6'h27 == select_56 ? io_inData_39 : _GEN_3622; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3624 = 6'h28 == select_56 ? io_inData_40 : _GEN_3623; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3625 = 6'h29 == select_56 ? io_inData_41 : _GEN_3624; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3626 = 6'h2a == select_56 ? io_inData_42 : _GEN_3625; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3627 = 6'h2b == select_56 ? io_inData_43 : _GEN_3626; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3628 = 6'h2c == select_56 ? io_inData_44 : _GEN_3627; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3629 = 6'h2d == select_56 ? io_inData_45 : _GEN_3628; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3630 = 6'h2e == select_56 ? io_inData_46 : _GEN_3629; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3631 = 6'h2f == select_56 ? io_inData_47 : _GEN_3630; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3632 = 6'h30 == select_56 ? io_inData_48 : _GEN_3631; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3633 = 6'h31 == select_56 ? io_inData_49 : _GEN_3632; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3634 = 6'h32 == select_56 ? io_inData_50 : _GEN_3633; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3635 = 6'h33 == select_56 ? io_inData_51 : _GEN_3634; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3636 = 6'h34 == select_56 ? io_inData_52 : _GEN_3635; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3637 = 6'h35 == select_56 ? io_inData_53 : _GEN_3636; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3638 = 6'h36 == select_56 ? io_inData_54 : _GEN_3637; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3639 = 6'h37 == select_56 ? io_inData_55 : _GEN_3638; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3640 = 6'h38 == select_56 ? io_inData_56 : _GEN_3639; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3641 = 6'h39 == select_56 ? io_inData_57 : _GEN_3640; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3642 = 6'h3a == select_56 ? io_inData_58 : _GEN_3641; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3643 = 6'h3b == select_56 ? io_inData_59 : _GEN_3642; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3644 = 6'h3c == select_56 ? io_inData_60 : _GEN_3643; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3645 = 6'h3d == select_56 ? io_inData_61 : _GEN_3644; // @[Switch.scala 33:19:@18298.4]
  assign _GEN_3646 = 6'h3e == select_56 ? io_inData_62 : _GEN_3645; // @[Switch.scala 33:19:@18298.4]
  assign _T_39539 = {valid_56_7,valid_56_6,valid_56_5,valid_56_4,valid_56_3,valid_56_2,valid_56_1,valid_56_0}; // @[Switch.scala 34:32:@18305.4]
  assign _T_39547 = {valid_56_15,valid_56_14,valid_56_13,valid_56_12,valid_56_11,valid_56_10,valid_56_9,valid_56_8,_T_39539}; // @[Switch.scala 34:32:@18313.4]
  assign _T_39554 = {valid_56_23,valid_56_22,valid_56_21,valid_56_20,valid_56_19,valid_56_18,valid_56_17,valid_56_16}; // @[Switch.scala 34:32:@18320.4]
  assign _T_39563 = {valid_56_31,valid_56_30,valid_56_29,valid_56_28,valid_56_27,valid_56_26,valid_56_25,valid_56_24,_T_39554,_T_39547}; // @[Switch.scala 34:32:@18329.4]
  assign _T_39570 = {valid_56_39,valid_56_38,valid_56_37,valid_56_36,valid_56_35,valid_56_34,valid_56_33,valid_56_32}; // @[Switch.scala 34:32:@18336.4]
  assign _T_39578 = {valid_56_47,valid_56_46,valid_56_45,valid_56_44,valid_56_43,valid_56_42,valid_56_41,valid_56_40,_T_39570}; // @[Switch.scala 34:32:@18344.4]
  assign _T_39585 = {valid_56_55,valid_56_54,valid_56_53,valid_56_52,valid_56_51,valid_56_50,valid_56_49,valid_56_48}; // @[Switch.scala 34:32:@18351.4]
  assign _T_39594 = {valid_56_63,valid_56_62,valid_56_61,valid_56_60,valid_56_59,valid_56_58,valid_56_57,valid_56_56,_T_39585,_T_39578}; // @[Switch.scala 34:32:@18360.4]
  assign _T_39595 = {_T_39594,_T_39563}; // @[Switch.scala 34:32:@18361.4]
  assign _T_39599 = io_inAddr_0 == 6'h39; // @[Switch.scala 30:53:@18364.4]
  assign valid_57_0 = io_inValid_0 & _T_39599; // @[Switch.scala 30:36:@18365.4]
  assign _T_39602 = io_inAddr_1 == 6'h39; // @[Switch.scala 30:53:@18367.4]
  assign valid_57_1 = io_inValid_1 & _T_39602; // @[Switch.scala 30:36:@18368.4]
  assign _T_39605 = io_inAddr_2 == 6'h39; // @[Switch.scala 30:53:@18370.4]
  assign valid_57_2 = io_inValid_2 & _T_39605; // @[Switch.scala 30:36:@18371.4]
  assign _T_39608 = io_inAddr_3 == 6'h39; // @[Switch.scala 30:53:@18373.4]
  assign valid_57_3 = io_inValid_3 & _T_39608; // @[Switch.scala 30:36:@18374.4]
  assign _T_39611 = io_inAddr_4 == 6'h39; // @[Switch.scala 30:53:@18376.4]
  assign valid_57_4 = io_inValid_4 & _T_39611; // @[Switch.scala 30:36:@18377.4]
  assign _T_39614 = io_inAddr_5 == 6'h39; // @[Switch.scala 30:53:@18379.4]
  assign valid_57_5 = io_inValid_5 & _T_39614; // @[Switch.scala 30:36:@18380.4]
  assign _T_39617 = io_inAddr_6 == 6'h39; // @[Switch.scala 30:53:@18382.4]
  assign valid_57_6 = io_inValid_6 & _T_39617; // @[Switch.scala 30:36:@18383.4]
  assign _T_39620 = io_inAddr_7 == 6'h39; // @[Switch.scala 30:53:@18385.4]
  assign valid_57_7 = io_inValid_7 & _T_39620; // @[Switch.scala 30:36:@18386.4]
  assign _T_39623 = io_inAddr_8 == 6'h39; // @[Switch.scala 30:53:@18388.4]
  assign valid_57_8 = io_inValid_8 & _T_39623; // @[Switch.scala 30:36:@18389.4]
  assign _T_39626 = io_inAddr_9 == 6'h39; // @[Switch.scala 30:53:@18391.4]
  assign valid_57_9 = io_inValid_9 & _T_39626; // @[Switch.scala 30:36:@18392.4]
  assign _T_39629 = io_inAddr_10 == 6'h39; // @[Switch.scala 30:53:@18394.4]
  assign valid_57_10 = io_inValid_10 & _T_39629; // @[Switch.scala 30:36:@18395.4]
  assign _T_39632 = io_inAddr_11 == 6'h39; // @[Switch.scala 30:53:@18397.4]
  assign valid_57_11 = io_inValid_11 & _T_39632; // @[Switch.scala 30:36:@18398.4]
  assign _T_39635 = io_inAddr_12 == 6'h39; // @[Switch.scala 30:53:@18400.4]
  assign valid_57_12 = io_inValid_12 & _T_39635; // @[Switch.scala 30:36:@18401.4]
  assign _T_39638 = io_inAddr_13 == 6'h39; // @[Switch.scala 30:53:@18403.4]
  assign valid_57_13 = io_inValid_13 & _T_39638; // @[Switch.scala 30:36:@18404.4]
  assign _T_39641 = io_inAddr_14 == 6'h39; // @[Switch.scala 30:53:@18406.4]
  assign valid_57_14 = io_inValid_14 & _T_39641; // @[Switch.scala 30:36:@18407.4]
  assign _T_39644 = io_inAddr_15 == 6'h39; // @[Switch.scala 30:53:@18409.4]
  assign valid_57_15 = io_inValid_15 & _T_39644; // @[Switch.scala 30:36:@18410.4]
  assign _T_39647 = io_inAddr_16 == 6'h39; // @[Switch.scala 30:53:@18412.4]
  assign valid_57_16 = io_inValid_16 & _T_39647; // @[Switch.scala 30:36:@18413.4]
  assign _T_39650 = io_inAddr_17 == 6'h39; // @[Switch.scala 30:53:@18415.4]
  assign valid_57_17 = io_inValid_17 & _T_39650; // @[Switch.scala 30:36:@18416.4]
  assign _T_39653 = io_inAddr_18 == 6'h39; // @[Switch.scala 30:53:@18418.4]
  assign valid_57_18 = io_inValid_18 & _T_39653; // @[Switch.scala 30:36:@18419.4]
  assign _T_39656 = io_inAddr_19 == 6'h39; // @[Switch.scala 30:53:@18421.4]
  assign valid_57_19 = io_inValid_19 & _T_39656; // @[Switch.scala 30:36:@18422.4]
  assign _T_39659 = io_inAddr_20 == 6'h39; // @[Switch.scala 30:53:@18424.4]
  assign valid_57_20 = io_inValid_20 & _T_39659; // @[Switch.scala 30:36:@18425.4]
  assign _T_39662 = io_inAddr_21 == 6'h39; // @[Switch.scala 30:53:@18427.4]
  assign valid_57_21 = io_inValid_21 & _T_39662; // @[Switch.scala 30:36:@18428.4]
  assign _T_39665 = io_inAddr_22 == 6'h39; // @[Switch.scala 30:53:@18430.4]
  assign valid_57_22 = io_inValid_22 & _T_39665; // @[Switch.scala 30:36:@18431.4]
  assign _T_39668 = io_inAddr_23 == 6'h39; // @[Switch.scala 30:53:@18433.4]
  assign valid_57_23 = io_inValid_23 & _T_39668; // @[Switch.scala 30:36:@18434.4]
  assign _T_39671 = io_inAddr_24 == 6'h39; // @[Switch.scala 30:53:@18436.4]
  assign valid_57_24 = io_inValid_24 & _T_39671; // @[Switch.scala 30:36:@18437.4]
  assign _T_39674 = io_inAddr_25 == 6'h39; // @[Switch.scala 30:53:@18439.4]
  assign valid_57_25 = io_inValid_25 & _T_39674; // @[Switch.scala 30:36:@18440.4]
  assign _T_39677 = io_inAddr_26 == 6'h39; // @[Switch.scala 30:53:@18442.4]
  assign valid_57_26 = io_inValid_26 & _T_39677; // @[Switch.scala 30:36:@18443.4]
  assign _T_39680 = io_inAddr_27 == 6'h39; // @[Switch.scala 30:53:@18445.4]
  assign valid_57_27 = io_inValid_27 & _T_39680; // @[Switch.scala 30:36:@18446.4]
  assign _T_39683 = io_inAddr_28 == 6'h39; // @[Switch.scala 30:53:@18448.4]
  assign valid_57_28 = io_inValid_28 & _T_39683; // @[Switch.scala 30:36:@18449.4]
  assign _T_39686 = io_inAddr_29 == 6'h39; // @[Switch.scala 30:53:@18451.4]
  assign valid_57_29 = io_inValid_29 & _T_39686; // @[Switch.scala 30:36:@18452.4]
  assign _T_39689 = io_inAddr_30 == 6'h39; // @[Switch.scala 30:53:@18454.4]
  assign valid_57_30 = io_inValid_30 & _T_39689; // @[Switch.scala 30:36:@18455.4]
  assign _T_39692 = io_inAddr_31 == 6'h39; // @[Switch.scala 30:53:@18457.4]
  assign valid_57_31 = io_inValid_31 & _T_39692; // @[Switch.scala 30:36:@18458.4]
  assign _T_39695 = io_inAddr_32 == 6'h39; // @[Switch.scala 30:53:@18460.4]
  assign valid_57_32 = io_inValid_32 & _T_39695; // @[Switch.scala 30:36:@18461.4]
  assign _T_39698 = io_inAddr_33 == 6'h39; // @[Switch.scala 30:53:@18463.4]
  assign valid_57_33 = io_inValid_33 & _T_39698; // @[Switch.scala 30:36:@18464.4]
  assign _T_39701 = io_inAddr_34 == 6'h39; // @[Switch.scala 30:53:@18466.4]
  assign valid_57_34 = io_inValid_34 & _T_39701; // @[Switch.scala 30:36:@18467.4]
  assign _T_39704 = io_inAddr_35 == 6'h39; // @[Switch.scala 30:53:@18469.4]
  assign valid_57_35 = io_inValid_35 & _T_39704; // @[Switch.scala 30:36:@18470.4]
  assign _T_39707 = io_inAddr_36 == 6'h39; // @[Switch.scala 30:53:@18472.4]
  assign valid_57_36 = io_inValid_36 & _T_39707; // @[Switch.scala 30:36:@18473.4]
  assign _T_39710 = io_inAddr_37 == 6'h39; // @[Switch.scala 30:53:@18475.4]
  assign valid_57_37 = io_inValid_37 & _T_39710; // @[Switch.scala 30:36:@18476.4]
  assign _T_39713 = io_inAddr_38 == 6'h39; // @[Switch.scala 30:53:@18478.4]
  assign valid_57_38 = io_inValid_38 & _T_39713; // @[Switch.scala 30:36:@18479.4]
  assign _T_39716 = io_inAddr_39 == 6'h39; // @[Switch.scala 30:53:@18481.4]
  assign valid_57_39 = io_inValid_39 & _T_39716; // @[Switch.scala 30:36:@18482.4]
  assign _T_39719 = io_inAddr_40 == 6'h39; // @[Switch.scala 30:53:@18484.4]
  assign valid_57_40 = io_inValid_40 & _T_39719; // @[Switch.scala 30:36:@18485.4]
  assign _T_39722 = io_inAddr_41 == 6'h39; // @[Switch.scala 30:53:@18487.4]
  assign valid_57_41 = io_inValid_41 & _T_39722; // @[Switch.scala 30:36:@18488.4]
  assign _T_39725 = io_inAddr_42 == 6'h39; // @[Switch.scala 30:53:@18490.4]
  assign valid_57_42 = io_inValid_42 & _T_39725; // @[Switch.scala 30:36:@18491.4]
  assign _T_39728 = io_inAddr_43 == 6'h39; // @[Switch.scala 30:53:@18493.4]
  assign valid_57_43 = io_inValid_43 & _T_39728; // @[Switch.scala 30:36:@18494.4]
  assign _T_39731 = io_inAddr_44 == 6'h39; // @[Switch.scala 30:53:@18496.4]
  assign valid_57_44 = io_inValid_44 & _T_39731; // @[Switch.scala 30:36:@18497.4]
  assign _T_39734 = io_inAddr_45 == 6'h39; // @[Switch.scala 30:53:@18499.4]
  assign valid_57_45 = io_inValid_45 & _T_39734; // @[Switch.scala 30:36:@18500.4]
  assign _T_39737 = io_inAddr_46 == 6'h39; // @[Switch.scala 30:53:@18502.4]
  assign valid_57_46 = io_inValid_46 & _T_39737; // @[Switch.scala 30:36:@18503.4]
  assign _T_39740 = io_inAddr_47 == 6'h39; // @[Switch.scala 30:53:@18505.4]
  assign valid_57_47 = io_inValid_47 & _T_39740; // @[Switch.scala 30:36:@18506.4]
  assign _T_39743 = io_inAddr_48 == 6'h39; // @[Switch.scala 30:53:@18508.4]
  assign valid_57_48 = io_inValid_48 & _T_39743; // @[Switch.scala 30:36:@18509.4]
  assign _T_39746 = io_inAddr_49 == 6'h39; // @[Switch.scala 30:53:@18511.4]
  assign valid_57_49 = io_inValid_49 & _T_39746; // @[Switch.scala 30:36:@18512.4]
  assign _T_39749 = io_inAddr_50 == 6'h39; // @[Switch.scala 30:53:@18514.4]
  assign valid_57_50 = io_inValid_50 & _T_39749; // @[Switch.scala 30:36:@18515.4]
  assign _T_39752 = io_inAddr_51 == 6'h39; // @[Switch.scala 30:53:@18517.4]
  assign valid_57_51 = io_inValid_51 & _T_39752; // @[Switch.scala 30:36:@18518.4]
  assign _T_39755 = io_inAddr_52 == 6'h39; // @[Switch.scala 30:53:@18520.4]
  assign valid_57_52 = io_inValid_52 & _T_39755; // @[Switch.scala 30:36:@18521.4]
  assign _T_39758 = io_inAddr_53 == 6'h39; // @[Switch.scala 30:53:@18523.4]
  assign valid_57_53 = io_inValid_53 & _T_39758; // @[Switch.scala 30:36:@18524.4]
  assign _T_39761 = io_inAddr_54 == 6'h39; // @[Switch.scala 30:53:@18526.4]
  assign valid_57_54 = io_inValid_54 & _T_39761; // @[Switch.scala 30:36:@18527.4]
  assign _T_39764 = io_inAddr_55 == 6'h39; // @[Switch.scala 30:53:@18529.4]
  assign valid_57_55 = io_inValid_55 & _T_39764; // @[Switch.scala 30:36:@18530.4]
  assign _T_39767 = io_inAddr_56 == 6'h39; // @[Switch.scala 30:53:@18532.4]
  assign valid_57_56 = io_inValid_56 & _T_39767; // @[Switch.scala 30:36:@18533.4]
  assign _T_39770 = io_inAddr_57 == 6'h39; // @[Switch.scala 30:53:@18535.4]
  assign valid_57_57 = io_inValid_57 & _T_39770; // @[Switch.scala 30:36:@18536.4]
  assign _T_39773 = io_inAddr_58 == 6'h39; // @[Switch.scala 30:53:@18538.4]
  assign valid_57_58 = io_inValid_58 & _T_39773; // @[Switch.scala 30:36:@18539.4]
  assign _T_39776 = io_inAddr_59 == 6'h39; // @[Switch.scala 30:53:@18541.4]
  assign valid_57_59 = io_inValid_59 & _T_39776; // @[Switch.scala 30:36:@18542.4]
  assign _T_39779 = io_inAddr_60 == 6'h39; // @[Switch.scala 30:53:@18544.4]
  assign valid_57_60 = io_inValid_60 & _T_39779; // @[Switch.scala 30:36:@18545.4]
  assign _T_39782 = io_inAddr_61 == 6'h39; // @[Switch.scala 30:53:@18547.4]
  assign valid_57_61 = io_inValid_61 & _T_39782; // @[Switch.scala 30:36:@18548.4]
  assign _T_39785 = io_inAddr_62 == 6'h39; // @[Switch.scala 30:53:@18550.4]
  assign valid_57_62 = io_inValid_62 & _T_39785; // @[Switch.scala 30:36:@18551.4]
  assign _T_39788 = io_inAddr_63 == 6'h39; // @[Switch.scala 30:53:@18553.4]
  assign valid_57_63 = io_inValid_63 & _T_39788; // @[Switch.scala 30:36:@18554.4]
  assign _T_39854 = valid_57_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@18556.4]
  assign _T_39855 = valid_57_61 ? 6'h3d : _T_39854; // @[Mux.scala 31:69:@18557.4]
  assign _T_39856 = valid_57_60 ? 6'h3c : _T_39855; // @[Mux.scala 31:69:@18558.4]
  assign _T_39857 = valid_57_59 ? 6'h3b : _T_39856; // @[Mux.scala 31:69:@18559.4]
  assign _T_39858 = valid_57_58 ? 6'h3a : _T_39857; // @[Mux.scala 31:69:@18560.4]
  assign _T_39859 = valid_57_57 ? 6'h39 : _T_39858; // @[Mux.scala 31:69:@18561.4]
  assign _T_39860 = valid_57_56 ? 6'h38 : _T_39859; // @[Mux.scala 31:69:@18562.4]
  assign _T_39861 = valid_57_55 ? 6'h37 : _T_39860; // @[Mux.scala 31:69:@18563.4]
  assign _T_39862 = valid_57_54 ? 6'h36 : _T_39861; // @[Mux.scala 31:69:@18564.4]
  assign _T_39863 = valid_57_53 ? 6'h35 : _T_39862; // @[Mux.scala 31:69:@18565.4]
  assign _T_39864 = valid_57_52 ? 6'h34 : _T_39863; // @[Mux.scala 31:69:@18566.4]
  assign _T_39865 = valid_57_51 ? 6'h33 : _T_39864; // @[Mux.scala 31:69:@18567.4]
  assign _T_39866 = valid_57_50 ? 6'h32 : _T_39865; // @[Mux.scala 31:69:@18568.4]
  assign _T_39867 = valid_57_49 ? 6'h31 : _T_39866; // @[Mux.scala 31:69:@18569.4]
  assign _T_39868 = valid_57_48 ? 6'h30 : _T_39867; // @[Mux.scala 31:69:@18570.4]
  assign _T_39869 = valid_57_47 ? 6'h2f : _T_39868; // @[Mux.scala 31:69:@18571.4]
  assign _T_39870 = valid_57_46 ? 6'h2e : _T_39869; // @[Mux.scala 31:69:@18572.4]
  assign _T_39871 = valid_57_45 ? 6'h2d : _T_39870; // @[Mux.scala 31:69:@18573.4]
  assign _T_39872 = valid_57_44 ? 6'h2c : _T_39871; // @[Mux.scala 31:69:@18574.4]
  assign _T_39873 = valid_57_43 ? 6'h2b : _T_39872; // @[Mux.scala 31:69:@18575.4]
  assign _T_39874 = valid_57_42 ? 6'h2a : _T_39873; // @[Mux.scala 31:69:@18576.4]
  assign _T_39875 = valid_57_41 ? 6'h29 : _T_39874; // @[Mux.scala 31:69:@18577.4]
  assign _T_39876 = valid_57_40 ? 6'h28 : _T_39875; // @[Mux.scala 31:69:@18578.4]
  assign _T_39877 = valid_57_39 ? 6'h27 : _T_39876; // @[Mux.scala 31:69:@18579.4]
  assign _T_39878 = valid_57_38 ? 6'h26 : _T_39877; // @[Mux.scala 31:69:@18580.4]
  assign _T_39879 = valid_57_37 ? 6'h25 : _T_39878; // @[Mux.scala 31:69:@18581.4]
  assign _T_39880 = valid_57_36 ? 6'h24 : _T_39879; // @[Mux.scala 31:69:@18582.4]
  assign _T_39881 = valid_57_35 ? 6'h23 : _T_39880; // @[Mux.scala 31:69:@18583.4]
  assign _T_39882 = valid_57_34 ? 6'h22 : _T_39881; // @[Mux.scala 31:69:@18584.4]
  assign _T_39883 = valid_57_33 ? 6'h21 : _T_39882; // @[Mux.scala 31:69:@18585.4]
  assign _T_39884 = valid_57_32 ? 6'h20 : _T_39883; // @[Mux.scala 31:69:@18586.4]
  assign _T_39885 = valid_57_31 ? 6'h1f : _T_39884; // @[Mux.scala 31:69:@18587.4]
  assign _T_39886 = valid_57_30 ? 6'h1e : _T_39885; // @[Mux.scala 31:69:@18588.4]
  assign _T_39887 = valid_57_29 ? 6'h1d : _T_39886; // @[Mux.scala 31:69:@18589.4]
  assign _T_39888 = valid_57_28 ? 6'h1c : _T_39887; // @[Mux.scala 31:69:@18590.4]
  assign _T_39889 = valid_57_27 ? 6'h1b : _T_39888; // @[Mux.scala 31:69:@18591.4]
  assign _T_39890 = valid_57_26 ? 6'h1a : _T_39889; // @[Mux.scala 31:69:@18592.4]
  assign _T_39891 = valid_57_25 ? 6'h19 : _T_39890; // @[Mux.scala 31:69:@18593.4]
  assign _T_39892 = valid_57_24 ? 6'h18 : _T_39891; // @[Mux.scala 31:69:@18594.4]
  assign _T_39893 = valid_57_23 ? 6'h17 : _T_39892; // @[Mux.scala 31:69:@18595.4]
  assign _T_39894 = valid_57_22 ? 6'h16 : _T_39893; // @[Mux.scala 31:69:@18596.4]
  assign _T_39895 = valid_57_21 ? 6'h15 : _T_39894; // @[Mux.scala 31:69:@18597.4]
  assign _T_39896 = valid_57_20 ? 6'h14 : _T_39895; // @[Mux.scala 31:69:@18598.4]
  assign _T_39897 = valid_57_19 ? 6'h13 : _T_39896; // @[Mux.scala 31:69:@18599.4]
  assign _T_39898 = valid_57_18 ? 6'h12 : _T_39897; // @[Mux.scala 31:69:@18600.4]
  assign _T_39899 = valid_57_17 ? 6'h11 : _T_39898; // @[Mux.scala 31:69:@18601.4]
  assign _T_39900 = valid_57_16 ? 6'h10 : _T_39899; // @[Mux.scala 31:69:@18602.4]
  assign _T_39901 = valid_57_15 ? 6'hf : _T_39900; // @[Mux.scala 31:69:@18603.4]
  assign _T_39902 = valid_57_14 ? 6'he : _T_39901; // @[Mux.scala 31:69:@18604.4]
  assign _T_39903 = valid_57_13 ? 6'hd : _T_39902; // @[Mux.scala 31:69:@18605.4]
  assign _T_39904 = valid_57_12 ? 6'hc : _T_39903; // @[Mux.scala 31:69:@18606.4]
  assign _T_39905 = valid_57_11 ? 6'hb : _T_39904; // @[Mux.scala 31:69:@18607.4]
  assign _T_39906 = valid_57_10 ? 6'ha : _T_39905; // @[Mux.scala 31:69:@18608.4]
  assign _T_39907 = valid_57_9 ? 6'h9 : _T_39906; // @[Mux.scala 31:69:@18609.4]
  assign _T_39908 = valid_57_8 ? 6'h8 : _T_39907; // @[Mux.scala 31:69:@18610.4]
  assign _T_39909 = valid_57_7 ? 6'h7 : _T_39908; // @[Mux.scala 31:69:@18611.4]
  assign _T_39910 = valid_57_6 ? 6'h6 : _T_39909; // @[Mux.scala 31:69:@18612.4]
  assign _T_39911 = valid_57_5 ? 6'h5 : _T_39910; // @[Mux.scala 31:69:@18613.4]
  assign _T_39912 = valid_57_4 ? 6'h4 : _T_39911; // @[Mux.scala 31:69:@18614.4]
  assign _T_39913 = valid_57_3 ? 6'h3 : _T_39912; // @[Mux.scala 31:69:@18615.4]
  assign _T_39914 = valid_57_2 ? 6'h2 : _T_39913; // @[Mux.scala 31:69:@18616.4]
  assign _T_39915 = valid_57_1 ? 6'h1 : _T_39914; // @[Mux.scala 31:69:@18617.4]
  assign select_57 = valid_57_0 ? 6'h0 : _T_39915; // @[Mux.scala 31:69:@18618.4]
  assign _GEN_3649 = 6'h1 == select_57 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3650 = 6'h2 == select_57 ? io_inData_2 : _GEN_3649; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3651 = 6'h3 == select_57 ? io_inData_3 : _GEN_3650; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3652 = 6'h4 == select_57 ? io_inData_4 : _GEN_3651; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3653 = 6'h5 == select_57 ? io_inData_5 : _GEN_3652; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3654 = 6'h6 == select_57 ? io_inData_6 : _GEN_3653; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3655 = 6'h7 == select_57 ? io_inData_7 : _GEN_3654; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3656 = 6'h8 == select_57 ? io_inData_8 : _GEN_3655; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3657 = 6'h9 == select_57 ? io_inData_9 : _GEN_3656; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3658 = 6'ha == select_57 ? io_inData_10 : _GEN_3657; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3659 = 6'hb == select_57 ? io_inData_11 : _GEN_3658; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3660 = 6'hc == select_57 ? io_inData_12 : _GEN_3659; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3661 = 6'hd == select_57 ? io_inData_13 : _GEN_3660; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3662 = 6'he == select_57 ? io_inData_14 : _GEN_3661; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3663 = 6'hf == select_57 ? io_inData_15 : _GEN_3662; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3664 = 6'h10 == select_57 ? io_inData_16 : _GEN_3663; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3665 = 6'h11 == select_57 ? io_inData_17 : _GEN_3664; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3666 = 6'h12 == select_57 ? io_inData_18 : _GEN_3665; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3667 = 6'h13 == select_57 ? io_inData_19 : _GEN_3666; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3668 = 6'h14 == select_57 ? io_inData_20 : _GEN_3667; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3669 = 6'h15 == select_57 ? io_inData_21 : _GEN_3668; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3670 = 6'h16 == select_57 ? io_inData_22 : _GEN_3669; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3671 = 6'h17 == select_57 ? io_inData_23 : _GEN_3670; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3672 = 6'h18 == select_57 ? io_inData_24 : _GEN_3671; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3673 = 6'h19 == select_57 ? io_inData_25 : _GEN_3672; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3674 = 6'h1a == select_57 ? io_inData_26 : _GEN_3673; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3675 = 6'h1b == select_57 ? io_inData_27 : _GEN_3674; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3676 = 6'h1c == select_57 ? io_inData_28 : _GEN_3675; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3677 = 6'h1d == select_57 ? io_inData_29 : _GEN_3676; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3678 = 6'h1e == select_57 ? io_inData_30 : _GEN_3677; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3679 = 6'h1f == select_57 ? io_inData_31 : _GEN_3678; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3680 = 6'h20 == select_57 ? io_inData_32 : _GEN_3679; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3681 = 6'h21 == select_57 ? io_inData_33 : _GEN_3680; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3682 = 6'h22 == select_57 ? io_inData_34 : _GEN_3681; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3683 = 6'h23 == select_57 ? io_inData_35 : _GEN_3682; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3684 = 6'h24 == select_57 ? io_inData_36 : _GEN_3683; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3685 = 6'h25 == select_57 ? io_inData_37 : _GEN_3684; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3686 = 6'h26 == select_57 ? io_inData_38 : _GEN_3685; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3687 = 6'h27 == select_57 ? io_inData_39 : _GEN_3686; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3688 = 6'h28 == select_57 ? io_inData_40 : _GEN_3687; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3689 = 6'h29 == select_57 ? io_inData_41 : _GEN_3688; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3690 = 6'h2a == select_57 ? io_inData_42 : _GEN_3689; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3691 = 6'h2b == select_57 ? io_inData_43 : _GEN_3690; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3692 = 6'h2c == select_57 ? io_inData_44 : _GEN_3691; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3693 = 6'h2d == select_57 ? io_inData_45 : _GEN_3692; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3694 = 6'h2e == select_57 ? io_inData_46 : _GEN_3693; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3695 = 6'h2f == select_57 ? io_inData_47 : _GEN_3694; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3696 = 6'h30 == select_57 ? io_inData_48 : _GEN_3695; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3697 = 6'h31 == select_57 ? io_inData_49 : _GEN_3696; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3698 = 6'h32 == select_57 ? io_inData_50 : _GEN_3697; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3699 = 6'h33 == select_57 ? io_inData_51 : _GEN_3698; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3700 = 6'h34 == select_57 ? io_inData_52 : _GEN_3699; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3701 = 6'h35 == select_57 ? io_inData_53 : _GEN_3700; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3702 = 6'h36 == select_57 ? io_inData_54 : _GEN_3701; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3703 = 6'h37 == select_57 ? io_inData_55 : _GEN_3702; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3704 = 6'h38 == select_57 ? io_inData_56 : _GEN_3703; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3705 = 6'h39 == select_57 ? io_inData_57 : _GEN_3704; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3706 = 6'h3a == select_57 ? io_inData_58 : _GEN_3705; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3707 = 6'h3b == select_57 ? io_inData_59 : _GEN_3706; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3708 = 6'h3c == select_57 ? io_inData_60 : _GEN_3707; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3709 = 6'h3d == select_57 ? io_inData_61 : _GEN_3708; // @[Switch.scala 33:19:@18620.4]
  assign _GEN_3710 = 6'h3e == select_57 ? io_inData_62 : _GEN_3709; // @[Switch.scala 33:19:@18620.4]
  assign _T_39924 = {valid_57_7,valid_57_6,valid_57_5,valid_57_4,valid_57_3,valid_57_2,valid_57_1,valid_57_0}; // @[Switch.scala 34:32:@18627.4]
  assign _T_39932 = {valid_57_15,valid_57_14,valid_57_13,valid_57_12,valid_57_11,valid_57_10,valid_57_9,valid_57_8,_T_39924}; // @[Switch.scala 34:32:@18635.4]
  assign _T_39939 = {valid_57_23,valid_57_22,valid_57_21,valid_57_20,valid_57_19,valid_57_18,valid_57_17,valid_57_16}; // @[Switch.scala 34:32:@18642.4]
  assign _T_39948 = {valid_57_31,valid_57_30,valid_57_29,valid_57_28,valid_57_27,valid_57_26,valid_57_25,valid_57_24,_T_39939,_T_39932}; // @[Switch.scala 34:32:@18651.4]
  assign _T_39955 = {valid_57_39,valid_57_38,valid_57_37,valid_57_36,valid_57_35,valid_57_34,valid_57_33,valid_57_32}; // @[Switch.scala 34:32:@18658.4]
  assign _T_39963 = {valid_57_47,valid_57_46,valid_57_45,valid_57_44,valid_57_43,valid_57_42,valid_57_41,valid_57_40,_T_39955}; // @[Switch.scala 34:32:@18666.4]
  assign _T_39970 = {valid_57_55,valid_57_54,valid_57_53,valid_57_52,valid_57_51,valid_57_50,valid_57_49,valid_57_48}; // @[Switch.scala 34:32:@18673.4]
  assign _T_39979 = {valid_57_63,valid_57_62,valid_57_61,valid_57_60,valid_57_59,valid_57_58,valid_57_57,valid_57_56,_T_39970,_T_39963}; // @[Switch.scala 34:32:@18682.4]
  assign _T_39980 = {_T_39979,_T_39948}; // @[Switch.scala 34:32:@18683.4]
  assign _T_39984 = io_inAddr_0 == 6'h3a; // @[Switch.scala 30:53:@18686.4]
  assign valid_58_0 = io_inValid_0 & _T_39984; // @[Switch.scala 30:36:@18687.4]
  assign _T_39987 = io_inAddr_1 == 6'h3a; // @[Switch.scala 30:53:@18689.4]
  assign valid_58_1 = io_inValid_1 & _T_39987; // @[Switch.scala 30:36:@18690.4]
  assign _T_39990 = io_inAddr_2 == 6'h3a; // @[Switch.scala 30:53:@18692.4]
  assign valid_58_2 = io_inValid_2 & _T_39990; // @[Switch.scala 30:36:@18693.4]
  assign _T_39993 = io_inAddr_3 == 6'h3a; // @[Switch.scala 30:53:@18695.4]
  assign valid_58_3 = io_inValid_3 & _T_39993; // @[Switch.scala 30:36:@18696.4]
  assign _T_39996 = io_inAddr_4 == 6'h3a; // @[Switch.scala 30:53:@18698.4]
  assign valid_58_4 = io_inValid_4 & _T_39996; // @[Switch.scala 30:36:@18699.4]
  assign _T_39999 = io_inAddr_5 == 6'h3a; // @[Switch.scala 30:53:@18701.4]
  assign valid_58_5 = io_inValid_5 & _T_39999; // @[Switch.scala 30:36:@18702.4]
  assign _T_40002 = io_inAddr_6 == 6'h3a; // @[Switch.scala 30:53:@18704.4]
  assign valid_58_6 = io_inValid_6 & _T_40002; // @[Switch.scala 30:36:@18705.4]
  assign _T_40005 = io_inAddr_7 == 6'h3a; // @[Switch.scala 30:53:@18707.4]
  assign valid_58_7 = io_inValid_7 & _T_40005; // @[Switch.scala 30:36:@18708.4]
  assign _T_40008 = io_inAddr_8 == 6'h3a; // @[Switch.scala 30:53:@18710.4]
  assign valid_58_8 = io_inValid_8 & _T_40008; // @[Switch.scala 30:36:@18711.4]
  assign _T_40011 = io_inAddr_9 == 6'h3a; // @[Switch.scala 30:53:@18713.4]
  assign valid_58_9 = io_inValid_9 & _T_40011; // @[Switch.scala 30:36:@18714.4]
  assign _T_40014 = io_inAddr_10 == 6'h3a; // @[Switch.scala 30:53:@18716.4]
  assign valid_58_10 = io_inValid_10 & _T_40014; // @[Switch.scala 30:36:@18717.4]
  assign _T_40017 = io_inAddr_11 == 6'h3a; // @[Switch.scala 30:53:@18719.4]
  assign valid_58_11 = io_inValid_11 & _T_40017; // @[Switch.scala 30:36:@18720.4]
  assign _T_40020 = io_inAddr_12 == 6'h3a; // @[Switch.scala 30:53:@18722.4]
  assign valid_58_12 = io_inValid_12 & _T_40020; // @[Switch.scala 30:36:@18723.4]
  assign _T_40023 = io_inAddr_13 == 6'h3a; // @[Switch.scala 30:53:@18725.4]
  assign valid_58_13 = io_inValid_13 & _T_40023; // @[Switch.scala 30:36:@18726.4]
  assign _T_40026 = io_inAddr_14 == 6'h3a; // @[Switch.scala 30:53:@18728.4]
  assign valid_58_14 = io_inValid_14 & _T_40026; // @[Switch.scala 30:36:@18729.4]
  assign _T_40029 = io_inAddr_15 == 6'h3a; // @[Switch.scala 30:53:@18731.4]
  assign valid_58_15 = io_inValid_15 & _T_40029; // @[Switch.scala 30:36:@18732.4]
  assign _T_40032 = io_inAddr_16 == 6'h3a; // @[Switch.scala 30:53:@18734.4]
  assign valid_58_16 = io_inValid_16 & _T_40032; // @[Switch.scala 30:36:@18735.4]
  assign _T_40035 = io_inAddr_17 == 6'h3a; // @[Switch.scala 30:53:@18737.4]
  assign valid_58_17 = io_inValid_17 & _T_40035; // @[Switch.scala 30:36:@18738.4]
  assign _T_40038 = io_inAddr_18 == 6'h3a; // @[Switch.scala 30:53:@18740.4]
  assign valid_58_18 = io_inValid_18 & _T_40038; // @[Switch.scala 30:36:@18741.4]
  assign _T_40041 = io_inAddr_19 == 6'h3a; // @[Switch.scala 30:53:@18743.4]
  assign valid_58_19 = io_inValid_19 & _T_40041; // @[Switch.scala 30:36:@18744.4]
  assign _T_40044 = io_inAddr_20 == 6'h3a; // @[Switch.scala 30:53:@18746.4]
  assign valid_58_20 = io_inValid_20 & _T_40044; // @[Switch.scala 30:36:@18747.4]
  assign _T_40047 = io_inAddr_21 == 6'h3a; // @[Switch.scala 30:53:@18749.4]
  assign valid_58_21 = io_inValid_21 & _T_40047; // @[Switch.scala 30:36:@18750.4]
  assign _T_40050 = io_inAddr_22 == 6'h3a; // @[Switch.scala 30:53:@18752.4]
  assign valid_58_22 = io_inValid_22 & _T_40050; // @[Switch.scala 30:36:@18753.4]
  assign _T_40053 = io_inAddr_23 == 6'h3a; // @[Switch.scala 30:53:@18755.4]
  assign valid_58_23 = io_inValid_23 & _T_40053; // @[Switch.scala 30:36:@18756.4]
  assign _T_40056 = io_inAddr_24 == 6'h3a; // @[Switch.scala 30:53:@18758.4]
  assign valid_58_24 = io_inValid_24 & _T_40056; // @[Switch.scala 30:36:@18759.4]
  assign _T_40059 = io_inAddr_25 == 6'h3a; // @[Switch.scala 30:53:@18761.4]
  assign valid_58_25 = io_inValid_25 & _T_40059; // @[Switch.scala 30:36:@18762.4]
  assign _T_40062 = io_inAddr_26 == 6'h3a; // @[Switch.scala 30:53:@18764.4]
  assign valid_58_26 = io_inValid_26 & _T_40062; // @[Switch.scala 30:36:@18765.4]
  assign _T_40065 = io_inAddr_27 == 6'h3a; // @[Switch.scala 30:53:@18767.4]
  assign valid_58_27 = io_inValid_27 & _T_40065; // @[Switch.scala 30:36:@18768.4]
  assign _T_40068 = io_inAddr_28 == 6'h3a; // @[Switch.scala 30:53:@18770.4]
  assign valid_58_28 = io_inValid_28 & _T_40068; // @[Switch.scala 30:36:@18771.4]
  assign _T_40071 = io_inAddr_29 == 6'h3a; // @[Switch.scala 30:53:@18773.4]
  assign valid_58_29 = io_inValid_29 & _T_40071; // @[Switch.scala 30:36:@18774.4]
  assign _T_40074 = io_inAddr_30 == 6'h3a; // @[Switch.scala 30:53:@18776.4]
  assign valid_58_30 = io_inValid_30 & _T_40074; // @[Switch.scala 30:36:@18777.4]
  assign _T_40077 = io_inAddr_31 == 6'h3a; // @[Switch.scala 30:53:@18779.4]
  assign valid_58_31 = io_inValid_31 & _T_40077; // @[Switch.scala 30:36:@18780.4]
  assign _T_40080 = io_inAddr_32 == 6'h3a; // @[Switch.scala 30:53:@18782.4]
  assign valid_58_32 = io_inValid_32 & _T_40080; // @[Switch.scala 30:36:@18783.4]
  assign _T_40083 = io_inAddr_33 == 6'h3a; // @[Switch.scala 30:53:@18785.4]
  assign valid_58_33 = io_inValid_33 & _T_40083; // @[Switch.scala 30:36:@18786.4]
  assign _T_40086 = io_inAddr_34 == 6'h3a; // @[Switch.scala 30:53:@18788.4]
  assign valid_58_34 = io_inValid_34 & _T_40086; // @[Switch.scala 30:36:@18789.4]
  assign _T_40089 = io_inAddr_35 == 6'h3a; // @[Switch.scala 30:53:@18791.4]
  assign valid_58_35 = io_inValid_35 & _T_40089; // @[Switch.scala 30:36:@18792.4]
  assign _T_40092 = io_inAddr_36 == 6'h3a; // @[Switch.scala 30:53:@18794.4]
  assign valid_58_36 = io_inValid_36 & _T_40092; // @[Switch.scala 30:36:@18795.4]
  assign _T_40095 = io_inAddr_37 == 6'h3a; // @[Switch.scala 30:53:@18797.4]
  assign valid_58_37 = io_inValid_37 & _T_40095; // @[Switch.scala 30:36:@18798.4]
  assign _T_40098 = io_inAddr_38 == 6'h3a; // @[Switch.scala 30:53:@18800.4]
  assign valid_58_38 = io_inValid_38 & _T_40098; // @[Switch.scala 30:36:@18801.4]
  assign _T_40101 = io_inAddr_39 == 6'h3a; // @[Switch.scala 30:53:@18803.4]
  assign valid_58_39 = io_inValid_39 & _T_40101; // @[Switch.scala 30:36:@18804.4]
  assign _T_40104 = io_inAddr_40 == 6'h3a; // @[Switch.scala 30:53:@18806.4]
  assign valid_58_40 = io_inValid_40 & _T_40104; // @[Switch.scala 30:36:@18807.4]
  assign _T_40107 = io_inAddr_41 == 6'h3a; // @[Switch.scala 30:53:@18809.4]
  assign valid_58_41 = io_inValid_41 & _T_40107; // @[Switch.scala 30:36:@18810.4]
  assign _T_40110 = io_inAddr_42 == 6'h3a; // @[Switch.scala 30:53:@18812.4]
  assign valid_58_42 = io_inValid_42 & _T_40110; // @[Switch.scala 30:36:@18813.4]
  assign _T_40113 = io_inAddr_43 == 6'h3a; // @[Switch.scala 30:53:@18815.4]
  assign valid_58_43 = io_inValid_43 & _T_40113; // @[Switch.scala 30:36:@18816.4]
  assign _T_40116 = io_inAddr_44 == 6'h3a; // @[Switch.scala 30:53:@18818.4]
  assign valid_58_44 = io_inValid_44 & _T_40116; // @[Switch.scala 30:36:@18819.4]
  assign _T_40119 = io_inAddr_45 == 6'h3a; // @[Switch.scala 30:53:@18821.4]
  assign valid_58_45 = io_inValid_45 & _T_40119; // @[Switch.scala 30:36:@18822.4]
  assign _T_40122 = io_inAddr_46 == 6'h3a; // @[Switch.scala 30:53:@18824.4]
  assign valid_58_46 = io_inValid_46 & _T_40122; // @[Switch.scala 30:36:@18825.4]
  assign _T_40125 = io_inAddr_47 == 6'h3a; // @[Switch.scala 30:53:@18827.4]
  assign valid_58_47 = io_inValid_47 & _T_40125; // @[Switch.scala 30:36:@18828.4]
  assign _T_40128 = io_inAddr_48 == 6'h3a; // @[Switch.scala 30:53:@18830.4]
  assign valid_58_48 = io_inValid_48 & _T_40128; // @[Switch.scala 30:36:@18831.4]
  assign _T_40131 = io_inAddr_49 == 6'h3a; // @[Switch.scala 30:53:@18833.4]
  assign valid_58_49 = io_inValid_49 & _T_40131; // @[Switch.scala 30:36:@18834.4]
  assign _T_40134 = io_inAddr_50 == 6'h3a; // @[Switch.scala 30:53:@18836.4]
  assign valid_58_50 = io_inValid_50 & _T_40134; // @[Switch.scala 30:36:@18837.4]
  assign _T_40137 = io_inAddr_51 == 6'h3a; // @[Switch.scala 30:53:@18839.4]
  assign valid_58_51 = io_inValid_51 & _T_40137; // @[Switch.scala 30:36:@18840.4]
  assign _T_40140 = io_inAddr_52 == 6'h3a; // @[Switch.scala 30:53:@18842.4]
  assign valid_58_52 = io_inValid_52 & _T_40140; // @[Switch.scala 30:36:@18843.4]
  assign _T_40143 = io_inAddr_53 == 6'h3a; // @[Switch.scala 30:53:@18845.4]
  assign valid_58_53 = io_inValid_53 & _T_40143; // @[Switch.scala 30:36:@18846.4]
  assign _T_40146 = io_inAddr_54 == 6'h3a; // @[Switch.scala 30:53:@18848.4]
  assign valid_58_54 = io_inValid_54 & _T_40146; // @[Switch.scala 30:36:@18849.4]
  assign _T_40149 = io_inAddr_55 == 6'h3a; // @[Switch.scala 30:53:@18851.4]
  assign valid_58_55 = io_inValid_55 & _T_40149; // @[Switch.scala 30:36:@18852.4]
  assign _T_40152 = io_inAddr_56 == 6'h3a; // @[Switch.scala 30:53:@18854.4]
  assign valid_58_56 = io_inValid_56 & _T_40152; // @[Switch.scala 30:36:@18855.4]
  assign _T_40155 = io_inAddr_57 == 6'h3a; // @[Switch.scala 30:53:@18857.4]
  assign valid_58_57 = io_inValid_57 & _T_40155; // @[Switch.scala 30:36:@18858.4]
  assign _T_40158 = io_inAddr_58 == 6'h3a; // @[Switch.scala 30:53:@18860.4]
  assign valid_58_58 = io_inValid_58 & _T_40158; // @[Switch.scala 30:36:@18861.4]
  assign _T_40161 = io_inAddr_59 == 6'h3a; // @[Switch.scala 30:53:@18863.4]
  assign valid_58_59 = io_inValid_59 & _T_40161; // @[Switch.scala 30:36:@18864.4]
  assign _T_40164 = io_inAddr_60 == 6'h3a; // @[Switch.scala 30:53:@18866.4]
  assign valid_58_60 = io_inValid_60 & _T_40164; // @[Switch.scala 30:36:@18867.4]
  assign _T_40167 = io_inAddr_61 == 6'h3a; // @[Switch.scala 30:53:@18869.4]
  assign valid_58_61 = io_inValid_61 & _T_40167; // @[Switch.scala 30:36:@18870.4]
  assign _T_40170 = io_inAddr_62 == 6'h3a; // @[Switch.scala 30:53:@18872.4]
  assign valid_58_62 = io_inValid_62 & _T_40170; // @[Switch.scala 30:36:@18873.4]
  assign _T_40173 = io_inAddr_63 == 6'h3a; // @[Switch.scala 30:53:@18875.4]
  assign valid_58_63 = io_inValid_63 & _T_40173; // @[Switch.scala 30:36:@18876.4]
  assign _T_40239 = valid_58_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@18878.4]
  assign _T_40240 = valid_58_61 ? 6'h3d : _T_40239; // @[Mux.scala 31:69:@18879.4]
  assign _T_40241 = valid_58_60 ? 6'h3c : _T_40240; // @[Mux.scala 31:69:@18880.4]
  assign _T_40242 = valid_58_59 ? 6'h3b : _T_40241; // @[Mux.scala 31:69:@18881.4]
  assign _T_40243 = valid_58_58 ? 6'h3a : _T_40242; // @[Mux.scala 31:69:@18882.4]
  assign _T_40244 = valid_58_57 ? 6'h39 : _T_40243; // @[Mux.scala 31:69:@18883.4]
  assign _T_40245 = valid_58_56 ? 6'h38 : _T_40244; // @[Mux.scala 31:69:@18884.4]
  assign _T_40246 = valid_58_55 ? 6'h37 : _T_40245; // @[Mux.scala 31:69:@18885.4]
  assign _T_40247 = valid_58_54 ? 6'h36 : _T_40246; // @[Mux.scala 31:69:@18886.4]
  assign _T_40248 = valid_58_53 ? 6'h35 : _T_40247; // @[Mux.scala 31:69:@18887.4]
  assign _T_40249 = valid_58_52 ? 6'h34 : _T_40248; // @[Mux.scala 31:69:@18888.4]
  assign _T_40250 = valid_58_51 ? 6'h33 : _T_40249; // @[Mux.scala 31:69:@18889.4]
  assign _T_40251 = valid_58_50 ? 6'h32 : _T_40250; // @[Mux.scala 31:69:@18890.4]
  assign _T_40252 = valid_58_49 ? 6'h31 : _T_40251; // @[Mux.scala 31:69:@18891.4]
  assign _T_40253 = valid_58_48 ? 6'h30 : _T_40252; // @[Mux.scala 31:69:@18892.4]
  assign _T_40254 = valid_58_47 ? 6'h2f : _T_40253; // @[Mux.scala 31:69:@18893.4]
  assign _T_40255 = valid_58_46 ? 6'h2e : _T_40254; // @[Mux.scala 31:69:@18894.4]
  assign _T_40256 = valid_58_45 ? 6'h2d : _T_40255; // @[Mux.scala 31:69:@18895.4]
  assign _T_40257 = valid_58_44 ? 6'h2c : _T_40256; // @[Mux.scala 31:69:@18896.4]
  assign _T_40258 = valid_58_43 ? 6'h2b : _T_40257; // @[Mux.scala 31:69:@18897.4]
  assign _T_40259 = valid_58_42 ? 6'h2a : _T_40258; // @[Mux.scala 31:69:@18898.4]
  assign _T_40260 = valid_58_41 ? 6'h29 : _T_40259; // @[Mux.scala 31:69:@18899.4]
  assign _T_40261 = valid_58_40 ? 6'h28 : _T_40260; // @[Mux.scala 31:69:@18900.4]
  assign _T_40262 = valid_58_39 ? 6'h27 : _T_40261; // @[Mux.scala 31:69:@18901.4]
  assign _T_40263 = valid_58_38 ? 6'h26 : _T_40262; // @[Mux.scala 31:69:@18902.4]
  assign _T_40264 = valid_58_37 ? 6'h25 : _T_40263; // @[Mux.scala 31:69:@18903.4]
  assign _T_40265 = valid_58_36 ? 6'h24 : _T_40264; // @[Mux.scala 31:69:@18904.4]
  assign _T_40266 = valid_58_35 ? 6'h23 : _T_40265; // @[Mux.scala 31:69:@18905.4]
  assign _T_40267 = valid_58_34 ? 6'h22 : _T_40266; // @[Mux.scala 31:69:@18906.4]
  assign _T_40268 = valid_58_33 ? 6'h21 : _T_40267; // @[Mux.scala 31:69:@18907.4]
  assign _T_40269 = valid_58_32 ? 6'h20 : _T_40268; // @[Mux.scala 31:69:@18908.4]
  assign _T_40270 = valid_58_31 ? 6'h1f : _T_40269; // @[Mux.scala 31:69:@18909.4]
  assign _T_40271 = valid_58_30 ? 6'h1e : _T_40270; // @[Mux.scala 31:69:@18910.4]
  assign _T_40272 = valid_58_29 ? 6'h1d : _T_40271; // @[Mux.scala 31:69:@18911.4]
  assign _T_40273 = valid_58_28 ? 6'h1c : _T_40272; // @[Mux.scala 31:69:@18912.4]
  assign _T_40274 = valid_58_27 ? 6'h1b : _T_40273; // @[Mux.scala 31:69:@18913.4]
  assign _T_40275 = valid_58_26 ? 6'h1a : _T_40274; // @[Mux.scala 31:69:@18914.4]
  assign _T_40276 = valid_58_25 ? 6'h19 : _T_40275; // @[Mux.scala 31:69:@18915.4]
  assign _T_40277 = valid_58_24 ? 6'h18 : _T_40276; // @[Mux.scala 31:69:@18916.4]
  assign _T_40278 = valid_58_23 ? 6'h17 : _T_40277; // @[Mux.scala 31:69:@18917.4]
  assign _T_40279 = valid_58_22 ? 6'h16 : _T_40278; // @[Mux.scala 31:69:@18918.4]
  assign _T_40280 = valid_58_21 ? 6'h15 : _T_40279; // @[Mux.scala 31:69:@18919.4]
  assign _T_40281 = valid_58_20 ? 6'h14 : _T_40280; // @[Mux.scala 31:69:@18920.4]
  assign _T_40282 = valid_58_19 ? 6'h13 : _T_40281; // @[Mux.scala 31:69:@18921.4]
  assign _T_40283 = valid_58_18 ? 6'h12 : _T_40282; // @[Mux.scala 31:69:@18922.4]
  assign _T_40284 = valid_58_17 ? 6'h11 : _T_40283; // @[Mux.scala 31:69:@18923.4]
  assign _T_40285 = valid_58_16 ? 6'h10 : _T_40284; // @[Mux.scala 31:69:@18924.4]
  assign _T_40286 = valid_58_15 ? 6'hf : _T_40285; // @[Mux.scala 31:69:@18925.4]
  assign _T_40287 = valid_58_14 ? 6'he : _T_40286; // @[Mux.scala 31:69:@18926.4]
  assign _T_40288 = valid_58_13 ? 6'hd : _T_40287; // @[Mux.scala 31:69:@18927.4]
  assign _T_40289 = valid_58_12 ? 6'hc : _T_40288; // @[Mux.scala 31:69:@18928.4]
  assign _T_40290 = valid_58_11 ? 6'hb : _T_40289; // @[Mux.scala 31:69:@18929.4]
  assign _T_40291 = valid_58_10 ? 6'ha : _T_40290; // @[Mux.scala 31:69:@18930.4]
  assign _T_40292 = valid_58_9 ? 6'h9 : _T_40291; // @[Mux.scala 31:69:@18931.4]
  assign _T_40293 = valid_58_8 ? 6'h8 : _T_40292; // @[Mux.scala 31:69:@18932.4]
  assign _T_40294 = valid_58_7 ? 6'h7 : _T_40293; // @[Mux.scala 31:69:@18933.4]
  assign _T_40295 = valid_58_6 ? 6'h6 : _T_40294; // @[Mux.scala 31:69:@18934.4]
  assign _T_40296 = valid_58_5 ? 6'h5 : _T_40295; // @[Mux.scala 31:69:@18935.4]
  assign _T_40297 = valid_58_4 ? 6'h4 : _T_40296; // @[Mux.scala 31:69:@18936.4]
  assign _T_40298 = valid_58_3 ? 6'h3 : _T_40297; // @[Mux.scala 31:69:@18937.4]
  assign _T_40299 = valid_58_2 ? 6'h2 : _T_40298; // @[Mux.scala 31:69:@18938.4]
  assign _T_40300 = valid_58_1 ? 6'h1 : _T_40299; // @[Mux.scala 31:69:@18939.4]
  assign select_58 = valid_58_0 ? 6'h0 : _T_40300; // @[Mux.scala 31:69:@18940.4]
  assign _GEN_3713 = 6'h1 == select_58 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3714 = 6'h2 == select_58 ? io_inData_2 : _GEN_3713; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3715 = 6'h3 == select_58 ? io_inData_3 : _GEN_3714; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3716 = 6'h4 == select_58 ? io_inData_4 : _GEN_3715; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3717 = 6'h5 == select_58 ? io_inData_5 : _GEN_3716; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3718 = 6'h6 == select_58 ? io_inData_6 : _GEN_3717; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3719 = 6'h7 == select_58 ? io_inData_7 : _GEN_3718; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3720 = 6'h8 == select_58 ? io_inData_8 : _GEN_3719; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3721 = 6'h9 == select_58 ? io_inData_9 : _GEN_3720; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3722 = 6'ha == select_58 ? io_inData_10 : _GEN_3721; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3723 = 6'hb == select_58 ? io_inData_11 : _GEN_3722; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3724 = 6'hc == select_58 ? io_inData_12 : _GEN_3723; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3725 = 6'hd == select_58 ? io_inData_13 : _GEN_3724; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3726 = 6'he == select_58 ? io_inData_14 : _GEN_3725; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3727 = 6'hf == select_58 ? io_inData_15 : _GEN_3726; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3728 = 6'h10 == select_58 ? io_inData_16 : _GEN_3727; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3729 = 6'h11 == select_58 ? io_inData_17 : _GEN_3728; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3730 = 6'h12 == select_58 ? io_inData_18 : _GEN_3729; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3731 = 6'h13 == select_58 ? io_inData_19 : _GEN_3730; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3732 = 6'h14 == select_58 ? io_inData_20 : _GEN_3731; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3733 = 6'h15 == select_58 ? io_inData_21 : _GEN_3732; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3734 = 6'h16 == select_58 ? io_inData_22 : _GEN_3733; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3735 = 6'h17 == select_58 ? io_inData_23 : _GEN_3734; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3736 = 6'h18 == select_58 ? io_inData_24 : _GEN_3735; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3737 = 6'h19 == select_58 ? io_inData_25 : _GEN_3736; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3738 = 6'h1a == select_58 ? io_inData_26 : _GEN_3737; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3739 = 6'h1b == select_58 ? io_inData_27 : _GEN_3738; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3740 = 6'h1c == select_58 ? io_inData_28 : _GEN_3739; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3741 = 6'h1d == select_58 ? io_inData_29 : _GEN_3740; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3742 = 6'h1e == select_58 ? io_inData_30 : _GEN_3741; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3743 = 6'h1f == select_58 ? io_inData_31 : _GEN_3742; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3744 = 6'h20 == select_58 ? io_inData_32 : _GEN_3743; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3745 = 6'h21 == select_58 ? io_inData_33 : _GEN_3744; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3746 = 6'h22 == select_58 ? io_inData_34 : _GEN_3745; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3747 = 6'h23 == select_58 ? io_inData_35 : _GEN_3746; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3748 = 6'h24 == select_58 ? io_inData_36 : _GEN_3747; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3749 = 6'h25 == select_58 ? io_inData_37 : _GEN_3748; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3750 = 6'h26 == select_58 ? io_inData_38 : _GEN_3749; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3751 = 6'h27 == select_58 ? io_inData_39 : _GEN_3750; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3752 = 6'h28 == select_58 ? io_inData_40 : _GEN_3751; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3753 = 6'h29 == select_58 ? io_inData_41 : _GEN_3752; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3754 = 6'h2a == select_58 ? io_inData_42 : _GEN_3753; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3755 = 6'h2b == select_58 ? io_inData_43 : _GEN_3754; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3756 = 6'h2c == select_58 ? io_inData_44 : _GEN_3755; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3757 = 6'h2d == select_58 ? io_inData_45 : _GEN_3756; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3758 = 6'h2e == select_58 ? io_inData_46 : _GEN_3757; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3759 = 6'h2f == select_58 ? io_inData_47 : _GEN_3758; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3760 = 6'h30 == select_58 ? io_inData_48 : _GEN_3759; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3761 = 6'h31 == select_58 ? io_inData_49 : _GEN_3760; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3762 = 6'h32 == select_58 ? io_inData_50 : _GEN_3761; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3763 = 6'h33 == select_58 ? io_inData_51 : _GEN_3762; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3764 = 6'h34 == select_58 ? io_inData_52 : _GEN_3763; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3765 = 6'h35 == select_58 ? io_inData_53 : _GEN_3764; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3766 = 6'h36 == select_58 ? io_inData_54 : _GEN_3765; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3767 = 6'h37 == select_58 ? io_inData_55 : _GEN_3766; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3768 = 6'h38 == select_58 ? io_inData_56 : _GEN_3767; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3769 = 6'h39 == select_58 ? io_inData_57 : _GEN_3768; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3770 = 6'h3a == select_58 ? io_inData_58 : _GEN_3769; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3771 = 6'h3b == select_58 ? io_inData_59 : _GEN_3770; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3772 = 6'h3c == select_58 ? io_inData_60 : _GEN_3771; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3773 = 6'h3d == select_58 ? io_inData_61 : _GEN_3772; // @[Switch.scala 33:19:@18942.4]
  assign _GEN_3774 = 6'h3e == select_58 ? io_inData_62 : _GEN_3773; // @[Switch.scala 33:19:@18942.4]
  assign _T_40309 = {valid_58_7,valid_58_6,valid_58_5,valid_58_4,valid_58_3,valid_58_2,valid_58_1,valid_58_0}; // @[Switch.scala 34:32:@18949.4]
  assign _T_40317 = {valid_58_15,valid_58_14,valid_58_13,valid_58_12,valid_58_11,valid_58_10,valid_58_9,valid_58_8,_T_40309}; // @[Switch.scala 34:32:@18957.4]
  assign _T_40324 = {valid_58_23,valid_58_22,valid_58_21,valid_58_20,valid_58_19,valid_58_18,valid_58_17,valid_58_16}; // @[Switch.scala 34:32:@18964.4]
  assign _T_40333 = {valid_58_31,valid_58_30,valid_58_29,valid_58_28,valid_58_27,valid_58_26,valid_58_25,valid_58_24,_T_40324,_T_40317}; // @[Switch.scala 34:32:@18973.4]
  assign _T_40340 = {valid_58_39,valid_58_38,valid_58_37,valid_58_36,valid_58_35,valid_58_34,valid_58_33,valid_58_32}; // @[Switch.scala 34:32:@18980.4]
  assign _T_40348 = {valid_58_47,valid_58_46,valid_58_45,valid_58_44,valid_58_43,valid_58_42,valid_58_41,valid_58_40,_T_40340}; // @[Switch.scala 34:32:@18988.4]
  assign _T_40355 = {valid_58_55,valid_58_54,valid_58_53,valid_58_52,valid_58_51,valid_58_50,valid_58_49,valid_58_48}; // @[Switch.scala 34:32:@18995.4]
  assign _T_40364 = {valid_58_63,valid_58_62,valid_58_61,valid_58_60,valid_58_59,valid_58_58,valid_58_57,valid_58_56,_T_40355,_T_40348}; // @[Switch.scala 34:32:@19004.4]
  assign _T_40365 = {_T_40364,_T_40333}; // @[Switch.scala 34:32:@19005.4]
  assign _T_40369 = io_inAddr_0 == 6'h3b; // @[Switch.scala 30:53:@19008.4]
  assign valid_59_0 = io_inValid_0 & _T_40369; // @[Switch.scala 30:36:@19009.4]
  assign _T_40372 = io_inAddr_1 == 6'h3b; // @[Switch.scala 30:53:@19011.4]
  assign valid_59_1 = io_inValid_1 & _T_40372; // @[Switch.scala 30:36:@19012.4]
  assign _T_40375 = io_inAddr_2 == 6'h3b; // @[Switch.scala 30:53:@19014.4]
  assign valid_59_2 = io_inValid_2 & _T_40375; // @[Switch.scala 30:36:@19015.4]
  assign _T_40378 = io_inAddr_3 == 6'h3b; // @[Switch.scala 30:53:@19017.4]
  assign valid_59_3 = io_inValid_3 & _T_40378; // @[Switch.scala 30:36:@19018.4]
  assign _T_40381 = io_inAddr_4 == 6'h3b; // @[Switch.scala 30:53:@19020.4]
  assign valid_59_4 = io_inValid_4 & _T_40381; // @[Switch.scala 30:36:@19021.4]
  assign _T_40384 = io_inAddr_5 == 6'h3b; // @[Switch.scala 30:53:@19023.4]
  assign valid_59_5 = io_inValid_5 & _T_40384; // @[Switch.scala 30:36:@19024.4]
  assign _T_40387 = io_inAddr_6 == 6'h3b; // @[Switch.scala 30:53:@19026.4]
  assign valid_59_6 = io_inValid_6 & _T_40387; // @[Switch.scala 30:36:@19027.4]
  assign _T_40390 = io_inAddr_7 == 6'h3b; // @[Switch.scala 30:53:@19029.4]
  assign valid_59_7 = io_inValid_7 & _T_40390; // @[Switch.scala 30:36:@19030.4]
  assign _T_40393 = io_inAddr_8 == 6'h3b; // @[Switch.scala 30:53:@19032.4]
  assign valid_59_8 = io_inValid_8 & _T_40393; // @[Switch.scala 30:36:@19033.4]
  assign _T_40396 = io_inAddr_9 == 6'h3b; // @[Switch.scala 30:53:@19035.4]
  assign valid_59_9 = io_inValid_9 & _T_40396; // @[Switch.scala 30:36:@19036.4]
  assign _T_40399 = io_inAddr_10 == 6'h3b; // @[Switch.scala 30:53:@19038.4]
  assign valid_59_10 = io_inValid_10 & _T_40399; // @[Switch.scala 30:36:@19039.4]
  assign _T_40402 = io_inAddr_11 == 6'h3b; // @[Switch.scala 30:53:@19041.4]
  assign valid_59_11 = io_inValid_11 & _T_40402; // @[Switch.scala 30:36:@19042.4]
  assign _T_40405 = io_inAddr_12 == 6'h3b; // @[Switch.scala 30:53:@19044.4]
  assign valid_59_12 = io_inValid_12 & _T_40405; // @[Switch.scala 30:36:@19045.4]
  assign _T_40408 = io_inAddr_13 == 6'h3b; // @[Switch.scala 30:53:@19047.4]
  assign valid_59_13 = io_inValid_13 & _T_40408; // @[Switch.scala 30:36:@19048.4]
  assign _T_40411 = io_inAddr_14 == 6'h3b; // @[Switch.scala 30:53:@19050.4]
  assign valid_59_14 = io_inValid_14 & _T_40411; // @[Switch.scala 30:36:@19051.4]
  assign _T_40414 = io_inAddr_15 == 6'h3b; // @[Switch.scala 30:53:@19053.4]
  assign valid_59_15 = io_inValid_15 & _T_40414; // @[Switch.scala 30:36:@19054.4]
  assign _T_40417 = io_inAddr_16 == 6'h3b; // @[Switch.scala 30:53:@19056.4]
  assign valid_59_16 = io_inValid_16 & _T_40417; // @[Switch.scala 30:36:@19057.4]
  assign _T_40420 = io_inAddr_17 == 6'h3b; // @[Switch.scala 30:53:@19059.4]
  assign valid_59_17 = io_inValid_17 & _T_40420; // @[Switch.scala 30:36:@19060.4]
  assign _T_40423 = io_inAddr_18 == 6'h3b; // @[Switch.scala 30:53:@19062.4]
  assign valid_59_18 = io_inValid_18 & _T_40423; // @[Switch.scala 30:36:@19063.4]
  assign _T_40426 = io_inAddr_19 == 6'h3b; // @[Switch.scala 30:53:@19065.4]
  assign valid_59_19 = io_inValid_19 & _T_40426; // @[Switch.scala 30:36:@19066.4]
  assign _T_40429 = io_inAddr_20 == 6'h3b; // @[Switch.scala 30:53:@19068.4]
  assign valid_59_20 = io_inValid_20 & _T_40429; // @[Switch.scala 30:36:@19069.4]
  assign _T_40432 = io_inAddr_21 == 6'h3b; // @[Switch.scala 30:53:@19071.4]
  assign valid_59_21 = io_inValid_21 & _T_40432; // @[Switch.scala 30:36:@19072.4]
  assign _T_40435 = io_inAddr_22 == 6'h3b; // @[Switch.scala 30:53:@19074.4]
  assign valid_59_22 = io_inValid_22 & _T_40435; // @[Switch.scala 30:36:@19075.4]
  assign _T_40438 = io_inAddr_23 == 6'h3b; // @[Switch.scala 30:53:@19077.4]
  assign valid_59_23 = io_inValid_23 & _T_40438; // @[Switch.scala 30:36:@19078.4]
  assign _T_40441 = io_inAddr_24 == 6'h3b; // @[Switch.scala 30:53:@19080.4]
  assign valid_59_24 = io_inValid_24 & _T_40441; // @[Switch.scala 30:36:@19081.4]
  assign _T_40444 = io_inAddr_25 == 6'h3b; // @[Switch.scala 30:53:@19083.4]
  assign valid_59_25 = io_inValid_25 & _T_40444; // @[Switch.scala 30:36:@19084.4]
  assign _T_40447 = io_inAddr_26 == 6'h3b; // @[Switch.scala 30:53:@19086.4]
  assign valid_59_26 = io_inValid_26 & _T_40447; // @[Switch.scala 30:36:@19087.4]
  assign _T_40450 = io_inAddr_27 == 6'h3b; // @[Switch.scala 30:53:@19089.4]
  assign valid_59_27 = io_inValid_27 & _T_40450; // @[Switch.scala 30:36:@19090.4]
  assign _T_40453 = io_inAddr_28 == 6'h3b; // @[Switch.scala 30:53:@19092.4]
  assign valid_59_28 = io_inValid_28 & _T_40453; // @[Switch.scala 30:36:@19093.4]
  assign _T_40456 = io_inAddr_29 == 6'h3b; // @[Switch.scala 30:53:@19095.4]
  assign valid_59_29 = io_inValid_29 & _T_40456; // @[Switch.scala 30:36:@19096.4]
  assign _T_40459 = io_inAddr_30 == 6'h3b; // @[Switch.scala 30:53:@19098.4]
  assign valid_59_30 = io_inValid_30 & _T_40459; // @[Switch.scala 30:36:@19099.4]
  assign _T_40462 = io_inAddr_31 == 6'h3b; // @[Switch.scala 30:53:@19101.4]
  assign valid_59_31 = io_inValid_31 & _T_40462; // @[Switch.scala 30:36:@19102.4]
  assign _T_40465 = io_inAddr_32 == 6'h3b; // @[Switch.scala 30:53:@19104.4]
  assign valid_59_32 = io_inValid_32 & _T_40465; // @[Switch.scala 30:36:@19105.4]
  assign _T_40468 = io_inAddr_33 == 6'h3b; // @[Switch.scala 30:53:@19107.4]
  assign valid_59_33 = io_inValid_33 & _T_40468; // @[Switch.scala 30:36:@19108.4]
  assign _T_40471 = io_inAddr_34 == 6'h3b; // @[Switch.scala 30:53:@19110.4]
  assign valid_59_34 = io_inValid_34 & _T_40471; // @[Switch.scala 30:36:@19111.4]
  assign _T_40474 = io_inAddr_35 == 6'h3b; // @[Switch.scala 30:53:@19113.4]
  assign valid_59_35 = io_inValid_35 & _T_40474; // @[Switch.scala 30:36:@19114.4]
  assign _T_40477 = io_inAddr_36 == 6'h3b; // @[Switch.scala 30:53:@19116.4]
  assign valid_59_36 = io_inValid_36 & _T_40477; // @[Switch.scala 30:36:@19117.4]
  assign _T_40480 = io_inAddr_37 == 6'h3b; // @[Switch.scala 30:53:@19119.4]
  assign valid_59_37 = io_inValid_37 & _T_40480; // @[Switch.scala 30:36:@19120.4]
  assign _T_40483 = io_inAddr_38 == 6'h3b; // @[Switch.scala 30:53:@19122.4]
  assign valid_59_38 = io_inValid_38 & _T_40483; // @[Switch.scala 30:36:@19123.4]
  assign _T_40486 = io_inAddr_39 == 6'h3b; // @[Switch.scala 30:53:@19125.4]
  assign valid_59_39 = io_inValid_39 & _T_40486; // @[Switch.scala 30:36:@19126.4]
  assign _T_40489 = io_inAddr_40 == 6'h3b; // @[Switch.scala 30:53:@19128.4]
  assign valid_59_40 = io_inValid_40 & _T_40489; // @[Switch.scala 30:36:@19129.4]
  assign _T_40492 = io_inAddr_41 == 6'h3b; // @[Switch.scala 30:53:@19131.4]
  assign valid_59_41 = io_inValid_41 & _T_40492; // @[Switch.scala 30:36:@19132.4]
  assign _T_40495 = io_inAddr_42 == 6'h3b; // @[Switch.scala 30:53:@19134.4]
  assign valid_59_42 = io_inValid_42 & _T_40495; // @[Switch.scala 30:36:@19135.4]
  assign _T_40498 = io_inAddr_43 == 6'h3b; // @[Switch.scala 30:53:@19137.4]
  assign valid_59_43 = io_inValid_43 & _T_40498; // @[Switch.scala 30:36:@19138.4]
  assign _T_40501 = io_inAddr_44 == 6'h3b; // @[Switch.scala 30:53:@19140.4]
  assign valid_59_44 = io_inValid_44 & _T_40501; // @[Switch.scala 30:36:@19141.4]
  assign _T_40504 = io_inAddr_45 == 6'h3b; // @[Switch.scala 30:53:@19143.4]
  assign valid_59_45 = io_inValid_45 & _T_40504; // @[Switch.scala 30:36:@19144.4]
  assign _T_40507 = io_inAddr_46 == 6'h3b; // @[Switch.scala 30:53:@19146.4]
  assign valid_59_46 = io_inValid_46 & _T_40507; // @[Switch.scala 30:36:@19147.4]
  assign _T_40510 = io_inAddr_47 == 6'h3b; // @[Switch.scala 30:53:@19149.4]
  assign valid_59_47 = io_inValid_47 & _T_40510; // @[Switch.scala 30:36:@19150.4]
  assign _T_40513 = io_inAddr_48 == 6'h3b; // @[Switch.scala 30:53:@19152.4]
  assign valid_59_48 = io_inValid_48 & _T_40513; // @[Switch.scala 30:36:@19153.4]
  assign _T_40516 = io_inAddr_49 == 6'h3b; // @[Switch.scala 30:53:@19155.4]
  assign valid_59_49 = io_inValid_49 & _T_40516; // @[Switch.scala 30:36:@19156.4]
  assign _T_40519 = io_inAddr_50 == 6'h3b; // @[Switch.scala 30:53:@19158.4]
  assign valid_59_50 = io_inValid_50 & _T_40519; // @[Switch.scala 30:36:@19159.4]
  assign _T_40522 = io_inAddr_51 == 6'h3b; // @[Switch.scala 30:53:@19161.4]
  assign valid_59_51 = io_inValid_51 & _T_40522; // @[Switch.scala 30:36:@19162.4]
  assign _T_40525 = io_inAddr_52 == 6'h3b; // @[Switch.scala 30:53:@19164.4]
  assign valid_59_52 = io_inValid_52 & _T_40525; // @[Switch.scala 30:36:@19165.4]
  assign _T_40528 = io_inAddr_53 == 6'h3b; // @[Switch.scala 30:53:@19167.4]
  assign valid_59_53 = io_inValid_53 & _T_40528; // @[Switch.scala 30:36:@19168.4]
  assign _T_40531 = io_inAddr_54 == 6'h3b; // @[Switch.scala 30:53:@19170.4]
  assign valid_59_54 = io_inValid_54 & _T_40531; // @[Switch.scala 30:36:@19171.4]
  assign _T_40534 = io_inAddr_55 == 6'h3b; // @[Switch.scala 30:53:@19173.4]
  assign valid_59_55 = io_inValid_55 & _T_40534; // @[Switch.scala 30:36:@19174.4]
  assign _T_40537 = io_inAddr_56 == 6'h3b; // @[Switch.scala 30:53:@19176.4]
  assign valid_59_56 = io_inValid_56 & _T_40537; // @[Switch.scala 30:36:@19177.4]
  assign _T_40540 = io_inAddr_57 == 6'h3b; // @[Switch.scala 30:53:@19179.4]
  assign valid_59_57 = io_inValid_57 & _T_40540; // @[Switch.scala 30:36:@19180.4]
  assign _T_40543 = io_inAddr_58 == 6'h3b; // @[Switch.scala 30:53:@19182.4]
  assign valid_59_58 = io_inValid_58 & _T_40543; // @[Switch.scala 30:36:@19183.4]
  assign _T_40546 = io_inAddr_59 == 6'h3b; // @[Switch.scala 30:53:@19185.4]
  assign valid_59_59 = io_inValid_59 & _T_40546; // @[Switch.scala 30:36:@19186.4]
  assign _T_40549 = io_inAddr_60 == 6'h3b; // @[Switch.scala 30:53:@19188.4]
  assign valid_59_60 = io_inValid_60 & _T_40549; // @[Switch.scala 30:36:@19189.4]
  assign _T_40552 = io_inAddr_61 == 6'h3b; // @[Switch.scala 30:53:@19191.4]
  assign valid_59_61 = io_inValid_61 & _T_40552; // @[Switch.scala 30:36:@19192.4]
  assign _T_40555 = io_inAddr_62 == 6'h3b; // @[Switch.scala 30:53:@19194.4]
  assign valid_59_62 = io_inValid_62 & _T_40555; // @[Switch.scala 30:36:@19195.4]
  assign _T_40558 = io_inAddr_63 == 6'h3b; // @[Switch.scala 30:53:@19197.4]
  assign valid_59_63 = io_inValid_63 & _T_40558; // @[Switch.scala 30:36:@19198.4]
  assign _T_40624 = valid_59_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@19200.4]
  assign _T_40625 = valid_59_61 ? 6'h3d : _T_40624; // @[Mux.scala 31:69:@19201.4]
  assign _T_40626 = valid_59_60 ? 6'h3c : _T_40625; // @[Mux.scala 31:69:@19202.4]
  assign _T_40627 = valid_59_59 ? 6'h3b : _T_40626; // @[Mux.scala 31:69:@19203.4]
  assign _T_40628 = valid_59_58 ? 6'h3a : _T_40627; // @[Mux.scala 31:69:@19204.4]
  assign _T_40629 = valid_59_57 ? 6'h39 : _T_40628; // @[Mux.scala 31:69:@19205.4]
  assign _T_40630 = valid_59_56 ? 6'h38 : _T_40629; // @[Mux.scala 31:69:@19206.4]
  assign _T_40631 = valid_59_55 ? 6'h37 : _T_40630; // @[Mux.scala 31:69:@19207.4]
  assign _T_40632 = valid_59_54 ? 6'h36 : _T_40631; // @[Mux.scala 31:69:@19208.4]
  assign _T_40633 = valid_59_53 ? 6'h35 : _T_40632; // @[Mux.scala 31:69:@19209.4]
  assign _T_40634 = valid_59_52 ? 6'h34 : _T_40633; // @[Mux.scala 31:69:@19210.4]
  assign _T_40635 = valid_59_51 ? 6'h33 : _T_40634; // @[Mux.scala 31:69:@19211.4]
  assign _T_40636 = valid_59_50 ? 6'h32 : _T_40635; // @[Mux.scala 31:69:@19212.4]
  assign _T_40637 = valid_59_49 ? 6'h31 : _T_40636; // @[Mux.scala 31:69:@19213.4]
  assign _T_40638 = valid_59_48 ? 6'h30 : _T_40637; // @[Mux.scala 31:69:@19214.4]
  assign _T_40639 = valid_59_47 ? 6'h2f : _T_40638; // @[Mux.scala 31:69:@19215.4]
  assign _T_40640 = valid_59_46 ? 6'h2e : _T_40639; // @[Mux.scala 31:69:@19216.4]
  assign _T_40641 = valid_59_45 ? 6'h2d : _T_40640; // @[Mux.scala 31:69:@19217.4]
  assign _T_40642 = valid_59_44 ? 6'h2c : _T_40641; // @[Mux.scala 31:69:@19218.4]
  assign _T_40643 = valid_59_43 ? 6'h2b : _T_40642; // @[Mux.scala 31:69:@19219.4]
  assign _T_40644 = valid_59_42 ? 6'h2a : _T_40643; // @[Mux.scala 31:69:@19220.4]
  assign _T_40645 = valid_59_41 ? 6'h29 : _T_40644; // @[Mux.scala 31:69:@19221.4]
  assign _T_40646 = valid_59_40 ? 6'h28 : _T_40645; // @[Mux.scala 31:69:@19222.4]
  assign _T_40647 = valid_59_39 ? 6'h27 : _T_40646; // @[Mux.scala 31:69:@19223.4]
  assign _T_40648 = valid_59_38 ? 6'h26 : _T_40647; // @[Mux.scala 31:69:@19224.4]
  assign _T_40649 = valid_59_37 ? 6'h25 : _T_40648; // @[Mux.scala 31:69:@19225.4]
  assign _T_40650 = valid_59_36 ? 6'h24 : _T_40649; // @[Mux.scala 31:69:@19226.4]
  assign _T_40651 = valid_59_35 ? 6'h23 : _T_40650; // @[Mux.scala 31:69:@19227.4]
  assign _T_40652 = valid_59_34 ? 6'h22 : _T_40651; // @[Mux.scala 31:69:@19228.4]
  assign _T_40653 = valid_59_33 ? 6'h21 : _T_40652; // @[Mux.scala 31:69:@19229.4]
  assign _T_40654 = valid_59_32 ? 6'h20 : _T_40653; // @[Mux.scala 31:69:@19230.4]
  assign _T_40655 = valid_59_31 ? 6'h1f : _T_40654; // @[Mux.scala 31:69:@19231.4]
  assign _T_40656 = valid_59_30 ? 6'h1e : _T_40655; // @[Mux.scala 31:69:@19232.4]
  assign _T_40657 = valid_59_29 ? 6'h1d : _T_40656; // @[Mux.scala 31:69:@19233.4]
  assign _T_40658 = valid_59_28 ? 6'h1c : _T_40657; // @[Mux.scala 31:69:@19234.4]
  assign _T_40659 = valid_59_27 ? 6'h1b : _T_40658; // @[Mux.scala 31:69:@19235.4]
  assign _T_40660 = valid_59_26 ? 6'h1a : _T_40659; // @[Mux.scala 31:69:@19236.4]
  assign _T_40661 = valid_59_25 ? 6'h19 : _T_40660; // @[Mux.scala 31:69:@19237.4]
  assign _T_40662 = valid_59_24 ? 6'h18 : _T_40661; // @[Mux.scala 31:69:@19238.4]
  assign _T_40663 = valid_59_23 ? 6'h17 : _T_40662; // @[Mux.scala 31:69:@19239.4]
  assign _T_40664 = valid_59_22 ? 6'h16 : _T_40663; // @[Mux.scala 31:69:@19240.4]
  assign _T_40665 = valid_59_21 ? 6'h15 : _T_40664; // @[Mux.scala 31:69:@19241.4]
  assign _T_40666 = valid_59_20 ? 6'h14 : _T_40665; // @[Mux.scala 31:69:@19242.4]
  assign _T_40667 = valid_59_19 ? 6'h13 : _T_40666; // @[Mux.scala 31:69:@19243.4]
  assign _T_40668 = valid_59_18 ? 6'h12 : _T_40667; // @[Mux.scala 31:69:@19244.4]
  assign _T_40669 = valid_59_17 ? 6'h11 : _T_40668; // @[Mux.scala 31:69:@19245.4]
  assign _T_40670 = valid_59_16 ? 6'h10 : _T_40669; // @[Mux.scala 31:69:@19246.4]
  assign _T_40671 = valid_59_15 ? 6'hf : _T_40670; // @[Mux.scala 31:69:@19247.4]
  assign _T_40672 = valid_59_14 ? 6'he : _T_40671; // @[Mux.scala 31:69:@19248.4]
  assign _T_40673 = valid_59_13 ? 6'hd : _T_40672; // @[Mux.scala 31:69:@19249.4]
  assign _T_40674 = valid_59_12 ? 6'hc : _T_40673; // @[Mux.scala 31:69:@19250.4]
  assign _T_40675 = valid_59_11 ? 6'hb : _T_40674; // @[Mux.scala 31:69:@19251.4]
  assign _T_40676 = valid_59_10 ? 6'ha : _T_40675; // @[Mux.scala 31:69:@19252.4]
  assign _T_40677 = valid_59_9 ? 6'h9 : _T_40676; // @[Mux.scala 31:69:@19253.4]
  assign _T_40678 = valid_59_8 ? 6'h8 : _T_40677; // @[Mux.scala 31:69:@19254.4]
  assign _T_40679 = valid_59_7 ? 6'h7 : _T_40678; // @[Mux.scala 31:69:@19255.4]
  assign _T_40680 = valid_59_6 ? 6'h6 : _T_40679; // @[Mux.scala 31:69:@19256.4]
  assign _T_40681 = valid_59_5 ? 6'h5 : _T_40680; // @[Mux.scala 31:69:@19257.4]
  assign _T_40682 = valid_59_4 ? 6'h4 : _T_40681; // @[Mux.scala 31:69:@19258.4]
  assign _T_40683 = valid_59_3 ? 6'h3 : _T_40682; // @[Mux.scala 31:69:@19259.4]
  assign _T_40684 = valid_59_2 ? 6'h2 : _T_40683; // @[Mux.scala 31:69:@19260.4]
  assign _T_40685 = valid_59_1 ? 6'h1 : _T_40684; // @[Mux.scala 31:69:@19261.4]
  assign select_59 = valid_59_0 ? 6'h0 : _T_40685; // @[Mux.scala 31:69:@19262.4]
  assign _GEN_3777 = 6'h1 == select_59 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3778 = 6'h2 == select_59 ? io_inData_2 : _GEN_3777; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3779 = 6'h3 == select_59 ? io_inData_3 : _GEN_3778; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3780 = 6'h4 == select_59 ? io_inData_4 : _GEN_3779; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3781 = 6'h5 == select_59 ? io_inData_5 : _GEN_3780; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3782 = 6'h6 == select_59 ? io_inData_6 : _GEN_3781; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3783 = 6'h7 == select_59 ? io_inData_7 : _GEN_3782; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3784 = 6'h8 == select_59 ? io_inData_8 : _GEN_3783; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3785 = 6'h9 == select_59 ? io_inData_9 : _GEN_3784; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3786 = 6'ha == select_59 ? io_inData_10 : _GEN_3785; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3787 = 6'hb == select_59 ? io_inData_11 : _GEN_3786; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3788 = 6'hc == select_59 ? io_inData_12 : _GEN_3787; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3789 = 6'hd == select_59 ? io_inData_13 : _GEN_3788; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3790 = 6'he == select_59 ? io_inData_14 : _GEN_3789; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3791 = 6'hf == select_59 ? io_inData_15 : _GEN_3790; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3792 = 6'h10 == select_59 ? io_inData_16 : _GEN_3791; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3793 = 6'h11 == select_59 ? io_inData_17 : _GEN_3792; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3794 = 6'h12 == select_59 ? io_inData_18 : _GEN_3793; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3795 = 6'h13 == select_59 ? io_inData_19 : _GEN_3794; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3796 = 6'h14 == select_59 ? io_inData_20 : _GEN_3795; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3797 = 6'h15 == select_59 ? io_inData_21 : _GEN_3796; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3798 = 6'h16 == select_59 ? io_inData_22 : _GEN_3797; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3799 = 6'h17 == select_59 ? io_inData_23 : _GEN_3798; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3800 = 6'h18 == select_59 ? io_inData_24 : _GEN_3799; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3801 = 6'h19 == select_59 ? io_inData_25 : _GEN_3800; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3802 = 6'h1a == select_59 ? io_inData_26 : _GEN_3801; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3803 = 6'h1b == select_59 ? io_inData_27 : _GEN_3802; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3804 = 6'h1c == select_59 ? io_inData_28 : _GEN_3803; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3805 = 6'h1d == select_59 ? io_inData_29 : _GEN_3804; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3806 = 6'h1e == select_59 ? io_inData_30 : _GEN_3805; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3807 = 6'h1f == select_59 ? io_inData_31 : _GEN_3806; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3808 = 6'h20 == select_59 ? io_inData_32 : _GEN_3807; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3809 = 6'h21 == select_59 ? io_inData_33 : _GEN_3808; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3810 = 6'h22 == select_59 ? io_inData_34 : _GEN_3809; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3811 = 6'h23 == select_59 ? io_inData_35 : _GEN_3810; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3812 = 6'h24 == select_59 ? io_inData_36 : _GEN_3811; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3813 = 6'h25 == select_59 ? io_inData_37 : _GEN_3812; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3814 = 6'h26 == select_59 ? io_inData_38 : _GEN_3813; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3815 = 6'h27 == select_59 ? io_inData_39 : _GEN_3814; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3816 = 6'h28 == select_59 ? io_inData_40 : _GEN_3815; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3817 = 6'h29 == select_59 ? io_inData_41 : _GEN_3816; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3818 = 6'h2a == select_59 ? io_inData_42 : _GEN_3817; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3819 = 6'h2b == select_59 ? io_inData_43 : _GEN_3818; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3820 = 6'h2c == select_59 ? io_inData_44 : _GEN_3819; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3821 = 6'h2d == select_59 ? io_inData_45 : _GEN_3820; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3822 = 6'h2e == select_59 ? io_inData_46 : _GEN_3821; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3823 = 6'h2f == select_59 ? io_inData_47 : _GEN_3822; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3824 = 6'h30 == select_59 ? io_inData_48 : _GEN_3823; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3825 = 6'h31 == select_59 ? io_inData_49 : _GEN_3824; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3826 = 6'h32 == select_59 ? io_inData_50 : _GEN_3825; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3827 = 6'h33 == select_59 ? io_inData_51 : _GEN_3826; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3828 = 6'h34 == select_59 ? io_inData_52 : _GEN_3827; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3829 = 6'h35 == select_59 ? io_inData_53 : _GEN_3828; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3830 = 6'h36 == select_59 ? io_inData_54 : _GEN_3829; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3831 = 6'h37 == select_59 ? io_inData_55 : _GEN_3830; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3832 = 6'h38 == select_59 ? io_inData_56 : _GEN_3831; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3833 = 6'h39 == select_59 ? io_inData_57 : _GEN_3832; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3834 = 6'h3a == select_59 ? io_inData_58 : _GEN_3833; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3835 = 6'h3b == select_59 ? io_inData_59 : _GEN_3834; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3836 = 6'h3c == select_59 ? io_inData_60 : _GEN_3835; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3837 = 6'h3d == select_59 ? io_inData_61 : _GEN_3836; // @[Switch.scala 33:19:@19264.4]
  assign _GEN_3838 = 6'h3e == select_59 ? io_inData_62 : _GEN_3837; // @[Switch.scala 33:19:@19264.4]
  assign _T_40694 = {valid_59_7,valid_59_6,valid_59_5,valid_59_4,valid_59_3,valid_59_2,valid_59_1,valid_59_0}; // @[Switch.scala 34:32:@19271.4]
  assign _T_40702 = {valid_59_15,valid_59_14,valid_59_13,valid_59_12,valid_59_11,valid_59_10,valid_59_9,valid_59_8,_T_40694}; // @[Switch.scala 34:32:@19279.4]
  assign _T_40709 = {valid_59_23,valid_59_22,valid_59_21,valid_59_20,valid_59_19,valid_59_18,valid_59_17,valid_59_16}; // @[Switch.scala 34:32:@19286.4]
  assign _T_40718 = {valid_59_31,valid_59_30,valid_59_29,valid_59_28,valid_59_27,valid_59_26,valid_59_25,valid_59_24,_T_40709,_T_40702}; // @[Switch.scala 34:32:@19295.4]
  assign _T_40725 = {valid_59_39,valid_59_38,valid_59_37,valid_59_36,valid_59_35,valid_59_34,valid_59_33,valid_59_32}; // @[Switch.scala 34:32:@19302.4]
  assign _T_40733 = {valid_59_47,valid_59_46,valid_59_45,valid_59_44,valid_59_43,valid_59_42,valid_59_41,valid_59_40,_T_40725}; // @[Switch.scala 34:32:@19310.4]
  assign _T_40740 = {valid_59_55,valid_59_54,valid_59_53,valid_59_52,valid_59_51,valid_59_50,valid_59_49,valid_59_48}; // @[Switch.scala 34:32:@19317.4]
  assign _T_40749 = {valid_59_63,valid_59_62,valid_59_61,valid_59_60,valid_59_59,valid_59_58,valid_59_57,valid_59_56,_T_40740,_T_40733}; // @[Switch.scala 34:32:@19326.4]
  assign _T_40750 = {_T_40749,_T_40718}; // @[Switch.scala 34:32:@19327.4]
  assign _T_40754 = io_inAddr_0 == 6'h3c; // @[Switch.scala 30:53:@19330.4]
  assign valid_60_0 = io_inValid_0 & _T_40754; // @[Switch.scala 30:36:@19331.4]
  assign _T_40757 = io_inAddr_1 == 6'h3c; // @[Switch.scala 30:53:@19333.4]
  assign valid_60_1 = io_inValid_1 & _T_40757; // @[Switch.scala 30:36:@19334.4]
  assign _T_40760 = io_inAddr_2 == 6'h3c; // @[Switch.scala 30:53:@19336.4]
  assign valid_60_2 = io_inValid_2 & _T_40760; // @[Switch.scala 30:36:@19337.4]
  assign _T_40763 = io_inAddr_3 == 6'h3c; // @[Switch.scala 30:53:@19339.4]
  assign valid_60_3 = io_inValid_3 & _T_40763; // @[Switch.scala 30:36:@19340.4]
  assign _T_40766 = io_inAddr_4 == 6'h3c; // @[Switch.scala 30:53:@19342.4]
  assign valid_60_4 = io_inValid_4 & _T_40766; // @[Switch.scala 30:36:@19343.4]
  assign _T_40769 = io_inAddr_5 == 6'h3c; // @[Switch.scala 30:53:@19345.4]
  assign valid_60_5 = io_inValid_5 & _T_40769; // @[Switch.scala 30:36:@19346.4]
  assign _T_40772 = io_inAddr_6 == 6'h3c; // @[Switch.scala 30:53:@19348.4]
  assign valid_60_6 = io_inValid_6 & _T_40772; // @[Switch.scala 30:36:@19349.4]
  assign _T_40775 = io_inAddr_7 == 6'h3c; // @[Switch.scala 30:53:@19351.4]
  assign valid_60_7 = io_inValid_7 & _T_40775; // @[Switch.scala 30:36:@19352.4]
  assign _T_40778 = io_inAddr_8 == 6'h3c; // @[Switch.scala 30:53:@19354.4]
  assign valid_60_8 = io_inValid_8 & _T_40778; // @[Switch.scala 30:36:@19355.4]
  assign _T_40781 = io_inAddr_9 == 6'h3c; // @[Switch.scala 30:53:@19357.4]
  assign valid_60_9 = io_inValid_9 & _T_40781; // @[Switch.scala 30:36:@19358.4]
  assign _T_40784 = io_inAddr_10 == 6'h3c; // @[Switch.scala 30:53:@19360.4]
  assign valid_60_10 = io_inValid_10 & _T_40784; // @[Switch.scala 30:36:@19361.4]
  assign _T_40787 = io_inAddr_11 == 6'h3c; // @[Switch.scala 30:53:@19363.4]
  assign valid_60_11 = io_inValid_11 & _T_40787; // @[Switch.scala 30:36:@19364.4]
  assign _T_40790 = io_inAddr_12 == 6'h3c; // @[Switch.scala 30:53:@19366.4]
  assign valid_60_12 = io_inValid_12 & _T_40790; // @[Switch.scala 30:36:@19367.4]
  assign _T_40793 = io_inAddr_13 == 6'h3c; // @[Switch.scala 30:53:@19369.4]
  assign valid_60_13 = io_inValid_13 & _T_40793; // @[Switch.scala 30:36:@19370.4]
  assign _T_40796 = io_inAddr_14 == 6'h3c; // @[Switch.scala 30:53:@19372.4]
  assign valid_60_14 = io_inValid_14 & _T_40796; // @[Switch.scala 30:36:@19373.4]
  assign _T_40799 = io_inAddr_15 == 6'h3c; // @[Switch.scala 30:53:@19375.4]
  assign valid_60_15 = io_inValid_15 & _T_40799; // @[Switch.scala 30:36:@19376.4]
  assign _T_40802 = io_inAddr_16 == 6'h3c; // @[Switch.scala 30:53:@19378.4]
  assign valid_60_16 = io_inValid_16 & _T_40802; // @[Switch.scala 30:36:@19379.4]
  assign _T_40805 = io_inAddr_17 == 6'h3c; // @[Switch.scala 30:53:@19381.4]
  assign valid_60_17 = io_inValid_17 & _T_40805; // @[Switch.scala 30:36:@19382.4]
  assign _T_40808 = io_inAddr_18 == 6'h3c; // @[Switch.scala 30:53:@19384.4]
  assign valid_60_18 = io_inValid_18 & _T_40808; // @[Switch.scala 30:36:@19385.4]
  assign _T_40811 = io_inAddr_19 == 6'h3c; // @[Switch.scala 30:53:@19387.4]
  assign valid_60_19 = io_inValid_19 & _T_40811; // @[Switch.scala 30:36:@19388.4]
  assign _T_40814 = io_inAddr_20 == 6'h3c; // @[Switch.scala 30:53:@19390.4]
  assign valid_60_20 = io_inValid_20 & _T_40814; // @[Switch.scala 30:36:@19391.4]
  assign _T_40817 = io_inAddr_21 == 6'h3c; // @[Switch.scala 30:53:@19393.4]
  assign valid_60_21 = io_inValid_21 & _T_40817; // @[Switch.scala 30:36:@19394.4]
  assign _T_40820 = io_inAddr_22 == 6'h3c; // @[Switch.scala 30:53:@19396.4]
  assign valid_60_22 = io_inValid_22 & _T_40820; // @[Switch.scala 30:36:@19397.4]
  assign _T_40823 = io_inAddr_23 == 6'h3c; // @[Switch.scala 30:53:@19399.4]
  assign valid_60_23 = io_inValid_23 & _T_40823; // @[Switch.scala 30:36:@19400.4]
  assign _T_40826 = io_inAddr_24 == 6'h3c; // @[Switch.scala 30:53:@19402.4]
  assign valid_60_24 = io_inValid_24 & _T_40826; // @[Switch.scala 30:36:@19403.4]
  assign _T_40829 = io_inAddr_25 == 6'h3c; // @[Switch.scala 30:53:@19405.4]
  assign valid_60_25 = io_inValid_25 & _T_40829; // @[Switch.scala 30:36:@19406.4]
  assign _T_40832 = io_inAddr_26 == 6'h3c; // @[Switch.scala 30:53:@19408.4]
  assign valid_60_26 = io_inValid_26 & _T_40832; // @[Switch.scala 30:36:@19409.4]
  assign _T_40835 = io_inAddr_27 == 6'h3c; // @[Switch.scala 30:53:@19411.4]
  assign valid_60_27 = io_inValid_27 & _T_40835; // @[Switch.scala 30:36:@19412.4]
  assign _T_40838 = io_inAddr_28 == 6'h3c; // @[Switch.scala 30:53:@19414.4]
  assign valid_60_28 = io_inValid_28 & _T_40838; // @[Switch.scala 30:36:@19415.4]
  assign _T_40841 = io_inAddr_29 == 6'h3c; // @[Switch.scala 30:53:@19417.4]
  assign valid_60_29 = io_inValid_29 & _T_40841; // @[Switch.scala 30:36:@19418.4]
  assign _T_40844 = io_inAddr_30 == 6'h3c; // @[Switch.scala 30:53:@19420.4]
  assign valid_60_30 = io_inValid_30 & _T_40844; // @[Switch.scala 30:36:@19421.4]
  assign _T_40847 = io_inAddr_31 == 6'h3c; // @[Switch.scala 30:53:@19423.4]
  assign valid_60_31 = io_inValid_31 & _T_40847; // @[Switch.scala 30:36:@19424.4]
  assign _T_40850 = io_inAddr_32 == 6'h3c; // @[Switch.scala 30:53:@19426.4]
  assign valid_60_32 = io_inValid_32 & _T_40850; // @[Switch.scala 30:36:@19427.4]
  assign _T_40853 = io_inAddr_33 == 6'h3c; // @[Switch.scala 30:53:@19429.4]
  assign valid_60_33 = io_inValid_33 & _T_40853; // @[Switch.scala 30:36:@19430.4]
  assign _T_40856 = io_inAddr_34 == 6'h3c; // @[Switch.scala 30:53:@19432.4]
  assign valid_60_34 = io_inValid_34 & _T_40856; // @[Switch.scala 30:36:@19433.4]
  assign _T_40859 = io_inAddr_35 == 6'h3c; // @[Switch.scala 30:53:@19435.4]
  assign valid_60_35 = io_inValid_35 & _T_40859; // @[Switch.scala 30:36:@19436.4]
  assign _T_40862 = io_inAddr_36 == 6'h3c; // @[Switch.scala 30:53:@19438.4]
  assign valid_60_36 = io_inValid_36 & _T_40862; // @[Switch.scala 30:36:@19439.4]
  assign _T_40865 = io_inAddr_37 == 6'h3c; // @[Switch.scala 30:53:@19441.4]
  assign valid_60_37 = io_inValid_37 & _T_40865; // @[Switch.scala 30:36:@19442.4]
  assign _T_40868 = io_inAddr_38 == 6'h3c; // @[Switch.scala 30:53:@19444.4]
  assign valid_60_38 = io_inValid_38 & _T_40868; // @[Switch.scala 30:36:@19445.4]
  assign _T_40871 = io_inAddr_39 == 6'h3c; // @[Switch.scala 30:53:@19447.4]
  assign valid_60_39 = io_inValid_39 & _T_40871; // @[Switch.scala 30:36:@19448.4]
  assign _T_40874 = io_inAddr_40 == 6'h3c; // @[Switch.scala 30:53:@19450.4]
  assign valid_60_40 = io_inValid_40 & _T_40874; // @[Switch.scala 30:36:@19451.4]
  assign _T_40877 = io_inAddr_41 == 6'h3c; // @[Switch.scala 30:53:@19453.4]
  assign valid_60_41 = io_inValid_41 & _T_40877; // @[Switch.scala 30:36:@19454.4]
  assign _T_40880 = io_inAddr_42 == 6'h3c; // @[Switch.scala 30:53:@19456.4]
  assign valid_60_42 = io_inValid_42 & _T_40880; // @[Switch.scala 30:36:@19457.4]
  assign _T_40883 = io_inAddr_43 == 6'h3c; // @[Switch.scala 30:53:@19459.4]
  assign valid_60_43 = io_inValid_43 & _T_40883; // @[Switch.scala 30:36:@19460.4]
  assign _T_40886 = io_inAddr_44 == 6'h3c; // @[Switch.scala 30:53:@19462.4]
  assign valid_60_44 = io_inValid_44 & _T_40886; // @[Switch.scala 30:36:@19463.4]
  assign _T_40889 = io_inAddr_45 == 6'h3c; // @[Switch.scala 30:53:@19465.4]
  assign valid_60_45 = io_inValid_45 & _T_40889; // @[Switch.scala 30:36:@19466.4]
  assign _T_40892 = io_inAddr_46 == 6'h3c; // @[Switch.scala 30:53:@19468.4]
  assign valid_60_46 = io_inValid_46 & _T_40892; // @[Switch.scala 30:36:@19469.4]
  assign _T_40895 = io_inAddr_47 == 6'h3c; // @[Switch.scala 30:53:@19471.4]
  assign valid_60_47 = io_inValid_47 & _T_40895; // @[Switch.scala 30:36:@19472.4]
  assign _T_40898 = io_inAddr_48 == 6'h3c; // @[Switch.scala 30:53:@19474.4]
  assign valid_60_48 = io_inValid_48 & _T_40898; // @[Switch.scala 30:36:@19475.4]
  assign _T_40901 = io_inAddr_49 == 6'h3c; // @[Switch.scala 30:53:@19477.4]
  assign valid_60_49 = io_inValid_49 & _T_40901; // @[Switch.scala 30:36:@19478.4]
  assign _T_40904 = io_inAddr_50 == 6'h3c; // @[Switch.scala 30:53:@19480.4]
  assign valid_60_50 = io_inValid_50 & _T_40904; // @[Switch.scala 30:36:@19481.4]
  assign _T_40907 = io_inAddr_51 == 6'h3c; // @[Switch.scala 30:53:@19483.4]
  assign valid_60_51 = io_inValid_51 & _T_40907; // @[Switch.scala 30:36:@19484.4]
  assign _T_40910 = io_inAddr_52 == 6'h3c; // @[Switch.scala 30:53:@19486.4]
  assign valid_60_52 = io_inValid_52 & _T_40910; // @[Switch.scala 30:36:@19487.4]
  assign _T_40913 = io_inAddr_53 == 6'h3c; // @[Switch.scala 30:53:@19489.4]
  assign valid_60_53 = io_inValid_53 & _T_40913; // @[Switch.scala 30:36:@19490.4]
  assign _T_40916 = io_inAddr_54 == 6'h3c; // @[Switch.scala 30:53:@19492.4]
  assign valid_60_54 = io_inValid_54 & _T_40916; // @[Switch.scala 30:36:@19493.4]
  assign _T_40919 = io_inAddr_55 == 6'h3c; // @[Switch.scala 30:53:@19495.4]
  assign valid_60_55 = io_inValid_55 & _T_40919; // @[Switch.scala 30:36:@19496.4]
  assign _T_40922 = io_inAddr_56 == 6'h3c; // @[Switch.scala 30:53:@19498.4]
  assign valid_60_56 = io_inValid_56 & _T_40922; // @[Switch.scala 30:36:@19499.4]
  assign _T_40925 = io_inAddr_57 == 6'h3c; // @[Switch.scala 30:53:@19501.4]
  assign valid_60_57 = io_inValid_57 & _T_40925; // @[Switch.scala 30:36:@19502.4]
  assign _T_40928 = io_inAddr_58 == 6'h3c; // @[Switch.scala 30:53:@19504.4]
  assign valid_60_58 = io_inValid_58 & _T_40928; // @[Switch.scala 30:36:@19505.4]
  assign _T_40931 = io_inAddr_59 == 6'h3c; // @[Switch.scala 30:53:@19507.4]
  assign valid_60_59 = io_inValid_59 & _T_40931; // @[Switch.scala 30:36:@19508.4]
  assign _T_40934 = io_inAddr_60 == 6'h3c; // @[Switch.scala 30:53:@19510.4]
  assign valid_60_60 = io_inValid_60 & _T_40934; // @[Switch.scala 30:36:@19511.4]
  assign _T_40937 = io_inAddr_61 == 6'h3c; // @[Switch.scala 30:53:@19513.4]
  assign valid_60_61 = io_inValid_61 & _T_40937; // @[Switch.scala 30:36:@19514.4]
  assign _T_40940 = io_inAddr_62 == 6'h3c; // @[Switch.scala 30:53:@19516.4]
  assign valid_60_62 = io_inValid_62 & _T_40940; // @[Switch.scala 30:36:@19517.4]
  assign _T_40943 = io_inAddr_63 == 6'h3c; // @[Switch.scala 30:53:@19519.4]
  assign valid_60_63 = io_inValid_63 & _T_40943; // @[Switch.scala 30:36:@19520.4]
  assign _T_41009 = valid_60_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@19522.4]
  assign _T_41010 = valid_60_61 ? 6'h3d : _T_41009; // @[Mux.scala 31:69:@19523.4]
  assign _T_41011 = valid_60_60 ? 6'h3c : _T_41010; // @[Mux.scala 31:69:@19524.4]
  assign _T_41012 = valid_60_59 ? 6'h3b : _T_41011; // @[Mux.scala 31:69:@19525.4]
  assign _T_41013 = valid_60_58 ? 6'h3a : _T_41012; // @[Mux.scala 31:69:@19526.4]
  assign _T_41014 = valid_60_57 ? 6'h39 : _T_41013; // @[Mux.scala 31:69:@19527.4]
  assign _T_41015 = valid_60_56 ? 6'h38 : _T_41014; // @[Mux.scala 31:69:@19528.4]
  assign _T_41016 = valid_60_55 ? 6'h37 : _T_41015; // @[Mux.scala 31:69:@19529.4]
  assign _T_41017 = valid_60_54 ? 6'h36 : _T_41016; // @[Mux.scala 31:69:@19530.4]
  assign _T_41018 = valid_60_53 ? 6'h35 : _T_41017; // @[Mux.scala 31:69:@19531.4]
  assign _T_41019 = valid_60_52 ? 6'h34 : _T_41018; // @[Mux.scala 31:69:@19532.4]
  assign _T_41020 = valid_60_51 ? 6'h33 : _T_41019; // @[Mux.scala 31:69:@19533.4]
  assign _T_41021 = valid_60_50 ? 6'h32 : _T_41020; // @[Mux.scala 31:69:@19534.4]
  assign _T_41022 = valid_60_49 ? 6'h31 : _T_41021; // @[Mux.scala 31:69:@19535.4]
  assign _T_41023 = valid_60_48 ? 6'h30 : _T_41022; // @[Mux.scala 31:69:@19536.4]
  assign _T_41024 = valid_60_47 ? 6'h2f : _T_41023; // @[Mux.scala 31:69:@19537.4]
  assign _T_41025 = valid_60_46 ? 6'h2e : _T_41024; // @[Mux.scala 31:69:@19538.4]
  assign _T_41026 = valid_60_45 ? 6'h2d : _T_41025; // @[Mux.scala 31:69:@19539.4]
  assign _T_41027 = valid_60_44 ? 6'h2c : _T_41026; // @[Mux.scala 31:69:@19540.4]
  assign _T_41028 = valid_60_43 ? 6'h2b : _T_41027; // @[Mux.scala 31:69:@19541.4]
  assign _T_41029 = valid_60_42 ? 6'h2a : _T_41028; // @[Mux.scala 31:69:@19542.4]
  assign _T_41030 = valid_60_41 ? 6'h29 : _T_41029; // @[Mux.scala 31:69:@19543.4]
  assign _T_41031 = valid_60_40 ? 6'h28 : _T_41030; // @[Mux.scala 31:69:@19544.4]
  assign _T_41032 = valid_60_39 ? 6'h27 : _T_41031; // @[Mux.scala 31:69:@19545.4]
  assign _T_41033 = valid_60_38 ? 6'h26 : _T_41032; // @[Mux.scala 31:69:@19546.4]
  assign _T_41034 = valid_60_37 ? 6'h25 : _T_41033; // @[Mux.scala 31:69:@19547.4]
  assign _T_41035 = valid_60_36 ? 6'h24 : _T_41034; // @[Mux.scala 31:69:@19548.4]
  assign _T_41036 = valid_60_35 ? 6'h23 : _T_41035; // @[Mux.scala 31:69:@19549.4]
  assign _T_41037 = valid_60_34 ? 6'h22 : _T_41036; // @[Mux.scala 31:69:@19550.4]
  assign _T_41038 = valid_60_33 ? 6'h21 : _T_41037; // @[Mux.scala 31:69:@19551.4]
  assign _T_41039 = valid_60_32 ? 6'h20 : _T_41038; // @[Mux.scala 31:69:@19552.4]
  assign _T_41040 = valid_60_31 ? 6'h1f : _T_41039; // @[Mux.scala 31:69:@19553.4]
  assign _T_41041 = valid_60_30 ? 6'h1e : _T_41040; // @[Mux.scala 31:69:@19554.4]
  assign _T_41042 = valid_60_29 ? 6'h1d : _T_41041; // @[Mux.scala 31:69:@19555.4]
  assign _T_41043 = valid_60_28 ? 6'h1c : _T_41042; // @[Mux.scala 31:69:@19556.4]
  assign _T_41044 = valid_60_27 ? 6'h1b : _T_41043; // @[Mux.scala 31:69:@19557.4]
  assign _T_41045 = valid_60_26 ? 6'h1a : _T_41044; // @[Mux.scala 31:69:@19558.4]
  assign _T_41046 = valid_60_25 ? 6'h19 : _T_41045; // @[Mux.scala 31:69:@19559.4]
  assign _T_41047 = valid_60_24 ? 6'h18 : _T_41046; // @[Mux.scala 31:69:@19560.4]
  assign _T_41048 = valid_60_23 ? 6'h17 : _T_41047; // @[Mux.scala 31:69:@19561.4]
  assign _T_41049 = valid_60_22 ? 6'h16 : _T_41048; // @[Mux.scala 31:69:@19562.4]
  assign _T_41050 = valid_60_21 ? 6'h15 : _T_41049; // @[Mux.scala 31:69:@19563.4]
  assign _T_41051 = valid_60_20 ? 6'h14 : _T_41050; // @[Mux.scala 31:69:@19564.4]
  assign _T_41052 = valid_60_19 ? 6'h13 : _T_41051; // @[Mux.scala 31:69:@19565.4]
  assign _T_41053 = valid_60_18 ? 6'h12 : _T_41052; // @[Mux.scala 31:69:@19566.4]
  assign _T_41054 = valid_60_17 ? 6'h11 : _T_41053; // @[Mux.scala 31:69:@19567.4]
  assign _T_41055 = valid_60_16 ? 6'h10 : _T_41054; // @[Mux.scala 31:69:@19568.4]
  assign _T_41056 = valid_60_15 ? 6'hf : _T_41055; // @[Mux.scala 31:69:@19569.4]
  assign _T_41057 = valid_60_14 ? 6'he : _T_41056; // @[Mux.scala 31:69:@19570.4]
  assign _T_41058 = valid_60_13 ? 6'hd : _T_41057; // @[Mux.scala 31:69:@19571.4]
  assign _T_41059 = valid_60_12 ? 6'hc : _T_41058; // @[Mux.scala 31:69:@19572.4]
  assign _T_41060 = valid_60_11 ? 6'hb : _T_41059; // @[Mux.scala 31:69:@19573.4]
  assign _T_41061 = valid_60_10 ? 6'ha : _T_41060; // @[Mux.scala 31:69:@19574.4]
  assign _T_41062 = valid_60_9 ? 6'h9 : _T_41061; // @[Mux.scala 31:69:@19575.4]
  assign _T_41063 = valid_60_8 ? 6'h8 : _T_41062; // @[Mux.scala 31:69:@19576.4]
  assign _T_41064 = valid_60_7 ? 6'h7 : _T_41063; // @[Mux.scala 31:69:@19577.4]
  assign _T_41065 = valid_60_6 ? 6'h6 : _T_41064; // @[Mux.scala 31:69:@19578.4]
  assign _T_41066 = valid_60_5 ? 6'h5 : _T_41065; // @[Mux.scala 31:69:@19579.4]
  assign _T_41067 = valid_60_4 ? 6'h4 : _T_41066; // @[Mux.scala 31:69:@19580.4]
  assign _T_41068 = valid_60_3 ? 6'h3 : _T_41067; // @[Mux.scala 31:69:@19581.4]
  assign _T_41069 = valid_60_2 ? 6'h2 : _T_41068; // @[Mux.scala 31:69:@19582.4]
  assign _T_41070 = valid_60_1 ? 6'h1 : _T_41069; // @[Mux.scala 31:69:@19583.4]
  assign select_60 = valid_60_0 ? 6'h0 : _T_41070; // @[Mux.scala 31:69:@19584.4]
  assign _GEN_3841 = 6'h1 == select_60 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3842 = 6'h2 == select_60 ? io_inData_2 : _GEN_3841; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3843 = 6'h3 == select_60 ? io_inData_3 : _GEN_3842; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3844 = 6'h4 == select_60 ? io_inData_4 : _GEN_3843; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3845 = 6'h5 == select_60 ? io_inData_5 : _GEN_3844; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3846 = 6'h6 == select_60 ? io_inData_6 : _GEN_3845; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3847 = 6'h7 == select_60 ? io_inData_7 : _GEN_3846; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3848 = 6'h8 == select_60 ? io_inData_8 : _GEN_3847; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3849 = 6'h9 == select_60 ? io_inData_9 : _GEN_3848; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3850 = 6'ha == select_60 ? io_inData_10 : _GEN_3849; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3851 = 6'hb == select_60 ? io_inData_11 : _GEN_3850; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3852 = 6'hc == select_60 ? io_inData_12 : _GEN_3851; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3853 = 6'hd == select_60 ? io_inData_13 : _GEN_3852; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3854 = 6'he == select_60 ? io_inData_14 : _GEN_3853; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3855 = 6'hf == select_60 ? io_inData_15 : _GEN_3854; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3856 = 6'h10 == select_60 ? io_inData_16 : _GEN_3855; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3857 = 6'h11 == select_60 ? io_inData_17 : _GEN_3856; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3858 = 6'h12 == select_60 ? io_inData_18 : _GEN_3857; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3859 = 6'h13 == select_60 ? io_inData_19 : _GEN_3858; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3860 = 6'h14 == select_60 ? io_inData_20 : _GEN_3859; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3861 = 6'h15 == select_60 ? io_inData_21 : _GEN_3860; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3862 = 6'h16 == select_60 ? io_inData_22 : _GEN_3861; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3863 = 6'h17 == select_60 ? io_inData_23 : _GEN_3862; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3864 = 6'h18 == select_60 ? io_inData_24 : _GEN_3863; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3865 = 6'h19 == select_60 ? io_inData_25 : _GEN_3864; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3866 = 6'h1a == select_60 ? io_inData_26 : _GEN_3865; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3867 = 6'h1b == select_60 ? io_inData_27 : _GEN_3866; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3868 = 6'h1c == select_60 ? io_inData_28 : _GEN_3867; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3869 = 6'h1d == select_60 ? io_inData_29 : _GEN_3868; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3870 = 6'h1e == select_60 ? io_inData_30 : _GEN_3869; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3871 = 6'h1f == select_60 ? io_inData_31 : _GEN_3870; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3872 = 6'h20 == select_60 ? io_inData_32 : _GEN_3871; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3873 = 6'h21 == select_60 ? io_inData_33 : _GEN_3872; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3874 = 6'h22 == select_60 ? io_inData_34 : _GEN_3873; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3875 = 6'h23 == select_60 ? io_inData_35 : _GEN_3874; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3876 = 6'h24 == select_60 ? io_inData_36 : _GEN_3875; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3877 = 6'h25 == select_60 ? io_inData_37 : _GEN_3876; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3878 = 6'h26 == select_60 ? io_inData_38 : _GEN_3877; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3879 = 6'h27 == select_60 ? io_inData_39 : _GEN_3878; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3880 = 6'h28 == select_60 ? io_inData_40 : _GEN_3879; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3881 = 6'h29 == select_60 ? io_inData_41 : _GEN_3880; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3882 = 6'h2a == select_60 ? io_inData_42 : _GEN_3881; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3883 = 6'h2b == select_60 ? io_inData_43 : _GEN_3882; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3884 = 6'h2c == select_60 ? io_inData_44 : _GEN_3883; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3885 = 6'h2d == select_60 ? io_inData_45 : _GEN_3884; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3886 = 6'h2e == select_60 ? io_inData_46 : _GEN_3885; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3887 = 6'h2f == select_60 ? io_inData_47 : _GEN_3886; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3888 = 6'h30 == select_60 ? io_inData_48 : _GEN_3887; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3889 = 6'h31 == select_60 ? io_inData_49 : _GEN_3888; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3890 = 6'h32 == select_60 ? io_inData_50 : _GEN_3889; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3891 = 6'h33 == select_60 ? io_inData_51 : _GEN_3890; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3892 = 6'h34 == select_60 ? io_inData_52 : _GEN_3891; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3893 = 6'h35 == select_60 ? io_inData_53 : _GEN_3892; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3894 = 6'h36 == select_60 ? io_inData_54 : _GEN_3893; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3895 = 6'h37 == select_60 ? io_inData_55 : _GEN_3894; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3896 = 6'h38 == select_60 ? io_inData_56 : _GEN_3895; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3897 = 6'h39 == select_60 ? io_inData_57 : _GEN_3896; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3898 = 6'h3a == select_60 ? io_inData_58 : _GEN_3897; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3899 = 6'h3b == select_60 ? io_inData_59 : _GEN_3898; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3900 = 6'h3c == select_60 ? io_inData_60 : _GEN_3899; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3901 = 6'h3d == select_60 ? io_inData_61 : _GEN_3900; // @[Switch.scala 33:19:@19586.4]
  assign _GEN_3902 = 6'h3e == select_60 ? io_inData_62 : _GEN_3901; // @[Switch.scala 33:19:@19586.4]
  assign _T_41079 = {valid_60_7,valid_60_6,valid_60_5,valid_60_4,valid_60_3,valid_60_2,valid_60_1,valid_60_0}; // @[Switch.scala 34:32:@19593.4]
  assign _T_41087 = {valid_60_15,valid_60_14,valid_60_13,valid_60_12,valid_60_11,valid_60_10,valid_60_9,valid_60_8,_T_41079}; // @[Switch.scala 34:32:@19601.4]
  assign _T_41094 = {valid_60_23,valid_60_22,valid_60_21,valid_60_20,valid_60_19,valid_60_18,valid_60_17,valid_60_16}; // @[Switch.scala 34:32:@19608.4]
  assign _T_41103 = {valid_60_31,valid_60_30,valid_60_29,valid_60_28,valid_60_27,valid_60_26,valid_60_25,valid_60_24,_T_41094,_T_41087}; // @[Switch.scala 34:32:@19617.4]
  assign _T_41110 = {valid_60_39,valid_60_38,valid_60_37,valid_60_36,valid_60_35,valid_60_34,valid_60_33,valid_60_32}; // @[Switch.scala 34:32:@19624.4]
  assign _T_41118 = {valid_60_47,valid_60_46,valid_60_45,valid_60_44,valid_60_43,valid_60_42,valid_60_41,valid_60_40,_T_41110}; // @[Switch.scala 34:32:@19632.4]
  assign _T_41125 = {valid_60_55,valid_60_54,valid_60_53,valid_60_52,valid_60_51,valid_60_50,valid_60_49,valid_60_48}; // @[Switch.scala 34:32:@19639.4]
  assign _T_41134 = {valid_60_63,valid_60_62,valid_60_61,valid_60_60,valid_60_59,valid_60_58,valid_60_57,valid_60_56,_T_41125,_T_41118}; // @[Switch.scala 34:32:@19648.4]
  assign _T_41135 = {_T_41134,_T_41103}; // @[Switch.scala 34:32:@19649.4]
  assign _T_41139 = io_inAddr_0 == 6'h3d; // @[Switch.scala 30:53:@19652.4]
  assign valid_61_0 = io_inValid_0 & _T_41139; // @[Switch.scala 30:36:@19653.4]
  assign _T_41142 = io_inAddr_1 == 6'h3d; // @[Switch.scala 30:53:@19655.4]
  assign valid_61_1 = io_inValid_1 & _T_41142; // @[Switch.scala 30:36:@19656.4]
  assign _T_41145 = io_inAddr_2 == 6'h3d; // @[Switch.scala 30:53:@19658.4]
  assign valid_61_2 = io_inValid_2 & _T_41145; // @[Switch.scala 30:36:@19659.4]
  assign _T_41148 = io_inAddr_3 == 6'h3d; // @[Switch.scala 30:53:@19661.4]
  assign valid_61_3 = io_inValid_3 & _T_41148; // @[Switch.scala 30:36:@19662.4]
  assign _T_41151 = io_inAddr_4 == 6'h3d; // @[Switch.scala 30:53:@19664.4]
  assign valid_61_4 = io_inValid_4 & _T_41151; // @[Switch.scala 30:36:@19665.4]
  assign _T_41154 = io_inAddr_5 == 6'h3d; // @[Switch.scala 30:53:@19667.4]
  assign valid_61_5 = io_inValid_5 & _T_41154; // @[Switch.scala 30:36:@19668.4]
  assign _T_41157 = io_inAddr_6 == 6'h3d; // @[Switch.scala 30:53:@19670.4]
  assign valid_61_6 = io_inValid_6 & _T_41157; // @[Switch.scala 30:36:@19671.4]
  assign _T_41160 = io_inAddr_7 == 6'h3d; // @[Switch.scala 30:53:@19673.4]
  assign valid_61_7 = io_inValid_7 & _T_41160; // @[Switch.scala 30:36:@19674.4]
  assign _T_41163 = io_inAddr_8 == 6'h3d; // @[Switch.scala 30:53:@19676.4]
  assign valid_61_8 = io_inValid_8 & _T_41163; // @[Switch.scala 30:36:@19677.4]
  assign _T_41166 = io_inAddr_9 == 6'h3d; // @[Switch.scala 30:53:@19679.4]
  assign valid_61_9 = io_inValid_9 & _T_41166; // @[Switch.scala 30:36:@19680.4]
  assign _T_41169 = io_inAddr_10 == 6'h3d; // @[Switch.scala 30:53:@19682.4]
  assign valid_61_10 = io_inValid_10 & _T_41169; // @[Switch.scala 30:36:@19683.4]
  assign _T_41172 = io_inAddr_11 == 6'h3d; // @[Switch.scala 30:53:@19685.4]
  assign valid_61_11 = io_inValid_11 & _T_41172; // @[Switch.scala 30:36:@19686.4]
  assign _T_41175 = io_inAddr_12 == 6'h3d; // @[Switch.scala 30:53:@19688.4]
  assign valid_61_12 = io_inValid_12 & _T_41175; // @[Switch.scala 30:36:@19689.4]
  assign _T_41178 = io_inAddr_13 == 6'h3d; // @[Switch.scala 30:53:@19691.4]
  assign valid_61_13 = io_inValid_13 & _T_41178; // @[Switch.scala 30:36:@19692.4]
  assign _T_41181 = io_inAddr_14 == 6'h3d; // @[Switch.scala 30:53:@19694.4]
  assign valid_61_14 = io_inValid_14 & _T_41181; // @[Switch.scala 30:36:@19695.4]
  assign _T_41184 = io_inAddr_15 == 6'h3d; // @[Switch.scala 30:53:@19697.4]
  assign valid_61_15 = io_inValid_15 & _T_41184; // @[Switch.scala 30:36:@19698.4]
  assign _T_41187 = io_inAddr_16 == 6'h3d; // @[Switch.scala 30:53:@19700.4]
  assign valid_61_16 = io_inValid_16 & _T_41187; // @[Switch.scala 30:36:@19701.4]
  assign _T_41190 = io_inAddr_17 == 6'h3d; // @[Switch.scala 30:53:@19703.4]
  assign valid_61_17 = io_inValid_17 & _T_41190; // @[Switch.scala 30:36:@19704.4]
  assign _T_41193 = io_inAddr_18 == 6'h3d; // @[Switch.scala 30:53:@19706.4]
  assign valid_61_18 = io_inValid_18 & _T_41193; // @[Switch.scala 30:36:@19707.4]
  assign _T_41196 = io_inAddr_19 == 6'h3d; // @[Switch.scala 30:53:@19709.4]
  assign valid_61_19 = io_inValid_19 & _T_41196; // @[Switch.scala 30:36:@19710.4]
  assign _T_41199 = io_inAddr_20 == 6'h3d; // @[Switch.scala 30:53:@19712.4]
  assign valid_61_20 = io_inValid_20 & _T_41199; // @[Switch.scala 30:36:@19713.4]
  assign _T_41202 = io_inAddr_21 == 6'h3d; // @[Switch.scala 30:53:@19715.4]
  assign valid_61_21 = io_inValid_21 & _T_41202; // @[Switch.scala 30:36:@19716.4]
  assign _T_41205 = io_inAddr_22 == 6'h3d; // @[Switch.scala 30:53:@19718.4]
  assign valid_61_22 = io_inValid_22 & _T_41205; // @[Switch.scala 30:36:@19719.4]
  assign _T_41208 = io_inAddr_23 == 6'h3d; // @[Switch.scala 30:53:@19721.4]
  assign valid_61_23 = io_inValid_23 & _T_41208; // @[Switch.scala 30:36:@19722.4]
  assign _T_41211 = io_inAddr_24 == 6'h3d; // @[Switch.scala 30:53:@19724.4]
  assign valid_61_24 = io_inValid_24 & _T_41211; // @[Switch.scala 30:36:@19725.4]
  assign _T_41214 = io_inAddr_25 == 6'h3d; // @[Switch.scala 30:53:@19727.4]
  assign valid_61_25 = io_inValid_25 & _T_41214; // @[Switch.scala 30:36:@19728.4]
  assign _T_41217 = io_inAddr_26 == 6'h3d; // @[Switch.scala 30:53:@19730.4]
  assign valid_61_26 = io_inValid_26 & _T_41217; // @[Switch.scala 30:36:@19731.4]
  assign _T_41220 = io_inAddr_27 == 6'h3d; // @[Switch.scala 30:53:@19733.4]
  assign valid_61_27 = io_inValid_27 & _T_41220; // @[Switch.scala 30:36:@19734.4]
  assign _T_41223 = io_inAddr_28 == 6'h3d; // @[Switch.scala 30:53:@19736.4]
  assign valid_61_28 = io_inValid_28 & _T_41223; // @[Switch.scala 30:36:@19737.4]
  assign _T_41226 = io_inAddr_29 == 6'h3d; // @[Switch.scala 30:53:@19739.4]
  assign valid_61_29 = io_inValid_29 & _T_41226; // @[Switch.scala 30:36:@19740.4]
  assign _T_41229 = io_inAddr_30 == 6'h3d; // @[Switch.scala 30:53:@19742.4]
  assign valid_61_30 = io_inValid_30 & _T_41229; // @[Switch.scala 30:36:@19743.4]
  assign _T_41232 = io_inAddr_31 == 6'h3d; // @[Switch.scala 30:53:@19745.4]
  assign valid_61_31 = io_inValid_31 & _T_41232; // @[Switch.scala 30:36:@19746.4]
  assign _T_41235 = io_inAddr_32 == 6'h3d; // @[Switch.scala 30:53:@19748.4]
  assign valid_61_32 = io_inValid_32 & _T_41235; // @[Switch.scala 30:36:@19749.4]
  assign _T_41238 = io_inAddr_33 == 6'h3d; // @[Switch.scala 30:53:@19751.4]
  assign valid_61_33 = io_inValid_33 & _T_41238; // @[Switch.scala 30:36:@19752.4]
  assign _T_41241 = io_inAddr_34 == 6'h3d; // @[Switch.scala 30:53:@19754.4]
  assign valid_61_34 = io_inValid_34 & _T_41241; // @[Switch.scala 30:36:@19755.4]
  assign _T_41244 = io_inAddr_35 == 6'h3d; // @[Switch.scala 30:53:@19757.4]
  assign valid_61_35 = io_inValid_35 & _T_41244; // @[Switch.scala 30:36:@19758.4]
  assign _T_41247 = io_inAddr_36 == 6'h3d; // @[Switch.scala 30:53:@19760.4]
  assign valid_61_36 = io_inValid_36 & _T_41247; // @[Switch.scala 30:36:@19761.4]
  assign _T_41250 = io_inAddr_37 == 6'h3d; // @[Switch.scala 30:53:@19763.4]
  assign valid_61_37 = io_inValid_37 & _T_41250; // @[Switch.scala 30:36:@19764.4]
  assign _T_41253 = io_inAddr_38 == 6'h3d; // @[Switch.scala 30:53:@19766.4]
  assign valid_61_38 = io_inValid_38 & _T_41253; // @[Switch.scala 30:36:@19767.4]
  assign _T_41256 = io_inAddr_39 == 6'h3d; // @[Switch.scala 30:53:@19769.4]
  assign valid_61_39 = io_inValid_39 & _T_41256; // @[Switch.scala 30:36:@19770.4]
  assign _T_41259 = io_inAddr_40 == 6'h3d; // @[Switch.scala 30:53:@19772.4]
  assign valid_61_40 = io_inValid_40 & _T_41259; // @[Switch.scala 30:36:@19773.4]
  assign _T_41262 = io_inAddr_41 == 6'h3d; // @[Switch.scala 30:53:@19775.4]
  assign valid_61_41 = io_inValid_41 & _T_41262; // @[Switch.scala 30:36:@19776.4]
  assign _T_41265 = io_inAddr_42 == 6'h3d; // @[Switch.scala 30:53:@19778.4]
  assign valid_61_42 = io_inValid_42 & _T_41265; // @[Switch.scala 30:36:@19779.4]
  assign _T_41268 = io_inAddr_43 == 6'h3d; // @[Switch.scala 30:53:@19781.4]
  assign valid_61_43 = io_inValid_43 & _T_41268; // @[Switch.scala 30:36:@19782.4]
  assign _T_41271 = io_inAddr_44 == 6'h3d; // @[Switch.scala 30:53:@19784.4]
  assign valid_61_44 = io_inValid_44 & _T_41271; // @[Switch.scala 30:36:@19785.4]
  assign _T_41274 = io_inAddr_45 == 6'h3d; // @[Switch.scala 30:53:@19787.4]
  assign valid_61_45 = io_inValid_45 & _T_41274; // @[Switch.scala 30:36:@19788.4]
  assign _T_41277 = io_inAddr_46 == 6'h3d; // @[Switch.scala 30:53:@19790.4]
  assign valid_61_46 = io_inValid_46 & _T_41277; // @[Switch.scala 30:36:@19791.4]
  assign _T_41280 = io_inAddr_47 == 6'h3d; // @[Switch.scala 30:53:@19793.4]
  assign valid_61_47 = io_inValid_47 & _T_41280; // @[Switch.scala 30:36:@19794.4]
  assign _T_41283 = io_inAddr_48 == 6'h3d; // @[Switch.scala 30:53:@19796.4]
  assign valid_61_48 = io_inValid_48 & _T_41283; // @[Switch.scala 30:36:@19797.4]
  assign _T_41286 = io_inAddr_49 == 6'h3d; // @[Switch.scala 30:53:@19799.4]
  assign valid_61_49 = io_inValid_49 & _T_41286; // @[Switch.scala 30:36:@19800.4]
  assign _T_41289 = io_inAddr_50 == 6'h3d; // @[Switch.scala 30:53:@19802.4]
  assign valid_61_50 = io_inValid_50 & _T_41289; // @[Switch.scala 30:36:@19803.4]
  assign _T_41292 = io_inAddr_51 == 6'h3d; // @[Switch.scala 30:53:@19805.4]
  assign valid_61_51 = io_inValid_51 & _T_41292; // @[Switch.scala 30:36:@19806.4]
  assign _T_41295 = io_inAddr_52 == 6'h3d; // @[Switch.scala 30:53:@19808.4]
  assign valid_61_52 = io_inValid_52 & _T_41295; // @[Switch.scala 30:36:@19809.4]
  assign _T_41298 = io_inAddr_53 == 6'h3d; // @[Switch.scala 30:53:@19811.4]
  assign valid_61_53 = io_inValid_53 & _T_41298; // @[Switch.scala 30:36:@19812.4]
  assign _T_41301 = io_inAddr_54 == 6'h3d; // @[Switch.scala 30:53:@19814.4]
  assign valid_61_54 = io_inValid_54 & _T_41301; // @[Switch.scala 30:36:@19815.4]
  assign _T_41304 = io_inAddr_55 == 6'h3d; // @[Switch.scala 30:53:@19817.4]
  assign valid_61_55 = io_inValid_55 & _T_41304; // @[Switch.scala 30:36:@19818.4]
  assign _T_41307 = io_inAddr_56 == 6'h3d; // @[Switch.scala 30:53:@19820.4]
  assign valid_61_56 = io_inValid_56 & _T_41307; // @[Switch.scala 30:36:@19821.4]
  assign _T_41310 = io_inAddr_57 == 6'h3d; // @[Switch.scala 30:53:@19823.4]
  assign valid_61_57 = io_inValid_57 & _T_41310; // @[Switch.scala 30:36:@19824.4]
  assign _T_41313 = io_inAddr_58 == 6'h3d; // @[Switch.scala 30:53:@19826.4]
  assign valid_61_58 = io_inValid_58 & _T_41313; // @[Switch.scala 30:36:@19827.4]
  assign _T_41316 = io_inAddr_59 == 6'h3d; // @[Switch.scala 30:53:@19829.4]
  assign valid_61_59 = io_inValid_59 & _T_41316; // @[Switch.scala 30:36:@19830.4]
  assign _T_41319 = io_inAddr_60 == 6'h3d; // @[Switch.scala 30:53:@19832.4]
  assign valid_61_60 = io_inValid_60 & _T_41319; // @[Switch.scala 30:36:@19833.4]
  assign _T_41322 = io_inAddr_61 == 6'h3d; // @[Switch.scala 30:53:@19835.4]
  assign valid_61_61 = io_inValid_61 & _T_41322; // @[Switch.scala 30:36:@19836.4]
  assign _T_41325 = io_inAddr_62 == 6'h3d; // @[Switch.scala 30:53:@19838.4]
  assign valid_61_62 = io_inValid_62 & _T_41325; // @[Switch.scala 30:36:@19839.4]
  assign _T_41328 = io_inAddr_63 == 6'h3d; // @[Switch.scala 30:53:@19841.4]
  assign valid_61_63 = io_inValid_63 & _T_41328; // @[Switch.scala 30:36:@19842.4]
  assign _T_41394 = valid_61_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@19844.4]
  assign _T_41395 = valid_61_61 ? 6'h3d : _T_41394; // @[Mux.scala 31:69:@19845.4]
  assign _T_41396 = valid_61_60 ? 6'h3c : _T_41395; // @[Mux.scala 31:69:@19846.4]
  assign _T_41397 = valid_61_59 ? 6'h3b : _T_41396; // @[Mux.scala 31:69:@19847.4]
  assign _T_41398 = valid_61_58 ? 6'h3a : _T_41397; // @[Mux.scala 31:69:@19848.4]
  assign _T_41399 = valid_61_57 ? 6'h39 : _T_41398; // @[Mux.scala 31:69:@19849.4]
  assign _T_41400 = valid_61_56 ? 6'h38 : _T_41399; // @[Mux.scala 31:69:@19850.4]
  assign _T_41401 = valid_61_55 ? 6'h37 : _T_41400; // @[Mux.scala 31:69:@19851.4]
  assign _T_41402 = valid_61_54 ? 6'h36 : _T_41401; // @[Mux.scala 31:69:@19852.4]
  assign _T_41403 = valid_61_53 ? 6'h35 : _T_41402; // @[Mux.scala 31:69:@19853.4]
  assign _T_41404 = valid_61_52 ? 6'h34 : _T_41403; // @[Mux.scala 31:69:@19854.4]
  assign _T_41405 = valid_61_51 ? 6'h33 : _T_41404; // @[Mux.scala 31:69:@19855.4]
  assign _T_41406 = valid_61_50 ? 6'h32 : _T_41405; // @[Mux.scala 31:69:@19856.4]
  assign _T_41407 = valid_61_49 ? 6'h31 : _T_41406; // @[Mux.scala 31:69:@19857.4]
  assign _T_41408 = valid_61_48 ? 6'h30 : _T_41407; // @[Mux.scala 31:69:@19858.4]
  assign _T_41409 = valid_61_47 ? 6'h2f : _T_41408; // @[Mux.scala 31:69:@19859.4]
  assign _T_41410 = valid_61_46 ? 6'h2e : _T_41409; // @[Mux.scala 31:69:@19860.4]
  assign _T_41411 = valid_61_45 ? 6'h2d : _T_41410; // @[Mux.scala 31:69:@19861.4]
  assign _T_41412 = valid_61_44 ? 6'h2c : _T_41411; // @[Mux.scala 31:69:@19862.4]
  assign _T_41413 = valid_61_43 ? 6'h2b : _T_41412; // @[Mux.scala 31:69:@19863.4]
  assign _T_41414 = valid_61_42 ? 6'h2a : _T_41413; // @[Mux.scala 31:69:@19864.4]
  assign _T_41415 = valid_61_41 ? 6'h29 : _T_41414; // @[Mux.scala 31:69:@19865.4]
  assign _T_41416 = valid_61_40 ? 6'h28 : _T_41415; // @[Mux.scala 31:69:@19866.4]
  assign _T_41417 = valid_61_39 ? 6'h27 : _T_41416; // @[Mux.scala 31:69:@19867.4]
  assign _T_41418 = valid_61_38 ? 6'h26 : _T_41417; // @[Mux.scala 31:69:@19868.4]
  assign _T_41419 = valid_61_37 ? 6'h25 : _T_41418; // @[Mux.scala 31:69:@19869.4]
  assign _T_41420 = valid_61_36 ? 6'h24 : _T_41419; // @[Mux.scala 31:69:@19870.4]
  assign _T_41421 = valid_61_35 ? 6'h23 : _T_41420; // @[Mux.scala 31:69:@19871.4]
  assign _T_41422 = valid_61_34 ? 6'h22 : _T_41421; // @[Mux.scala 31:69:@19872.4]
  assign _T_41423 = valid_61_33 ? 6'h21 : _T_41422; // @[Mux.scala 31:69:@19873.4]
  assign _T_41424 = valid_61_32 ? 6'h20 : _T_41423; // @[Mux.scala 31:69:@19874.4]
  assign _T_41425 = valid_61_31 ? 6'h1f : _T_41424; // @[Mux.scala 31:69:@19875.4]
  assign _T_41426 = valid_61_30 ? 6'h1e : _T_41425; // @[Mux.scala 31:69:@19876.4]
  assign _T_41427 = valid_61_29 ? 6'h1d : _T_41426; // @[Mux.scala 31:69:@19877.4]
  assign _T_41428 = valid_61_28 ? 6'h1c : _T_41427; // @[Mux.scala 31:69:@19878.4]
  assign _T_41429 = valid_61_27 ? 6'h1b : _T_41428; // @[Mux.scala 31:69:@19879.4]
  assign _T_41430 = valid_61_26 ? 6'h1a : _T_41429; // @[Mux.scala 31:69:@19880.4]
  assign _T_41431 = valid_61_25 ? 6'h19 : _T_41430; // @[Mux.scala 31:69:@19881.4]
  assign _T_41432 = valid_61_24 ? 6'h18 : _T_41431; // @[Mux.scala 31:69:@19882.4]
  assign _T_41433 = valid_61_23 ? 6'h17 : _T_41432; // @[Mux.scala 31:69:@19883.4]
  assign _T_41434 = valid_61_22 ? 6'h16 : _T_41433; // @[Mux.scala 31:69:@19884.4]
  assign _T_41435 = valid_61_21 ? 6'h15 : _T_41434; // @[Mux.scala 31:69:@19885.4]
  assign _T_41436 = valid_61_20 ? 6'h14 : _T_41435; // @[Mux.scala 31:69:@19886.4]
  assign _T_41437 = valid_61_19 ? 6'h13 : _T_41436; // @[Mux.scala 31:69:@19887.4]
  assign _T_41438 = valid_61_18 ? 6'h12 : _T_41437; // @[Mux.scala 31:69:@19888.4]
  assign _T_41439 = valid_61_17 ? 6'h11 : _T_41438; // @[Mux.scala 31:69:@19889.4]
  assign _T_41440 = valid_61_16 ? 6'h10 : _T_41439; // @[Mux.scala 31:69:@19890.4]
  assign _T_41441 = valid_61_15 ? 6'hf : _T_41440; // @[Mux.scala 31:69:@19891.4]
  assign _T_41442 = valid_61_14 ? 6'he : _T_41441; // @[Mux.scala 31:69:@19892.4]
  assign _T_41443 = valid_61_13 ? 6'hd : _T_41442; // @[Mux.scala 31:69:@19893.4]
  assign _T_41444 = valid_61_12 ? 6'hc : _T_41443; // @[Mux.scala 31:69:@19894.4]
  assign _T_41445 = valid_61_11 ? 6'hb : _T_41444; // @[Mux.scala 31:69:@19895.4]
  assign _T_41446 = valid_61_10 ? 6'ha : _T_41445; // @[Mux.scala 31:69:@19896.4]
  assign _T_41447 = valid_61_9 ? 6'h9 : _T_41446; // @[Mux.scala 31:69:@19897.4]
  assign _T_41448 = valid_61_8 ? 6'h8 : _T_41447; // @[Mux.scala 31:69:@19898.4]
  assign _T_41449 = valid_61_7 ? 6'h7 : _T_41448; // @[Mux.scala 31:69:@19899.4]
  assign _T_41450 = valid_61_6 ? 6'h6 : _T_41449; // @[Mux.scala 31:69:@19900.4]
  assign _T_41451 = valid_61_5 ? 6'h5 : _T_41450; // @[Mux.scala 31:69:@19901.4]
  assign _T_41452 = valid_61_4 ? 6'h4 : _T_41451; // @[Mux.scala 31:69:@19902.4]
  assign _T_41453 = valid_61_3 ? 6'h3 : _T_41452; // @[Mux.scala 31:69:@19903.4]
  assign _T_41454 = valid_61_2 ? 6'h2 : _T_41453; // @[Mux.scala 31:69:@19904.4]
  assign _T_41455 = valid_61_1 ? 6'h1 : _T_41454; // @[Mux.scala 31:69:@19905.4]
  assign select_61 = valid_61_0 ? 6'h0 : _T_41455; // @[Mux.scala 31:69:@19906.4]
  assign _GEN_3905 = 6'h1 == select_61 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3906 = 6'h2 == select_61 ? io_inData_2 : _GEN_3905; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3907 = 6'h3 == select_61 ? io_inData_3 : _GEN_3906; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3908 = 6'h4 == select_61 ? io_inData_4 : _GEN_3907; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3909 = 6'h5 == select_61 ? io_inData_5 : _GEN_3908; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3910 = 6'h6 == select_61 ? io_inData_6 : _GEN_3909; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3911 = 6'h7 == select_61 ? io_inData_7 : _GEN_3910; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3912 = 6'h8 == select_61 ? io_inData_8 : _GEN_3911; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3913 = 6'h9 == select_61 ? io_inData_9 : _GEN_3912; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3914 = 6'ha == select_61 ? io_inData_10 : _GEN_3913; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3915 = 6'hb == select_61 ? io_inData_11 : _GEN_3914; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3916 = 6'hc == select_61 ? io_inData_12 : _GEN_3915; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3917 = 6'hd == select_61 ? io_inData_13 : _GEN_3916; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3918 = 6'he == select_61 ? io_inData_14 : _GEN_3917; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3919 = 6'hf == select_61 ? io_inData_15 : _GEN_3918; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3920 = 6'h10 == select_61 ? io_inData_16 : _GEN_3919; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3921 = 6'h11 == select_61 ? io_inData_17 : _GEN_3920; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3922 = 6'h12 == select_61 ? io_inData_18 : _GEN_3921; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3923 = 6'h13 == select_61 ? io_inData_19 : _GEN_3922; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3924 = 6'h14 == select_61 ? io_inData_20 : _GEN_3923; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3925 = 6'h15 == select_61 ? io_inData_21 : _GEN_3924; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3926 = 6'h16 == select_61 ? io_inData_22 : _GEN_3925; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3927 = 6'h17 == select_61 ? io_inData_23 : _GEN_3926; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3928 = 6'h18 == select_61 ? io_inData_24 : _GEN_3927; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3929 = 6'h19 == select_61 ? io_inData_25 : _GEN_3928; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3930 = 6'h1a == select_61 ? io_inData_26 : _GEN_3929; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3931 = 6'h1b == select_61 ? io_inData_27 : _GEN_3930; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3932 = 6'h1c == select_61 ? io_inData_28 : _GEN_3931; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3933 = 6'h1d == select_61 ? io_inData_29 : _GEN_3932; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3934 = 6'h1e == select_61 ? io_inData_30 : _GEN_3933; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3935 = 6'h1f == select_61 ? io_inData_31 : _GEN_3934; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3936 = 6'h20 == select_61 ? io_inData_32 : _GEN_3935; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3937 = 6'h21 == select_61 ? io_inData_33 : _GEN_3936; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3938 = 6'h22 == select_61 ? io_inData_34 : _GEN_3937; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3939 = 6'h23 == select_61 ? io_inData_35 : _GEN_3938; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3940 = 6'h24 == select_61 ? io_inData_36 : _GEN_3939; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3941 = 6'h25 == select_61 ? io_inData_37 : _GEN_3940; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3942 = 6'h26 == select_61 ? io_inData_38 : _GEN_3941; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3943 = 6'h27 == select_61 ? io_inData_39 : _GEN_3942; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3944 = 6'h28 == select_61 ? io_inData_40 : _GEN_3943; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3945 = 6'h29 == select_61 ? io_inData_41 : _GEN_3944; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3946 = 6'h2a == select_61 ? io_inData_42 : _GEN_3945; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3947 = 6'h2b == select_61 ? io_inData_43 : _GEN_3946; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3948 = 6'h2c == select_61 ? io_inData_44 : _GEN_3947; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3949 = 6'h2d == select_61 ? io_inData_45 : _GEN_3948; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3950 = 6'h2e == select_61 ? io_inData_46 : _GEN_3949; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3951 = 6'h2f == select_61 ? io_inData_47 : _GEN_3950; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3952 = 6'h30 == select_61 ? io_inData_48 : _GEN_3951; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3953 = 6'h31 == select_61 ? io_inData_49 : _GEN_3952; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3954 = 6'h32 == select_61 ? io_inData_50 : _GEN_3953; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3955 = 6'h33 == select_61 ? io_inData_51 : _GEN_3954; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3956 = 6'h34 == select_61 ? io_inData_52 : _GEN_3955; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3957 = 6'h35 == select_61 ? io_inData_53 : _GEN_3956; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3958 = 6'h36 == select_61 ? io_inData_54 : _GEN_3957; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3959 = 6'h37 == select_61 ? io_inData_55 : _GEN_3958; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3960 = 6'h38 == select_61 ? io_inData_56 : _GEN_3959; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3961 = 6'h39 == select_61 ? io_inData_57 : _GEN_3960; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3962 = 6'h3a == select_61 ? io_inData_58 : _GEN_3961; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3963 = 6'h3b == select_61 ? io_inData_59 : _GEN_3962; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3964 = 6'h3c == select_61 ? io_inData_60 : _GEN_3963; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3965 = 6'h3d == select_61 ? io_inData_61 : _GEN_3964; // @[Switch.scala 33:19:@19908.4]
  assign _GEN_3966 = 6'h3e == select_61 ? io_inData_62 : _GEN_3965; // @[Switch.scala 33:19:@19908.4]
  assign _T_41464 = {valid_61_7,valid_61_6,valid_61_5,valid_61_4,valid_61_3,valid_61_2,valid_61_1,valid_61_0}; // @[Switch.scala 34:32:@19915.4]
  assign _T_41472 = {valid_61_15,valid_61_14,valid_61_13,valid_61_12,valid_61_11,valid_61_10,valid_61_9,valid_61_8,_T_41464}; // @[Switch.scala 34:32:@19923.4]
  assign _T_41479 = {valid_61_23,valid_61_22,valid_61_21,valid_61_20,valid_61_19,valid_61_18,valid_61_17,valid_61_16}; // @[Switch.scala 34:32:@19930.4]
  assign _T_41488 = {valid_61_31,valid_61_30,valid_61_29,valid_61_28,valid_61_27,valid_61_26,valid_61_25,valid_61_24,_T_41479,_T_41472}; // @[Switch.scala 34:32:@19939.4]
  assign _T_41495 = {valid_61_39,valid_61_38,valid_61_37,valid_61_36,valid_61_35,valid_61_34,valid_61_33,valid_61_32}; // @[Switch.scala 34:32:@19946.4]
  assign _T_41503 = {valid_61_47,valid_61_46,valid_61_45,valid_61_44,valid_61_43,valid_61_42,valid_61_41,valid_61_40,_T_41495}; // @[Switch.scala 34:32:@19954.4]
  assign _T_41510 = {valid_61_55,valid_61_54,valid_61_53,valid_61_52,valid_61_51,valid_61_50,valid_61_49,valid_61_48}; // @[Switch.scala 34:32:@19961.4]
  assign _T_41519 = {valid_61_63,valid_61_62,valid_61_61,valid_61_60,valid_61_59,valid_61_58,valid_61_57,valid_61_56,_T_41510,_T_41503}; // @[Switch.scala 34:32:@19970.4]
  assign _T_41520 = {_T_41519,_T_41488}; // @[Switch.scala 34:32:@19971.4]
  assign _T_41524 = io_inAddr_0 == 6'h3e; // @[Switch.scala 30:53:@19974.4]
  assign valid_62_0 = io_inValid_0 & _T_41524; // @[Switch.scala 30:36:@19975.4]
  assign _T_41527 = io_inAddr_1 == 6'h3e; // @[Switch.scala 30:53:@19977.4]
  assign valid_62_1 = io_inValid_1 & _T_41527; // @[Switch.scala 30:36:@19978.4]
  assign _T_41530 = io_inAddr_2 == 6'h3e; // @[Switch.scala 30:53:@19980.4]
  assign valid_62_2 = io_inValid_2 & _T_41530; // @[Switch.scala 30:36:@19981.4]
  assign _T_41533 = io_inAddr_3 == 6'h3e; // @[Switch.scala 30:53:@19983.4]
  assign valid_62_3 = io_inValid_3 & _T_41533; // @[Switch.scala 30:36:@19984.4]
  assign _T_41536 = io_inAddr_4 == 6'h3e; // @[Switch.scala 30:53:@19986.4]
  assign valid_62_4 = io_inValid_4 & _T_41536; // @[Switch.scala 30:36:@19987.4]
  assign _T_41539 = io_inAddr_5 == 6'h3e; // @[Switch.scala 30:53:@19989.4]
  assign valid_62_5 = io_inValid_5 & _T_41539; // @[Switch.scala 30:36:@19990.4]
  assign _T_41542 = io_inAddr_6 == 6'h3e; // @[Switch.scala 30:53:@19992.4]
  assign valid_62_6 = io_inValid_6 & _T_41542; // @[Switch.scala 30:36:@19993.4]
  assign _T_41545 = io_inAddr_7 == 6'h3e; // @[Switch.scala 30:53:@19995.4]
  assign valid_62_7 = io_inValid_7 & _T_41545; // @[Switch.scala 30:36:@19996.4]
  assign _T_41548 = io_inAddr_8 == 6'h3e; // @[Switch.scala 30:53:@19998.4]
  assign valid_62_8 = io_inValid_8 & _T_41548; // @[Switch.scala 30:36:@19999.4]
  assign _T_41551 = io_inAddr_9 == 6'h3e; // @[Switch.scala 30:53:@20001.4]
  assign valid_62_9 = io_inValid_9 & _T_41551; // @[Switch.scala 30:36:@20002.4]
  assign _T_41554 = io_inAddr_10 == 6'h3e; // @[Switch.scala 30:53:@20004.4]
  assign valid_62_10 = io_inValid_10 & _T_41554; // @[Switch.scala 30:36:@20005.4]
  assign _T_41557 = io_inAddr_11 == 6'h3e; // @[Switch.scala 30:53:@20007.4]
  assign valid_62_11 = io_inValid_11 & _T_41557; // @[Switch.scala 30:36:@20008.4]
  assign _T_41560 = io_inAddr_12 == 6'h3e; // @[Switch.scala 30:53:@20010.4]
  assign valid_62_12 = io_inValid_12 & _T_41560; // @[Switch.scala 30:36:@20011.4]
  assign _T_41563 = io_inAddr_13 == 6'h3e; // @[Switch.scala 30:53:@20013.4]
  assign valid_62_13 = io_inValid_13 & _T_41563; // @[Switch.scala 30:36:@20014.4]
  assign _T_41566 = io_inAddr_14 == 6'h3e; // @[Switch.scala 30:53:@20016.4]
  assign valid_62_14 = io_inValid_14 & _T_41566; // @[Switch.scala 30:36:@20017.4]
  assign _T_41569 = io_inAddr_15 == 6'h3e; // @[Switch.scala 30:53:@20019.4]
  assign valid_62_15 = io_inValid_15 & _T_41569; // @[Switch.scala 30:36:@20020.4]
  assign _T_41572 = io_inAddr_16 == 6'h3e; // @[Switch.scala 30:53:@20022.4]
  assign valid_62_16 = io_inValid_16 & _T_41572; // @[Switch.scala 30:36:@20023.4]
  assign _T_41575 = io_inAddr_17 == 6'h3e; // @[Switch.scala 30:53:@20025.4]
  assign valid_62_17 = io_inValid_17 & _T_41575; // @[Switch.scala 30:36:@20026.4]
  assign _T_41578 = io_inAddr_18 == 6'h3e; // @[Switch.scala 30:53:@20028.4]
  assign valid_62_18 = io_inValid_18 & _T_41578; // @[Switch.scala 30:36:@20029.4]
  assign _T_41581 = io_inAddr_19 == 6'h3e; // @[Switch.scala 30:53:@20031.4]
  assign valid_62_19 = io_inValid_19 & _T_41581; // @[Switch.scala 30:36:@20032.4]
  assign _T_41584 = io_inAddr_20 == 6'h3e; // @[Switch.scala 30:53:@20034.4]
  assign valid_62_20 = io_inValid_20 & _T_41584; // @[Switch.scala 30:36:@20035.4]
  assign _T_41587 = io_inAddr_21 == 6'h3e; // @[Switch.scala 30:53:@20037.4]
  assign valid_62_21 = io_inValid_21 & _T_41587; // @[Switch.scala 30:36:@20038.4]
  assign _T_41590 = io_inAddr_22 == 6'h3e; // @[Switch.scala 30:53:@20040.4]
  assign valid_62_22 = io_inValid_22 & _T_41590; // @[Switch.scala 30:36:@20041.4]
  assign _T_41593 = io_inAddr_23 == 6'h3e; // @[Switch.scala 30:53:@20043.4]
  assign valid_62_23 = io_inValid_23 & _T_41593; // @[Switch.scala 30:36:@20044.4]
  assign _T_41596 = io_inAddr_24 == 6'h3e; // @[Switch.scala 30:53:@20046.4]
  assign valid_62_24 = io_inValid_24 & _T_41596; // @[Switch.scala 30:36:@20047.4]
  assign _T_41599 = io_inAddr_25 == 6'h3e; // @[Switch.scala 30:53:@20049.4]
  assign valid_62_25 = io_inValid_25 & _T_41599; // @[Switch.scala 30:36:@20050.4]
  assign _T_41602 = io_inAddr_26 == 6'h3e; // @[Switch.scala 30:53:@20052.4]
  assign valid_62_26 = io_inValid_26 & _T_41602; // @[Switch.scala 30:36:@20053.4]
  assign _T_41605 = io_inAddr_27 == 6'h3e; // @[Switch.scala 30:53:@20055.4]
  assign valid_62_27 = io_inValid_27 & _T_41605; // @[Switch.scala 30:36:@20056.4]
  assign _T_41608 = io_inAddr_28 == 6'h3e; // @[Switch.scala 30:53:@20058.4]
  assign valid_62_28 = io_inValid_28 & _T_41608; // @[Switch.scala 30:36:@20059.4]
  assign _T_41611 = io_inAddr_29 == 6'h3e; // @[Switch.scala 30:53:@20061.4]
  assign valid_62_29 = io_inValid_29 & _T_41611; // @[Switch.scala 30:36:@20062.4]
  assign _T_41614 = io_inAddr_30 == 6'h3e; // @[Switch.scala 30:53:@20064.4]
  assign valid_62_30 = io_inValid_30 & _T_41614; // @[Switch.scala 30:36:@20065.4]
  assign _T_41617 = io_inAddr_31 == 6'h3e; // @[Switch.scala 30:53:@20067.4]
  assign valid_62_31 = io_inValid_31 & _T_41617; // @[Switch.scala 30:36:@20068.4]
  assign _T_41620 = io_inAddr_32 == 6'h3e; // @[Switch.scala 30:53:@20070.4]
  assign valid_62_32 = io_inValid_32 & _T_41620; // @[Switch.scala 30:36:@20071.4]
  assign _T_41623 = io_inAddr_33 == 6'h3e; // @[Switch.scala 30:53:@20073.4]
  assign valid_62_33 = io_inValid_33 & _T_41623; // @[Switch.scala 30:36:@20074.4]
  assign _T_41626 = io_inAddr_34 == 6'h3e; // @[Switch.scala 30:53:@20076.4]
  assign valid_62_34 = io_inValid_34 & _T_41626; // @[Switch.scala 30:36:@20077.4]
  assign _T_41629 = io_inAddr_35 == 6'h3e; // @[Switch.scala 30:53:@20079.4]
  assign valid_62_35 = io_inValid_35 & _T_41629; // @[Switch.scala 30:36:@20080.4]
  assign _T_41632 = io_inAddr_36 == 6'h3e; // @[Switch.scala 30:53:@20082.4]
  assign valid_62_36 = io_inValid_36 & _T_41632; // @[Switch.scala 30:36:@20083.4]
  assign _T_41635 = io_inAddr_37 == 6'h3e; // @[Switch.scala 30:53:@20085.4]
  assign valid_62_37 = io_inValid_37 & _T_41635; // @[Switch.scala 30:36:@20086.4]
  assign _T_41638 = io_inAddr_38 == 6'h3e; // @[Switch.scala 30:53:@20088.4]
  assign valid_62_38 = io_inValid_38 & _T_41638; // @[Switch.scala 30:36:@20089.4]
  assign _T_41641 = io_inAddr_39 == 6'h3e; // @[Switch.scala 30:53:@20091.4]
  assign valid_62_39 = io_inValid_39 & _T_41641; // @[Switch.scala 30:36:@20092.4]
  assign _T_41644 = io_inAddr_40 == 6'h3e; // @[Switch.scala 30:53:@20094.4]
  assign valid_62_40 = io_inValid_40 & _T_41644; // @[Switch.scala 30:36:@20095.4]
  assign _T_41647 = io_inAddr_41 == 6'h3e; // @[Switch.scala 30:53:@20097.4]
  assign valid_62_41 = io_inValid_41 & _T_41647; // @[Switch.scala 30:36:@20098.4]
  assign _T_41650 = io_inAddr_42 == 6'h3e; // @[Switch.scala 30:53:@20100.4]
  assign valid_62_42 = io_inValid_42 & _T_41650; // @[Switch.scala 30:36:@20101.4]
  assign _T_41653 = io_inAddr_43 == 6'h3e; // @[Switch.scala 30:53:@20103.4]
  assign valid_62_43 = io_inValid_43 & _T_41653; // @[Switch.scala 30:36:@20104.4]
  assign _T_41656 = io_inAddr_44 == 6'h3e; // @[Switch.scala 30:53:@20106.4]
  assign valid_62_44 = io_inValid_44 & _T_41656; // @[Switch.scala 30:36:@20107.4]
  assign _T_41659 = io_inAddr_45 == 6'h3e; // @[Switch.scala 30:53:@20109.4]
  assign valid_62_45 = io_inValid_45 & _T_41659; // @[Switch.scala 30:36:@20110.4]
  assign _T_41662 = io_inAddr_46 == 6'h3e; // @[Switch.scala 30:53:@20112.4]
  assign valid_62_46 = io_inValid_46 & _T_41662; // @[Switch.scala 30:36:@20113.4]
  assign _T_41665 = io_inAddr_47 == 6'h3e; // @[Switch.scala 30:53:@20115.4]
  assign valid_62_47 = io_inValid_47 & _T_41665; // @[Switch.scala 30:36:@20116.4]
  assign _T_41668 = io_inAddr_48 == 6'h3e; // @[Switch.scala 30:53:@20118.4]
  assign valid_62_48 = io_inValid_48 & _T_41668; // @[Switch.scala 30:36:@20119.4]
  assign _T_41671 = io_inAddr_49 == 6'h3e; // @[Switch.scala 30:53:@20121.4]
  assign valid_62_49 = io_inValid_49 & _T_41671; // @[Switch.scala 30:36:@20122.4]
  assign _T_41674 = io_inAddr_50 == 6'h3e; // @[Switch.scala 30:53:@20124.4]
  assign valid_62_50 = io_inValid_50 & _T_41674; // @[Switch.scala 30:36:@20125.4]
  assign _T_41677 = io_inAddr_51 == 6'h3e; // @[Switch.scala 30:53:@20127.4]
  assign valid_62_51 = io_inValid_51 & _T_41677; // @[Switch.scala 30:36:@20128.4]
  assign _T_41680 = io_inAddr_52 == 6'h3e; // @[Switch.scala 30:53:@20130.4]
  assign valid_62_52 = io_inValid_52 & _T_41680; // @[Switch.scala 30:36:@20131.4]
  assign _T_41683 = io_inAddr_53 == 6'h3e; // @[Switch.scala 30:53:@20133.4]
  assign valid_62_53 = io_inValid_53 & _T_41683; // @[Switch.scala 30:36:@20134.4]
  assign _T_41686 = io_inAddr_54 == 6'h3e; // @[Switch.scala 30:53:@20136.4]
  assign valid_62_54 = io_inValid_54 & _T_41686; // @[Switch.scala 30:36:@20137.4]
  assign _T_41689 = io_inAddr_55 == 6'h3e; // @[Switch.scala 30:53:@20139.4]
  assign valid_62_55 = io_inValid_55 & _T_41689; // @[Switch.scala 30:36:@20140.4]
  assign _T_41692 = io_inAddr_56 == 6'h3e; // @[Switch.scala 30:53:@20142.4]
  assign valid_62_56 = io_inValid_56 & _T_41692; // @[Switch.scala 30:36:@20143.4]
  assign _T_41695 = io_inAddr_57 == 6'h3e; // @[Switch.scala 30:53:@20145.4]
  assign valid_62_57 = io_inValid_57 & _T_41695; // @[Switch.scala 30:36:@20146.4]
  assign _T_41698 = io_inAddr_58 == 6'h3e; // @[Switch.scala 30:53:@20148.4]
  assign valid_62_58 = io_inValid_58 & _T_41698; // @[Switch.scala 30:36:@20149.4]
  assign _T_41701 = io_inAddr_59 == 6'h3e; // @[Switch.scala 30:53:@20151.4]
  assign valid_62_59 = io_inValid_59 & _T_41701; // @[Switch.scala 30:36:@20152.4]
  assign _T_41704 = io_inAddr_60 == 6'h3e; // @[Switch.scala 30:53:@20154.4]
  assign valid_62_60 = io_inValid_60 & _T_41704; // @[Switch.scala 30:36:@20155.4]
  assign _T_41707 = io_inAddr_61 == 6'h3e; // @[Switch.scala 30:53:@20157.4]
  assign valid_62_61 = io_inValid_61 & _T_41707; // @[Switch.scala 30:36:@20158.4]
  assign _T_41710 = io_inAddr_62 == 6'h3e; // @[Switch.scala 30:53:@20160.4]
  assign valid_62_62 = io_inValid_62 & _T_41710; // @[Switch.scala 30:36:@20161.4]
  assign _T_41713 = io_inAddr_63 == 6'h3e; // @[Switch.scala 30:53:@20163.4]
  assign valid_62_63 = io_inValid_63 & _T_41713; // @[Switch.scala 30:36:@20164.4]
  assign _T_41779 = valid_62_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@20166.4]
  assign _T_41780 = valid_62_61 ? 6'h3d : _T_41779; // @[Mux.scala 31:69:@20167.4]
  assign _T_41781 = valid_62_60 ? 6'h3c : _T_41780; // @[Mux.scala 31:69:@20168.4]
  assign _T_41782 = valid_62_59 ? 6'h3b : _T_41781; // @[Mux.scala 31:69:@20169.4]
  assign _T_41783 = valid_62_58 ? 6'h3a : _T_41782; // @[Mux.scala 31:69:@20170.4]
  assign _T_41784 = valid_62_57 ? 6'h39 : _T_41783; // @[Mux.scala 31:69:@20171.4]
  assign _T_41785 = valid_62_56 ? 6'h38 : _T_41784; // @[Mux.scala 31:69:@20172.4]
  assign _T_41786 = valid_62_55 ? 6'h37 : _T_41785; // @[Mux.scala 31:69:@20173.4]
  assign _T_41787 = valid_62_54 ? 6'h36 : _T_41786; // @[Mux.scala 31:69:@20174.4]
  assign _T_41788 = valid_62_53 ? 6'h35 : _T_41787; // @[Mux.scala 31:69:@20175.4]
  assign _T_41789 = valid_62_52 ? 6'h34 : _T_41788; // @[Mux.scala 31:69:@20176.4]
  assign _T_41790 = valid_62_51 ? 6'h33 : _T_41789; // @[Mux.scala 31:69:@20177.4]
  assign _T_41791 = valid_62_50 ? 6'h32 : _T_41790; // @[Mux.scala 31:69:@20178.4]
  assign _T_41792 = valid_62_49 ? 6'h31 : _T_41791; // @[Mux.scala 31:69:@20179.4]
  assign _T_41793 = valid_62_48 ? 6'h30 : _T_41792; // @[Mux.scala 31:69:@20180.4]
  assign _T_41794 = valid_62_47 ? 6'h2f : _T_41793; // @[Mux.scala 31:69:@20181.4]
  assign _T_41795 = valid_62_46 ? 6'h2e : _T_41794; // @[Mux.scala 31:69:@20182.4]
  assign _T_41796 = valid_62_45 ? 6'h2d : _T_41795; // @[Mux.scala 31:69:@20183.4]
  assign _T_41797 = valid_62_44 ? 6'h2c : _T_41796; // @[Mux.scala 31:69:@20184.4]
  assign _T_41798 = valid_62_43 ? 6'h2b : _T_41797; // @[Mux.scala 31:69:@20185.4]
  assign _T_41799 = valid_62_42 ? 6'h2a : _T_41798; // @[Mux.scala 31:69:@20186.4]
  assign _T_41800 = valid_62_41 ? 6'h29 : _T_41799; // @[Mux.scala 31:69:@20187.4]
  assign _T_41801 = valid_62_40 ? 6'h28 : _T_41800; // @[Mux.scala 31:69:@20188.4]
  assign _T_41802 = valid_62_39 ? 6'h27 : _T_41801; // @[Mux.scala 31:69:@20189.4]
  assign _T_41803 = valid_62_38 ? 6'h26 : _T_41802; // @[Mux.scala 31:69:@20190.4]
  assign _T_41804 = valid_62_37 ? 6'h25 : _T_41803; // @[Mux.scala 31:69:@20191.4]
  assign _T_41805 = valid_62_36 ? 6'h24 : _T_41804; // @[Mux.scala 31:69:@20192.4]
  assign _T_41806 = valid_62_35 ? 6'h23 : _T_41805; // @[Mux.scala 31:69:@20193.4]
  assign _T_41807 = valid_62_34 ? 6'h22 : _T_41806; // @[Mux.scala 31:69:@20194.4]
  assign _T_41808 = valid_62_33 ? 6'h21 : _T_41807; // @[Mux.scala 31:69:@20195.4]
  assign _T_41809 = valid_62_32 ? 6'h20 : _T_41808; // @[Mux.scala 31:69:@20196.4]
  assign _T_41810 = valid_62_31 ? 6'h1f : _T_41809; // @[Mux.scala 31:69:@20197.4]
  assign _T_41811 = valid_62_30 ? 6'h1e : _T_41810; // @[Mux.scala 31:69:@20198.4]
  assign _T_41812 = valid_62_29 ? 6'h1d : _T_41811; // @[Mux.scala 31:69:@20199.4]
  assign _T_41813 = valid_62_28 ? 6'h1c : _T_41812; // @[Mux.scala 31:69:@20200.4]
  assign _T_41814 = valid_62_27 ? 6'h1b : _T_41813; // @[Mux.scala 31:69:@20201.4]
  assign _T_41815 = valid_62_26 ? 6'h1a : _T_41814; // @[Mux.scala 31:69:@20202.4]
  assign _T_41816 = valid_62_25 ? 6'h19 : _T_41815; // @[Mux.scala 31:69:@20203.4]
  assign _T_41817 = valid_62_24 ? 6'h18 : _T_41816; // @[Mux.scala 31:69:@20204.4]
  assign _T_41818 = valid_62_23 ? 6'h17 : _T_41817; // @[Mux.scala 31:69:@20205.4]
  assign _T_41819 = valid_62_22 ? 6'h16 : _T_41818; // @[Mux.scala 31:69:@20206.4]
  assign _T_41820 = valid_62_21 ? 6'h15 : _T_41819; // @[Mux.scala 31:69:@20207.4]
  assign _T_41821 = valid_62_20 ? 6'h14 : _T_41820; // @[Mux.scala 31:69:@20208.4]
  assign _T_41822 = valid_62_19 ? 6'h13 : _T_41821; // @[Mux.scala 31:69:@20209.4]
  assign _T_41823 = valid_62_18 ? 6'h12 : _T_41822; // @[Mux.scala 31:69:@20210.4]
  assign _T_41824 = valid_62_17 ? 6'h11 : _T_41823; // @[Mux.scala 31:69:@20211.4]
  assign _T_41825 = valid_62_16 ? 6'h10 : _T_41824; // @[Mux.scala 31:69:@20212.4]
  assign _T_41826 = valid_62_15 ? 6'hf : _T_41825; // @[Mux.scala 31:69:@20213.4]
  assign _T_41827 = valid_62_14 ? 6'he : _T_41826; // @[Mux.scala 31:69:@20214.4]
  assign _T_41828 = valid_62_13 ? 6'hd : _T_41827; // @[Mux.scala 31:69:@20215.4]
  assign _T_41829 = valid_62_12 ? 6'hc : _T_41828; // @[Mux.scala 31:69:@20216.4]
  assign _T_41830 = valid_62_11 ? 6'hb : _T_41829; // @[Mux.scala 31:69:@20217.4]
  assign _T_41831 = valid_62_10 ? 6'ha : _T_41830; // @[Mux.scala 31:69:@20218.4]
  assign _T_41832 = valid_62_9 ? 6'h9 : _T_41831; // @[Mux.scala 31:69:@20219.4]
  assign _T_41833 = valid_62_8 ? 6'h8 : _T_41832; // @[Mux.scala 31:69:@20220.4]
  assign _T_41834 = valid_62_7 ? 6'h7 : _T_41833; // @[Mux.scala 31:69:@20221.4]
  assign _T_41835 = valid_62_6 ? 6'h6 : _T_41834; // @[Mux.scala 31:69:@20222.4]
  assign _T_41836 = valid_62_5 ? 6'h5 : _T_41835; // @[Mux.scala 31:69:@20223.4]
  assign _T_41837 = valid_62_4 ? 6'h4 : _T_41836; // @[Mux.scala 31:69:@20224.4]
  assign _T_41838 = valid_62_3 ? 6'h3 : _T_41837; // @[Mux.scala 31:69:@20225.4]
  assign _T_41839 = valid_62_2 ? 6'h2 : _T_41838; // @[Mux.scala 31:69:@20226.4]
  assign _T_41840 = valid_62_1 ? 6'h1 : _T_41839; // @[Mux.scala 31:69:@20227.4]
  assign select_62 = valid_62_0 ? 6'h0 : _T_41840; // @[Mux.scala 31:69:@20228.4]
  assign _GEN_3969 = 6'h1 == select_62 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_3970 = 6'h2 == select_62 ? io_inData_2 : _GEN_3969; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_3971 = 6'h3 == select_62 ? io_inData_3 : _GEN_3970; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_3972 = 6'h4 == select_62 ? io_inData_4 : _GEN_3971; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_3973 = 6'h5 == select_62 ? io_inData_5 : _GEN_3972; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_3974 = 6'h6 == select_62 ? io_inData_6 : _GEN_3973; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_3975 = 6'h7 == select_62 ? io_inData_7 : _GEN_3974; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_3976 = 6'h8 == select_62 ? io_inData_8 : _GEN_3975; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_3977 = 6'h9 == select_62 ? io_inData_9 : _GEN_3976; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_3978 = 6'ha == select_62 ? io_inData_10 : _GEN_3977; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_3979 = 6'hb == select_62 ? io_inData_11 : _GEN_3978; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_3980 = 6'hc == select_62 ? io_inData_12 : _GEN_3979; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_3981 = 6'hd == select_62 ? io_inData_13 : _GEN_3980; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_3982 = 6'he == select_62 ? io_inData_14 : _GEN_3981; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_3983 = 6'hf == select_62 ? io_inData_15 : _GEN_3982; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_3984 = 6'h10 == select_62 ? io_inData_16 : _GEN_3983; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_3985 = 6'h11 == select_62 ? io_inData_17 : _GEN_3984; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_3986 = 6'h12 == select_62 ? io_inData_18 : _GEN_3985; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_3987 = 6'h13 == select_62 ? io_inData_19 : _GEN_3986; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_3988 = 6'h14 == select_62 ? io_inData_20 : _GEN_3987; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_3989 = 6'h15 == select_62 ? io_inData_21 : _GEN_3988; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_3990 = 6'h16 == select_62 ? io_inData_22 : _GEN_3989; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_3991 = 6'h17 == select_62 ? io_inData_23 : _GEN_3990; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_3992 = 6'h18 == select_62 ? io_inData_24 : _GEN_3991; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_3993 = 6'h19 == select_62 ? io_inData_25 : _GEN_3992; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_3994 = 6'h1a == select_62 ? io_inData_26 : _GEN_3993; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_3995 = 6'h1b == select_62 ? io_inData_27 : _GEN_3994; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_3996 = 6'h1c == select_62 ? io_inData_28 : _GEN_3995; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_3997 = 6'h1d == select_62 ? io_inData_29 : _GEN_3996; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_3998 = 6'h1e == select_62 ? io_inData_30 : _GEN_3997; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_3999 = 6'h1f == select_62 ? io_inData_31 : _GEN_3998; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_4000 = 6'h20 == select_62 ? io_inData_32 : _GEN_3999; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_4001 = 6'h21 == select_62 ? io_inData_33 : _GEN_4000; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_4002 = 6'h22 == select_62 ? io_inData_34 : _GEN_4001; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_4003 = 6'h23 == select_62 ? io_inData_35 : _GEN_4002; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_4004 = 6'h24 == select_62 ? io_inData_36 : _GEN_4003; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_4005 = 6'h25 == select_62 ? io_inData_37 : _GEN_4004; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_4006 = 6'h26 == select_62 ? io_inData_38 : _GEN_4005; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_4007 = 6'h27 == select_62 ? io_inData_39 : _GEN_4006; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_4008 = 6'h28 == select_62 ? io_inData_40 : _GEN_4007; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_4009 = 6'h29 == select_62 ? io_inData_41 : _GEN_4008; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_4010 = 6'h2a == select_62 ? io_inData_42 : _GEN_4009; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_4011 = 6'h2b == select_62 ? io_inData_43 : _GEN_4010; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_4012 = 6'h2c == select_62 ? io_inData_44 : _GEN_4011; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_4013 = 6'h2d == select_62 ? io_inData_45 : _GEN_4012; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_4014 = 6'h2e == select_62 ? io_inData_46 : _GEN_4013; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_4015 = 6'h2f == select_62 ? io_inData_47 : _GEN_4014; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_4016 = 6'h30 == select_62 ? io_inData_48 : _GEN_4015; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_4017 = 6'h31 == select_62 ? io_inData_49 : _GEN_4016; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_4018 = 6'h32 == select_62 ? io_inData_50 : _GEN_4017; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_4019 = 6'h33 == select_62 ? io_inData_51 : _GEN_4018; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_4020 = 6'h34 == select_62 ? io_inData_52 : _GEN_4019; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_4021 = 6'h35 == select_62 ? io_inData_53 : _GEN_4020; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_4022 = 6'h36 == select_62 ? io_inData_54 : _GEN_4021; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_4023 = 6'h37 == select_62 ? io_inData_55 : _GEN_4022; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_4024 = 6'h38 == select_62 ? io_inData_56 : _GEN_4023; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_4025 = 6'h39 == select_62 ? io_inData_57 : _GEN_4024; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_4026 = 6'h3a == select_62 ? io_inData_58 : _GEN_4025; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_4027 = 6'h3b == select_62 ? io_inData_59 : _GEN_4026; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_4028 = 6'h3c == select_62 ? io_inData_60 : _GEN_4027; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_4029 = 6'h3d == select_62 ? io_inData_61 : _GEN_4028; // @[Switch.scala 33:19:@20230.4]
  assign _GEN_4030 = 6'h3e == select_62 ? io_inData_62 : _GEN_4029; // @[Switch.scala 33:19:@20230.4]
  assign _T_41849 = {valid_62_7,valid_62_6,valid_62_5,valid_62_4,valid_62_3,valid_62_2,valid_62_1,valid_62_0}; // @[Switch.scala 34:32:@20237.4]
  assign _T_41857 = {valid_62_15,valid_62_14,valid_62_13,valid_62_12,valid_62_11,valid_62_10,valid_62_9,valid_62_8,_T_41849}; // @[Switch.scala 34:32:@20245.4]
  assign _T_41864 = {valid_62_23,valid_62_22,valid_62_21,valid_62_20,valid_62_19,valid_62_18,valid_62_17,valid_62_16}; // @[Switch.scala 34:32:@20252.4]
  assign _T_41873 = {valid_62_31,valid_62_30,valid_62_29,valid_62_28,valid_62_27,valid_62_26,valid_62_25,valid_62_24,_T_41864,_T_41857}; // @[Switch.scala 34:32:@20261.4]
  assign _T_41880 = {valid_62_39,valid_62_38,valid_62_37,valid_62_36,valid_62_35,valid_62_34,valid_62_33,valid_62_32}; // @[Switch.scala 34:32:@20268.4]
  assign _T_41888 = {valid_62_47,valid_62_46,valid_62_45,valid_62_44,valid_62_43,valid_62_42,valid_62_41,valid_62_40,_T_41880}; // @[Switch.scala 34:32:@20276.4]
  assign _T_41895 = {valid_62_55,valid_62_54,valid_62_53,valid_62_52,valid_62_51,valid_62_50,valid_62_49,valid_62_48}; // @[Switch.scala 34:32:@20283.4]
  assign _T_41904 = {valid_62_63,valid_62_62,valid_62_61,valid_62_60,valid_62_59,valid_62_58,valid_62_57,valid_62_56,_T_41895,_T_41888}; // @[Switch.scala 34:32:@20292.4]
  assign _T_41905 = {_T_41904,_T_41873}; // @[Switch.scala 34:32:@20293.4]
  assign _T_41909 = io_inAddr_0 == 6'h3f; // @[Switch.scala 30:53:@20296.4]
  assign valid_63_0 = io_inValid_0 & _T_41909; // @[Switch.scala 30:36:@20297.4]
  assign _T_41912 = io_inAddr_1 == 6'h3f; // @[Switch.scala 30:53:@20299.4]
  assign valid_63_1 = io_inValid_1 & _T_41912; // @[Switch.scala 30:36:@20300.4]
  assign _T_41915 = io_inAddr_2 == 6'h3f; // @[Switch.scala 30:53:@20302.4]
  assign valid_63_2 = io_inValid_2 & _T_41915; // @[Switch.scala 30:36:@20303.4]
  assign _T_41918 = io_inAddr_3 == 6'h3f; // @[Switch.scala 30:53:@20305.4]
  assign valid_63_3 = io_inValid_3 & _T_41918; // @[Switch.scala 30:36:@20306.4]
  assign _T_41921 = io_inAddr_4 == 6'h3f; // @[Switch.scala 30:53:@20308.4]
  assign valid_63_4 = io_inValid_4 & _T_41921; // @[Switch.scala 30:36:@20309.4]
  assign _T_41924 = io_inAddr_5 == 6'h3f; // @[Switch.scala 30:53:@20311.4]
  assign valid_63_5 = io_inValid_5 & _T_41924; // @[Switch.scala 30:36:@20312.4]
  assign _T_41927 = io_inAddr_6 == 6'h3f; // @[Switch.scala 30:53:@20314.4]
  assign valid_63_6 = io_inValid_6 & _T_41927; // @[Switch.scala 30:36:@20315.4]
  assign _T_41930 = io_inAddr_7 == 6'h3f; // @[Switch.scala 30:53:@20317.4]
  assign valid_63_7 = io_inValid_7 & _T_41930; // @[Switch.scala 30:36:@20318.4]
  assign _T_41933 = io_inAddr_8 == 6'h3f; // @[Switch.scala 30:53:@20320.4]
  assign valid_63_8 = io_inValid_8 & _T_41933; // @[Switch.scala 30:36:@20321.4]
  assign _T_41936 = io_inAddr_9 == 6'h3f; // @[Switch.scala 30:53:@20323.4]
  assign valid_63_9 = io_inValid_9 & _T_41936; // @[Switch.scala 30:36:@20324.4]
  assign _T_41939 = io_inAddr_10 == 6'h3f; // @[Switch.scala 30:53:@20326.4]
  assign valid_63_10 = io_inValid_10 & _T_41939; // @[Switch.scala 30:36:@20327.4]
  assign _T_41942 = io_inAddr_11 == 6'h3f; // @[Switch.scala 30:53:@20329.4]
  assign valid_63_11 = io_inValid_11 & _T_41942; // @[Switch.scala 30:36:@20330.4]
  assign _T_41945 = io_inAddr_12 == 6'h3f; // @[Switch.scala 30:53:@20332.4]
  assign valid_63_12 = io_inValid_12 & _T_41945; // @[Switch.scala 30:36:@20333.4]
  assign _T_41948 = io_inAddr_13 == 6'h3f; // @[Switch.scala 30:53:@20335.4]
  assign valid_63_13 = io_inValid_13 & _T_41948; // @[Switch.scala 30:36:@20336.4]
  assign _T_41951 = io_inAddr_14 == 6'h3f; // @[Switch.scala 30:53:@20338.4]
  assign valid_63_14 = io_inValid_14 & _T_41951; // @[Switch.scala 30:36:@20339.4]
  assign _T_41954 = io_inAddr_15 == 6'h3f; // @[Switch.scala 30:53:@20341.4]
  assign valid_63_15 = io_inValid_15 & _T_41954; // @[Switch.scala 30:36:@20342.4]
  assign _T_41957 = io_inAddr_16 == 6'h3f; // @[Switch.scala 30:53:@20344.4]
  assign valid_63_16 = io_inValid_16 & _T_41957; // @[Switch.scala 30:36:@20345.4]
  assign _T_41960 = io_inAddr_17 == 6'h3f; // @[Switch.scala 30:53:@20347.4]
  assign valid_63_17 = io_inValid_17 & _T_41960; // @[Switch.scala 30:36:@20348.4]
  assign _T_41963 = io_inAddr_18 == 6'h3f; // @[Switch.scala 30:53:@20350.4]
  assign valid_63_18 = io_inValid_18 & _T_41963; // @[Switch.scala 30:36:@20351.4]
  assign _T_41966 = io_inAddr_19 == 6'h3f; // @[Switch.scala 30:53:@20353.4]
  assign valid_63_19 = io_inValid_19 & _T_41966; // @[Switch.scala 30:36:@20354.4]
  assign _T_41969 = io_inAddr_20 == 6'h3f; // @[Switch.scala 30:53:@20356.4]
  assign valid_63_20 = io_inValid_20 & _T_41969; // @[Switch.scala 30:36:@20357.4]
  assign _T_41972 = io_inAddr_21 == 6'h3f; // @[Switch.scala 30:53:@20359.4]
  assign valid_63_21 = io_inValid_21 & _T_41972; // @[Switch.scala 30:36:@20360.4]
  assign _T_41975 = io_inAddr_22 == 6'h3f; // @[Switch.scala 30:53:@20362.4]
  assign valid_63_22 = io_inValid_22 & _T_41975; // @[Switch.scala 30:36:@20363.4]
  assign _T_41978 = io_inAddr_23 == 6'h3f; // @[Switch.scala 30:53:@20365.4]
  assign valid_63_23 = io_inValid_23 & _T_41978; // @[Switch.scala 30:36:@20366.4]
  assign _T_41981 = io_inAddr_24 == 6'h3f; // @[Switch.scala 30:53:@20368.4]
  assign valid_63_24 = io_inValid_24 & _T_41981; // @[Switch.scala 30:36:@20369.4]
  assign _T_41984 = io_inAddr_25 == 6'h3f; // @[Switch.scala 30:53:@20371.4]
  assign valid_63_25 = io_inValid_25 & _T_41984; // @[Switch.scala 30:36:@20372.4]
  assign _T_41987 = io_inAddr_26 == 6'h3f; // @[Switch.scala 30:53:@20374.4]
  assign valid_63_26 = io_inValid_26 & _T_41987; // @[Switch.scala 30:36:@20375.4]
  assign _T_41990 = io_inAddr_27 == 6'h3f; // @[Switch.scala 30:53:@20377.4]
  assign valid_63_27 = io_inValid_27 & _T_41990; // @[Switch.scala 30:36:@20378.4]
  assign _T_41993 = io_inAddr_28 == 6'h3f; // @[Switch.scala 30:53:@20380.4]
  assign valid_63_28 = io_inValid_28 & _T_41993; // @[Switch.scala 30:36:@20381.4]
  assign _T_41996 = io_inAddr_29 == 6'h3f; // @[Switch.scala 30:53:@20383.4]
  assign valid_63_29 = io_inValid_29 & _T_41996; // @[Switch.scala 30:36:@20384.4]
  assign _T_41999 = io_inAddr_30 == 6'h3f; // @[Switch.scala 30:53:@20386.4]
  assign valid_63_30 = io_inValid_30 & _T_41999; // @[Switch.scala 30:36:@20387.4]
  assign _T_42002 = io_inAddr_31 == 6'h3f; // @[Switch.scala 30:53:@20389.4]
  assign valid_63_31 = io_inValid_31 & _T_42002; // @[Switch.scala 30:36:@20390.4]
  assign _T_42005 = io_inAddr_32 == 6'h3f; // @[Switch.scala 30:53:@20392.4]
  assign valid_63_32 = io_inValid_32 & _T_42005; // @[Switch.scala 30:36:@20393.4]
  assign _T_42008 = io_inAddr_33 == 6'h3f; // @[Switch.scala 30:53:@20395.4]
  assign valid_63_33 = io_inValid_33 & _T_42008; // @[Switch.scala 30:36:@20396.4]
  assign _T_42011 = io_inAddr_34 == 6'h3f; // @[Switch.scala 30:53:@20398.4]
  assign valid_63_34 = io_inValid_34 & _T_42011; // @[Switch.scala 30:36:@20399.4]
  assign _T_42014 = io_inAddr_35 == 6'h3f; // @[Switch.scala 30:53:@20401.4]
  assign valid_63_35 = io_inValid_35 & _T_42014; // @[Switch.scala 30:36:@20402.4]
  assign _T_42017 = io_inAddr_36 == 6'h3f; // @[Switch.scala 30:53:@20404.4]
  assign valid_63_36 = io_inValid_36 & _T_42017; // @[Switch.scala 30:36:@20405.4]
  assign _T_42020 = io_inAddr_37 == 6'h3f; // @[Switch.scala 30:53:@20407.4]
  assign valid_63_37 = io_inValid_37 & _T_42020; // @[Switch.scala 30:36:@20408.4]
  assign _T_42023 = io_inAddr_38 == 6'h3f; // @[Switch.scala 30:53:@20410.4]
  assign valid_63_38 = io_inValid_38 & _T_42023; // @[Switch.scala 30:36:@20411.4]
  assign _T_42026 = io_inAddr_39 == 6'h3f; // @[Switch.scala 30:53:@20413.4]
  assign valid_63_39 = io_inValid_39 & _T_42026; // @[Switch.scala 30:36:@20414.4]
  assign _T_42029 = io_inAddr_40 == 6'h3f; // @[Switch.scala 30:53:@20416.4]
  assign valid_63_40 = io_inValid_40 & _T_42029; // @[Switch.scala 30:36:@20417.4]
  assign _T_42032 = io_inAddr_41 == 6'h3f; // @[Switch.scala 30:53:@20419.4]
  assign valid_63_41 = io_inValid_41 & _T_42032; // @[Switch.scala 30:36:@20420.4]
  assign _T_42035 = io_inAddr_42 == 6'h3f; // @[Switch.scala 30:53:@20422.4]
  assign valid_63_42 = io_inValid_42 & _T_42035; // @[Switch.scala 30:36:@20423.4]
  assign _T_42038 = io_inAddr_43 == 6'h3f; // @[Switch.scala 30:53:@20425.4]
  assign valid_63_43 = io_inValid_43 & _T_42038; // @[Switch.scala 30:36:@20426.4]
  assign _T_42041 = io_inAddr_44 == 6'h3f; // @[Switch.scala 30:53:@20428.4]
  assign valid_63_44 = io_inValid_44 & _T_42041; // @[Switch.scala 30:36:@20429.4]
  assign _T_42044 = io_inAddr_45 == 6'h3f; // @[Switch.scala 30:53:@20431.4]
  assign valid_63_45 = io_inValid_45 & _T_42044; // @[Switch.scala 30:36:@20432.4]
  assign _T_42047 = io_inAddr_46 == 6'h3f; // @[Switch.scala 30:53:@20434.4]
  assign valid_63_46 = io_inValid_46 & _T_42047; // @[Switch.scala 30:36:@20435.4]
  assign _T_42050 = io_inAddr_47 == 6'h3f; // @[Switch.scala 30:53:@20437.4]
  assign valid_63_47 = io_inValid_47 & _T_42050; // @[Switch.scala 30:36:@20438.4]
  assign _T_42053 = io_inAddr_48 == 6'h3f; // @[Switch.scala 30:53:@20440.4]
  assign valid_63_48 = io_inValid_48 & _T_42053; // @[Switch.scala 30:36:@20441.4]
  assign _T_42056 = io_inAddr_49 == 6'h3f; // @[Switch.scala 30:53:@20443.4]
  assign valid_63_49 = io_inValid_49 & _T_42056; // @[Switch.scala 30:36:@20444.4]
  assign _T_42059 = io_inAddr_50 == 6'h3f; // @[Switch.scala 30:53:@20446.4]
  assign valid_63_50 = io_inValid_50 & _T_42059; // @[Switch.scala 30:36:@20447.4]
  assign _T_42062 = io_inAddr_51 == 6'h3f; // @[Switch.scala 30:53:@20449.4]
  assign valid_63_51 = io_inValid_51 & _T_42062; // @[Switch.scala 30:36:@20450.4]
  assign _T_42065 = io_inAddr_52 == 6'h3f; // @[Switch.scala 30:53:@20452.4]
  assign valid_63_52 = io_inValid_52 & _T_42065; // @[Switch.scala 30:36:@20453.4]
  assign _T_42068 = io_inAddr_53 == 6'h3f; // @[Switch.scala 30:53:@20455.4]
  assign valid_63_53 = io_inValid_53 & _T_42068; // @[Switch.scala 30:36:@20456.4]
  assign _T_42071 = io_inAddr_54 == 6'h3f; // @[Switch.scala 30:53:@20458.4]
  assign valid_63_54 = io_inValid_54 & _T_42071; // @[Switch.scala 30:36:@20459.4]
  assign _T_42074 = io_inAddr_55 == 6'h3f; // @[Switch.scala 30:53:@20461.4]
  assign valid_63_55 = io_inValid_55 & _T_42074; // @[Switch.scala 30:36:@20462.4]
  assign _T_42077 = io_inAddr_56 == 6'h3f; // @[Switch.scala 30:53:@20464.4]
  assign valid_63_56 = io_inValid_56 & _T_42077; // @[Switch.scala 30:36:@20465.4]
  assign _T_42080 = io_inAddr_57 == 6'h3f; // @[Switch.scala 30:53:@20467.4]
  assign valid_63_57 = io_inValid_57 & _T_42080; // @[Switch.scala 30:36:@20468.4]
  assign _T_42083 = io_inAddr_58 == 6'h3f; // @[Switch.scala 30:53:@20470.4]
  assign valid_63_58 = io_inValid_58 & _T_42083; // @[Switch.scala 30:36:@20471.4]
  assign _T_42086 = io_inAddr_59 == 6'h3f; // @[Switch.scala 30:53:@20473.4]
  assign valid_63_59 = io_inValid_59 & _T_42086; // @[Switch.scala 30:36:@20474.4]
  assign _T_42089 = io_inAddr_60 == 6'h3f; // @[Switch.scala 30:53:@20476.4]
  assign valid_63_60 = io_inValid_60 & _T_42089; // @[Switch.scala 30:36:@20477.4]
  assign _T_42092 = io_inAddr_61 == 6'h3f; // @[Switch.scala 30:53:@20479.4]
  assign valid_63_61 = io_inValid_61 & _T_42092; // @[Switch.scala 30:36:@20480.4]
  assign _T_42095 = io_inAddr_62 == 6'h3f; // @[Switch.scala 30:53:@20482.4]
  assign valid_63_62 = io_inValid_62 & _T_42095; // @[Switch.scala 30:36:@20483.4]
  assign _T_42098 = io_inAddr_63 == 6'h3f; // @[Switch.scala 30:53:@20485.4]
  assign valid_63_63 = io_inValid_63 & _T_42098; // @[Switch.scala 30:36:@20486.4]
  assign _T_42164 = valid_63_62 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@20488.4]
  assign _T_42165 = valid_63_61 ? 6'h3d : _T_42164; // @[Mux.scala 31:69:@20489.4]
  assign _T_42166 = valid_63_60 ? 6'h3c : _T_42165; // @[Mux.scala 31:69:@20490.4]
  assign _T_42167 = valid_63_59 ? 6'h3b : _T_42166; // @[Mux.scala 31:69:@20491.4]
  assign _T_42168 = valid_63_58 ? 6'h3a : _T_42167; // @[Mux.scala 31:69:@20492.4]
  assign _T_42169 = valid_63_57 ? 6'h39 : _T_42168; // @[Mux.scala 31:69:@20493.4]
  assign _T_42170 = valid_63_56 ? 6'h38 : _T_42169; // @[Mux.scala 31:69:@20494.4]
  assign _T_42171 = valid_63_55 ? 6'h37 : _T_42170; // @[Mux.scala 31:69:@20495.4]
  assign _T_42172 = valid_63_54 ? 6'h36 : _T_42171; // @[Mux.scala 31:69:@20496.4]
  assign _T_42173 = valid_63_53 ? 6'h35 : _T_42172; // @[Mux.scala 31:69:@20497.4]
  assign _T_42174 = valid_63_52 ? 6'h34 : _T_42173; // @[Mux.scala 31:69:@20498.4]
  assign _T_42175 = valid_63_51 ? 6'h33 : _T_42174; // @[Mux.scala 31:69:@20499.4]
  assign _T_42176 = valid_63_50 ? 6'h32 : _T_42175; // @[Mux.scala 31:69:@20500.4]
  assign _T_42177 = valid_63_49 ? 6'h31 : _T_42176; // @[Mux.scala 31:69:@20501.4]
  assign _T_42178 = valid_63_48 ? 6'h30 : _T_42177; // @[Mux.scala 31:69:@20502.4]
  assign _T_42179 = valid_63_47 ? 6'h2f : _T_42178; // @[Mux.scala 31:69:@20503.4]
  assign _T_42180 = valid_63_46 ? 6'h2e : _T_42179; // @[Mux.scala 31:69:@20504.4]
  assign _T_42181 = valid_63_45 ? 6'h2d : _T_42180; // @[Mux.scala 31:69:@20505.4]
  assign _T_42182 = valid_63_44 ? 6'h2c : _T_42181; // @[Mux.scala 31:69:@20506.4]
  assign _T_42183 = valid_63_43 ? 6'h2b : _T_42182; // @[Mux.scala 31:69:@20507.4]
  assign _T_42184 = valid_63_42 ? 6'h2a : _T_42183; // @[Mux.scala 31:69:@20508.4]
  assign _T_42185 = valid_63_41 ? 6'h29 : _T_42184; // @[Mux.scala 31:69:@20509.4]
  assign _T_42186 = valid_63_40 ? 6'h28 : _T_42185; // @[Mux.scala 31:69:@20510.4]
  assign _T_42187 = valid_63_39 ? 6'h27 : _T_42186; // @[Mux.scala 31:69:@20511.4]
  assign _T_42188 = valid_63_38 ? 6'h26 : _T_42187; // @[Mux.scala 31:69:@20512.4]
  assign _T_42189 = valid_63_37 ? 6'h25 : _T_42188; // @[Mux.scala 31:69:@20513.4]
  assign _T_42190 = valid_63_36 ? 6'h24 : _T_42189; // @[Mux.scala 31:69:@20514.4]
  assign _T_42191 = valid_63_35 ? 6'h23 : _T_42190; // @[Mux.scala 31:69:@20515.4]
  assign _T_42192 = valid_63_34 ? 6'h22 : _T_42191; // @[Mux.scala 31:69:@20516.4]
  assign _T_42193 = valid_63_33 ? 6'h21 : _T_42192; // @[Mux.scala 31:69:@20517.4]
  assign _T_42194 = valid_63_32 ? 6'h20 : _T_42193; // @[Mux.scala 31:69:@20518.4]
  assign _T_42195 = valid_63_31 ? 6'h1f : _T_42194; // @[Mux.scala 31:69:@20519.4]
  assign _T_42196 = valid_63_30 ? 6'h1e : _T_42195; // @[Mux.scala 31:69:@20520.4]
  assign _T_42197 = valid_63_29 ? 6'h1d : _T_42196; // @[Mux.scala 31:69:@20521.4]
  assign _T_42198 = valid_63_28 ? 6'h1c : _T_42197; // @[Mux.scala 31:69:@20522.4]
  assign _T_42199 = valid_63_27 ? 6'h1b : _T_42198; // @[Mux.scala 31:69:@20523.4]
  assign _T_42200 = valid_63_26 ? 6'h1a : _T_42199; // @[Mux.scala 31:69:@20524.4]
  assign _T_42201 = valid_63_25 ? 6'h19 : _T_42200; // @[Mux.scala 31:69:@20525.4]
  assign _T_42202 = valid_63_24 ? 6'h18 : _T_42201; // @[Mux.scala 31:69:@20526.4]
  assign _T_42203 = valid_63_23 ? 6'h17 : _T_42202; // @[Mux.scala 31:69:@20527.4]
  assign _T_42204 = valid_63_22 ? 6'h16 : _T_42203; // @[Mux.scala 31:69:@20528.4]
  assign _T_42205 = valid_63_21 ? 6'h15 : _T_42204; // @[Mux.scala 31:69:@20529.4]
  assign _T_42206 = valid_63_20 ? 6'h14 : _T_42205; // @[Mux.scala 31:69:@20530.4]
  assign _T_42207 = valid_63_19 ? 6'h13 : _T_42206; // @[Mux.scala 31:69:@20531.4]
  assign _T_42208 = valid_63_18 ? 6'h12 : _T_42207; // @[Mux.scala 31:69:@20532.4]
  assign _T_42209 = valid_63_17 ? 6'h11 : _T_42208; // @[Mux.scala 31:69:@20533.4]
  assign _T_42210 = valid_63_16 ? 6'h10 : _T_42209; // @[Mux.scala 31:69:@20534.4]
  assign _T_42211 = valid_63_15 ? 6'hf : _T_42210; // @[Mux.scala 31:69:@20535.4]
  assign _T_42212 = valid_63_14 ? 6'he : _T_42211; // @[Mux.scala 31:69:@20536.4]
  assign _T_42213 = valid_63_13 ? 6'hd : _T_42212; // @[Mux.scala 31:69:@20537.4]
  assign _T_42214 = valid_63_12 ? 6'hc : _T_42213; // @[Mux.scala 31:69:@20538.4]
  assign _T_42215 = valid_63_11 ? 6'hb : _T_42214; // @[Mux.scala 31:69:@20539.4]
  assign _T_42216 = valid_63_10 ? 6'ha : _T_42215; // @[Mux.scala 31:69:@20540.4]
  assign _T_42217 = valid_63_9 ? 6'h9 : _T_42216; // @[Mux.scala 31:69:@20541.4]
  assign _T_42218 = valid_63_8 ? 6'h8 : _T_42217; // @[Mux.scala 31:69:@20542.4]
  assign _T_42219 = valid_63_7 ? 6'h7 : _T_42218; // @[Mux.scala 31:69:@20543.4]
  assign _T_42220 = valid_63_6 ? 6'h6 : _T_42219; // @[Mux.scala 31:69:@20544.4]
  assign _T_42221 = valid_63_5 ? 6'h5 : _T_42220; // @[Mux.scala 31:69:@20545.4]
  assign _T_42222 = valid_63_4 ? 6'h4 : _T_42221; // @[Mux.scala 31:69:@20546.4]
  assign _T_42223 = valid_63_3 ? 6'h3 : _T_42222; // @[Mux.scala 31:69:@20547.4]
  assign _T_42224 = valid_63_2 ? 6'h2 : _T_42223; // @[Mux.scala 31:69:@20548.4]
  assign _T_42225 = valid_63_1 ? 6'h1 : _T_42224; // @[Mux.scala 31:69:@20549.4]
  assign select_63 = valid_63_0 ? 6'h0 : _T_42225; // @[Mux.scala 31:69:@20550.4]
  assign _GEN_4033 = 6'h1 == select_63 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4034 = 6'h2 == select_63 ? io_inData_2 : _GEN_4033; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4035 = 6'h3 == select_63 ? io_inData_3 : _GEN_4034; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4036 = 6'h4 == select_63 ? io_inData_4 : _GEN_4035; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4037 = 6'h5 == select_63 ? io_inData_5 : _GEN_4036; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4038 = 6'h6 == select_63 ? io_inData_6 : _GEN_4037; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4039 = 6'h7 == select_63 ? io_inData_7 : _GEN_4038; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4040 = 6'h8 == select_63 ? io_inData_8 : _GEN_4039; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4041 = 6'h9 == select_63 ? io_inData_9 : _GEN_4040; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4042 = 6'ha == select_63 ? io_inData_10 : _GEN_4041; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4043 = 6'hb == select_63 ? io_inData_11 : _GEN_4042; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4044 = 6'hc == select_63 ? io_inData_12 : _GEN_4043; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4045 = 6'hd == select_63 ? io_inData_13 : _GEN_4044; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4046 = 6'he == select_63 ? io_inData_14 : _GEN_4045; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4047 = 6'hf == select_63 ? io_inData_15 : _GEN_4046; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4048 = 6'h10 == select_63 ? io_inData_16 : _GEN_4047; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4049 = 6'h11 == select_63 ? io_inData_17 : _GEN_4048; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4050 = 6'h12 == select_63 ? io_inData_18 : _GEN_4049; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4051 = 6'h13 == select_63 ? io_inData_19 : _GEN_4050; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4052 = 6'h14 == select_63 ? io_inData_20 : _GEN_4051; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4053 = 6'h15 == select_63 ? io_inData_21 : _GEN_4052; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4054 = 6'h16 == select_63 ? io_inData_22 : _GEN_4053; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4055 = 6'h17 == select_63 ? io_inData_23 : _GEN_4054; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4056 = 6'h18 == select_63 ? io_inData_24 : _GEN_4055; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4057 = 6'h19 == select_63 ? io_inData_25 : _GEN_4056; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4058 = 6'h1a == select_63 ? io_inData_26 : _GEN_4057; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4059 = 6'h1b == select_63 ? io_inData_27 : _GEN_4058; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4060 = 6'h1c == select_63 ? io_inData_28 : _GEN_4059; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4061 = 6'h1d == select_63 ? io_inData_29 : _GEN_4060; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4062 = 6'h1e == select_63 ? io_inData_30 : _GEN_4061; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4063 = 6'h1f == select_63 ? io_inData_31 : _GEN_4062; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4064 = 6'h20 == select_63 ? io_inData_32 : _GEN_4063; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4065 = 6'h21 == select_63 ? io_inData_33 : _GEN_4064; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4066 = 6'h22 == select_63 ? io_inData_34 : _GEN_4065; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4067 = 6'h23 == select_63 ? io_inData_35 : _GEN_4066; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4068 = 6'h24 == select_63 ? io_inData_36 : _GEN_4067; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4069 = 6'h25 == select_63 ? io_inData_37 : _GEN_4068; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4070 = 6'h26 == select_63 ? io_inData_38 : _GEN_4069; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4071 = 6'h27 == select_63 ? io_inData_39 : _GEN_4070; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4072 = 6'h28 == select_63 ? io_inData_40 : _GEN_4071; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4073 = 6'h29 == select_63 ? io_inData_41 : _GEN_4072; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4074 = 6'h2a == select_63 ? io_inData_42 : _GEN_4073; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4075 = 6'h2b == select_63 ? io_inData_43 : _GEN_4074; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4076 = 6'h2c == select_63 ? io_inData_44 : _GEN_4075; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4077 = 6'h2d == select_63 ? io_inData_45 : _GEN_4076; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4078 = 6'h2e == select_63 ? io_inData_46 : _GEN_4077; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4079 = 6'h2f == select_63 ? io_inData_47 : _GEN_4078; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4080 = 6'h30 == select_63 ? io_inData_48 : _GEN_4079; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4081 = 6'h31 == select_63 ? io_inData_49 : _GEN_4080; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4082 = 6'h32 == select_63 ? io_inData_50 : _GEN_4081; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4083 = 6'h33 == select_63 ? io_inData_51 : _GEN_4082; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4084 = 6'h34 == select_63 ? io_inData_52 : _GEN_4083; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4085 = 6'h35 == select_63 ? io_inData_53 : _GEN_4084; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4086 = 6'h36 == select_63 ? io_inData_54 : _GEN_4085; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4087 = 6'h37 == select_63 ? io_inData_55 : _GEN_4086; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4088 = 6'h38 == select_63 ? io_inData_56 : _GEN_4087; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4089 = 6'h39 == select_63 ? io_inData_57 : _GEN_4088; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4090 = 6'h3a == select_63 ? io_inData_58 : _GEN_4089; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4091 = 6'h3b == select_63 ? io_inData_59 : _GEN_4090; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4092 = 6'h3c == select_63 ? io_inData_60 : _GEN_4091; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4093 = 6'h3d == select_63 ? io_inData_61 : _GEN_4092; // @[Switch.scala 33:19:@20552.4]
  assign _GEN_4094 = 6'h3e == select_63 ? io_inData_62 : _GEN_4093; // @[Switch.scala 33:19:@20552.4]
  assign _T_42234 = {valid_63_7,valid_63_6,valid_63_5,valid_63_4,valid_63_3,valid_63_2,valid_63_1,valid_63_0}; // @[Switch.scala 34:32:@20559.4]
  assign _T_42242 = {valid_63_15,valid_63_14,valid_63_13,valid_63_12,valid_63_11,valid_63_10,valid_63_9,valid_63_8,_T_42234}; // @[Switch.scala 34:32:@20567.4]
  assign _T_42249 = {valid_63_23,valid_63_22,valid_63_21,valid_63_20,valid_63_19,valid_63_18,valid_63_17,valid_63_16}; // @[Switch.scala 34:32:@20574.4]
  assign _T_42258 = {valid_63_31,valid_63_30,valid_63_29,valid_63_28,valid_63_27,valid_63_26,valid_63_25,valid_63_24,_T_42249,_T_42242}; // @[Switch.scala 34:32:@20583.4]
  assign _T_42265 = {valid_63_39,valid_63_38,valid_63_37,valid_63_36,valid_63_35,valid_63_34,valid_63_33,valid_63_32}; // @[Switch.scala 34:32:@20590.4]
  assign _T_42273 = {valid_63_47,valid_63_46,valid_63_45,valid_63_44,valid_63_43,valid_63_42,valid_63_41,valid_63_40,_T_42265}; // @[Switch.scala 34:32:@20598.4]
  assign _T_42280 = {valid_63_55,valid_63_54,valid_63_53,valid_63_52,valid_63_51,valid_63_50,valid_63_49,valid_63_48}; // @[Switch.scala 34:32:@20605.4]
  assign _T_42289 = {valid_63_63,valid_63_62,valid_63_61,valid_63_60,valid_63_59,valid_63_58,valid_63_57,valid_63_56,_T_42280,_T_42273}; // @[Switch.scala 34:32:@20614.4]
  assign _T_42290 = {_T_42289,_T_42258}; // @[Switch.scala 34:32:@20615.4]
  assign _T_59460 = select_0 == 6'h0; // @[Switch.scala 41:52:@20619.4]
  assign output_0_0 = io_outValid_0 & _T_59460; // @[Switch.scala 41:38:@20620.4]
  assign _T_59463 = select_1 == 6'h0; // @[Switch.scala 41:52:@20622.4]
  assign output_0_1 = io_outValid_1 & _T_59463; // @[Switch.scala 41:38:@20623.4]
  assign _T_59466 = select_2 == 6'h0; // @[Switch.scala 41:52:@20625.4]
  assign output_0_2 = io_outValid_2 & _T_59466; // @[Switch.scala 41:38:@20626.4]
  assign _T_59469 = select_3 == 6'h0; // @[Switch.scala 41:52:@20628.4]
  assign output_0_3 = io_outValid_3 & _T_59469; // @[Switch.scala 41:38:@20629.4]
  assign _T_59472 = select_4 == 6'h0; // @[Switch.scala 41:52:@20631.4]
  assign output_0_4 = io_outValid_4 & _T_59472; // @[Switch.scala 41:38:@20632.4]
  assign _T_59475 = select_5 == 6'h0; // @[Switch.scala 41:52:@20634.4]
  assign output_0_5 = io_outValid_5 & _T_59475; // @[Switch.scala 41:38:@20635.4]
  assign _T_59478 = select_6 == 6'h0; // @[Switch.scala 41:52:@20637.4]
  assign output_0_6 = io_outValid_6 & _T_59478; // @[Switch.scala 41:38:@20638.4]
  assign _T_59481 = select_7 == 6'h0; // @[Switch.scala 41:52:@20640.4]
  assign output_0_7 = io_outValid_7 & _T_59481; // @[Switch.scala 41:38:@20641.4]
  assign _T_59484 = select_8 == 6'h0; // @[Switch.scala 41:52:@20643.4]
  assign output_0_8 = io_outValid_8 & _T_59484; // @[Switch.scala 41:38:@20644.4]
  assign _T_59487 = select_9 == 6'h0; // @[Switch.scala 41:52:@20646.4]
  assign output_0_9 = io_outValid_9 & _T_59487; // @[Switch.scala 41:38:@20647.4]
  assign _T_59490 = select_10 == 6'h0; // @[Switch.scala 41:52:@20649.4]
  assign output_0_10 = io_outValid_10 & _T_59490; // @[Switch.scala 41:38:@20650.4]
  assign _T_59493 = select_11 == 6'h0; // @[Switch.scala 41:52:@20652.4]
  assign output_0_11 = io_outValid_11 & _T_59493; // @[Switch.scala 41:38:@20653.4]
  assign _T_59496 = select_12 == 6'h0; // @[Switch.scala 41:52:@20655.4]
  assign output_0_12 = io_outValid_12 & _T_59496; // @[Switch.scala 41:38:@20656.4]
  assign _T_59499 = select_13 == 6'h0; // @[Switch.scala 41:52:@20658.4]
  assign output_0_13 = io_outValid_13 & _T_59499; // @[Switch.scala 41:38:@20659.4]
  assign _T_59502 = select_14 == 6'h0; // @[Switch.scala 41:52:@20661.4]
  assign output_0_14 = io_outValid_14 & _T_59502; // @[Switch.scala 41:38:@20662.4]
  assign _T_59505 = select_15 == 6'h0; // @[Switch.scala 41:52:@20664.4]
  assign output_0_15 = io_outValid_15 & _T_59505; // @[Switch.scala 41:38:@20665.4]
  assign _T_59508 = select_16 == 6'h0; // @[Switch.scala 41:52:@20667.4]
  assign output_0_16 = io_outValid_16 & _T_59508; // @[Switch.scala 41:38:@20668.4]
  assign _T_59511 = select_17 == 6'h0; // @[Switch.scala 41:52:@20670.4]
  assign output_0_17 = io_outValid_17 & _T_59511; // @[Switch.scala 41:38:@20671.4]
  assign _T_59514 = select_18 == 6'h0; // @[Switch.scala 41:52:@20673.4]
  assign output_0_18 = io_outValid_18 & _T_59514; // @[Switch.scala 41:38:@20674.4]
  assign _T_59517 = select_19 == 6'h0; // @[Switch.scala 41:52:@20676.4]
  assign output_0_19 = io_outValid_19 & _T_59517; // @[Switch.scala 41:38:@20677.4]
  assign _T_59520 = select_20 == 6'h0; // @[Switch.scala 41:52:@20679.4]
  assign output_0_20 = io_outValid_20 & _T_59520; // @[Switch.scala 41:38:@20680.4]
  assign _T_59523 = select_21 == 6'h0; // @[Switch.scala 41:52:@20682.4]
  assign output_0_21 = io_outValid_21 & _T_59523; // @[Switch.scala 41:38:@20683.4]
  assign _T_59526 = select_22 == 6'h0; // @[Switch.scala 41:52:@20685.4]
  assign output_0_22 = io_outValid_22 & _T_59526; // @[Switch.scala 41:38:@20686.4]
  assign _T_59529 = select_23 == 6'h0; // @[Switch.scala 41:52:@20688.4]
  assign output_0_23 = io_outValid_23 & _T_59529; // @[Switch.scala 41:38:@20689.4]
  assign _T_59532 = select_24 == 6'h0; // @[Switch.scala 41:52:@20691.4]
  assign output_0_24 = io_outValid_24 & _T_59532; // @[Switch.scala 41:38:@20692.4]
  assign _T_59535 = select_25 == 6'h0; // @[Switch.scala 41:52:@20694.4]
  assign output_0_25 = io_outValid_25 & _T_59535; // @[Switch.scala 41:38:@20695.4]
  assign _T_59538 = select_26 == 6'h0; // @[Switch.scala 41:52:@20697.4]
  assign output_0_26 = io_outValid_26 & _T_59538; // @[Switch.scala 41:38:@20698.4]
  assign _T_59541 = select_27 == 6'h0; // @[Switch.scala 41:52:@20700.4]
  assign output_0_27 = io_outValid_27 & _T_59541; // @[Switch.scala 41:38:@20701.4]
  assign _T_59544 = select_28 == 6'h0; // @[Switch.scala 41:52:@20703.4]
  assign output_0_28 = io_outValid_28 & _T_59544; // @[Switch.scala 41:38:@20704.4]
  assign _T_59547 = select_29 == 6'h0; // @[Switch.scala 41:52:@20706.4]
  assign output_0_29 = io_outValid_29 & _T_59547; // @[Switch.scala 41:38:@20707.4]
  assign _T_59550 = select_30 == 6'h0; // @[Switch.scala 41:52:@20709.4]
  assign output_0_30 = io_outValid_30 & _T_59550; // @[Switch.scala 41:38:@20710.4]
  assign _T_59553 = select_31 == 6'h0; // @[Switch.scala 41:52:@20712.4]
  assign output_0_31 = io_outValid_31 & _T_59553; // @[Switch.scala 41:38:@20713.4]
  assign _T_59556 = select_32 == 6'h0; // @[Switch.scala 41:52:@20715.4]
  assign output_0_32 = io_outValid_32 & _T_59556; // @[Switch.scala 41:38:@20716.4]
  assign _T_59559 = select_33 == 6'h0; // @[Switch.scala 41:52:@20718.4]
  assign output_0_33 = io_outValid_33 & _T_59559; // @[Switch.scala 41:38:@20719.4]
  assign _T_59562 = select_34 == 6'h0; // @[Switch.scala 41:52:@20721.4]
  assign output_0_34 = io_outValid_34 & _T_59562; // @[Switch.scala 41:38:@20722.4]
  assign _T_59565 = select_35 == 6'h0; // @[Switch.scala 41:52:@20724.4]
  assign output_0_35 = io_outValid_35 & _T_59565; // @[Switch.scala 41:38:@20725.4]
  assign _T_59568 = select_36 == 6'h0; // @[Switch.scala 41:52:@20727.4]
  assign output_0_36 = io_outValid_36 & _T_59568; // @[Switch.scala 41:38:@20728.4]
  assign _T_59571 = select_37 == 6'h0; // @[Switch.scala 41:52:@20730.4]
  assign output_0_37 = io_outValid_37 & _T_59571; // @[Switch.scala 41:38:@20731.4]
  assign _T_59574 = select_38 == 6'h0; // @[Switch.scala 41:52:@20733.4]
  assign output_0_38 = io_outValid_38 & _T_59574; // @[Switch.scala 41:38:@20734.4]
  assign _T_59577 = select_39 == 6'h0; // @[Switch.scala 41:52:@20736.4]
  assign output_0_39 = io_outValid_39 & _T_59577; // @[Switch.scala 41:38:@20737.4]
  assign _T_59580 = select_40 == 6'h0; // @[Switch.scala 41:52:@20739.4]
  assign output_0_40 = io_outValid_40 & _T_59580; // @[Switch.scala 41:38:@20740.4]
  assign _T_59583 = select_41 == 6'h0; // @[Switch.scala 41:52:@20742.4]
  assign output_0_41 = io_outValid_41 & _T_59583; // @[Switch.scala 41:38:@20743.4]
  assign _T_59586 = select_42 == 6'h0; // @[Switch.scala 41:52:@20745.4]
  assign output_0_42 = io_outValid_42 & _T_59586; // @[Switch.scala 41:38:@20746.4]
  assign _T_59589 = select_43 == 6'h0; // @[Switch.scala 41:52:@20748.4]
  assign output_0_43 = io_outValid_43 & _T_59589; // @[Switch.scala 41:38:@20749.4]
  assign _T_59592 = select_44 == 6'h0; // @[Switch.scala 41:52:@20751.4]
  assign output_0_44 = io_outValid_44 & _T_59592; // @[Switch.scala 41:38:@20752.4]
  assign _T_59595 = select_45 == 6'h0; // @[Switch.scala 41:52:@20754.4]
  assign output_0_45 = io_outValid_45 & _T_59595; // @[Switch.scala 41:38:@20755.4]
  assign _T_59598 = select_46 == 6'h0; // @[Switch.scala 41:52:@20757.4]
  assign output_0_46 = io_outValid_46 & _T_59598; // @[Switch.scala 41:38:@20758.4]
  assign _T_59601 = select_47 == 6'h0; // @[Switch.scala 41:52:@20760.4]
  assign output_0_47 = io_outValid_47 & _T_59601; // @[Switch.scala 41:38:@20761.4]
  assign _T_59604 = select_48 == 6'h0; // @[Switch.scala 41:52:@20763.4]
  assign output_0_48 = io_outValid_48 & _T_59604; // @[Switch.scala 41:38:@20764.4]
  assign _T_59607 = select_49 == 6'h0; // @[Switch.scala 41:52:@20766.4]
  assign output_0_49 = io_outValid_49 & _T_59607; // @[Switch.scala 41:38:@20767.4]
  assign _T_59610 = select_50 == 6'h0; // @[Switch.scala 41:52:@20769.4]
  assign output_0_50 = io_outValid_50 & _T_59610; // @[Switch.scala 41:38:@20770.4]
  assign _T_59613 = select_51 == 6'h0; // @[Switch.scala 41:52:@20772.4]
  assign output_0_51 = io_outValid_51 & _T_59613; // @[Switch.scala 41:38:@20773.4]
  assign _T_59616 = select_52 == 6'h0; // @[Switch.scala 41:52:@20775.4]
  assign output_0_52 = io_outValid_52 & _T_59616; // @[Switch.scala 41:38:@20776.4]
  assign _T_59619 = select_53 == 6'h0; // @[Switch.scala 41:52:@20778.4]
  assign output_0_53 = io_outValid_53 & _T_59619; // @[Switch.scala 41:38:@20779.4]
  assign _T_59622 = select_54 == 6'h0; // @[Switch.scala 41:52:@20781.4]
  assign output_0_54 = io_outValid_54 & _T_59622; // @[Switch.scala 41:38:@20782.4]
  assign _T_59625 = select_55 == 6'h0; // @[Switch.scala 41:52:@20784.4]
  assign output_0_55 = io_outValid_55 & _T_59625; // @[Switch.scala 41:38:@20785.4]
  assign _T_59628 = select_56 == 6'h0; // @[Switch.scala 41:52:@20787.4]
  assign output_0_56 = io_outValid_56 & _T_59628; // @[Switch.scala 41:38:@20788.4]
  assign _T_59631 = select_57 == 6'h0; // @[Switch.scala 41:52:@20790.4]
  assign output_0_57 = io_outValid_57 & _T_59631; // @[Switch.scala 41:38:@20791.4]
  assign _T_59634 = select_58 == 6'h0; // @[Switch.scala 41:52:@20793.4]
  assign output_0_58 = io_outValid_58 & _T_59634; // @[Switch.scala 41:38:@20794.4]
  assign _T_59637 = select_59 == 6'h0; // @[Switch.scala 41:52:@20796.4]
  assign output_0_59 = io_outValid_59 & _T_59637; // @[Switch.scala 41:38:@20797.4]
  assign _T_59640 = select_60 == 6'h0; // @[Switch.scala 41:52:@20799.4]
  assign output_0_60 = io_outValid_60 & _T_59640; // @[Switch.scala 41:38:@20800.4]
  assign _T_59643 = select_61 == 6'h0; // @[Switch.scala 41:52:@20802.4]
  assign output_0_61 = io_outValid_61 & _T_59643; // @[Switch.scala 41:38:@20803.4]
  assign _T_59646 = select_62 == 6'h0; // @[Switch.scala 41:52:@20805.4]
  assign output_0_62 = io_outValid_62 & _T_59646; // @[Switch.scala 41:38:@20806.4]
  assign _T_59649 = select_63 == 6'h0; // @[Switch.scala 41:52:@20808.4]
  assign output_0_63 = io_outValid_63 & _T_59649; // @[Switch.scala 41:38:@20809.4]
  assign _T_59657 = {output_0_7,output_0_6,output_0_5,output_0_4,output_0_3,output_0_2,output_0_1,output_0_0}; // @[Switch.scala 43:31:@20817.4]
  assign _T_59665 = {output_0_15,output_0_14,output_0_13,output_0_12,output_0_11,output_0_10,output_0_9,output_0_8,_T_59657}; // @[Switch.scala 43:31:@20825.4]
  assign _T_59672 = {output_0_23,output_0_22,output_0_21,output_0_20,output_0_19,output_0_18,output_0_17,output_0_16}; // @[Switch.scala 43:31:@20832.4]
  assign _T_59681 = {output_0_31,output_0_30,output_0_29,output_0_28,output_0_27,output_0_26,output_0_25,output_0_24,_T_59672,_T_59665}; // @[Switch.scala 43:31:@20841.4]
  assign _T_59688 = {output_0_39,output_0_38,output_0_37,output_0_36,output_0_35,output_0_34,output_0_33,output_0_32}; // @[Switch.scala 43:31:@20848.4]
  assign _T_59696 = {output_0_47,output_0_46,output_0_45,output_0_44,output_0_43,output_0_42,output_0_41,output_0_40,_T_59688}; // @[Switch.scala 43:31:@20856.4]
  assign _T_59703 = {output_0_55,output_0_54,output_0_53,output_0_52,output_0_51,output_0_50,output_0_49,output_0_48}; // @[Switch.scala 43:31:@20863.4]
  assign _T_59712 = {output_0_63,output_0_62,output_0_61,output_0_60,output_0_59,output_0_58,output_0_57,output_0_56,_T_59703,_T_59696}; // @[Switch.scala 43:31:@20872.4]
  assign _T_59713 = {_T_59712,_T_59681}; // @[Switch.scala 43:31:@20873.4]
  assign _T_59717 = select_0 == 6'h1; // @[Switch.scala 41:52:@20876.4]
  assign output_1_0 = io_outValid_0 & _T_59717; // @[Switch.scala 41:38:@20877.4]
  assign _T_59720 = select_1 == 6'h1; // @[Switch.scala 41:52:@20879.4]
  assign output_1_1 = io_outValid_1 & _T_59720; // @[Switch.scala 41:38:@20880.4]
  assign _T_59723 = select_2 == 6'h1; // @[Switch.scala 41:52:@20882.4]
  assign output_1_2 = io_outValid_2 & _T_59723; // @[Switch.scala 41:38:@20883.4]
  assign _T_59726 = select_3 == 6'h1; // @[Switch.scala 41:52:@20885.4]
  assign output_1_3 = io_outValid_3 & _T_59726; // @[Switch.scala 41:38:@20886.4]
  assign _T_59729 = select_4 == 6'h1; // @[Switch.scala 41:52:@20888.4]
  assign output_1_4 = io_outValid_4 & _T_59729; // @[Switch.scala 41:38:@20889.4]
  assign _T_59732 = select_5 == 6'h1; // @[Switch.scala 41:52:@20891.4]
  assign output_1_5 = io_outValid_5 & _T_59732; // @[Switch.scala 41:38:@20892.4]
  assign _T_59735 = select_6 == 6'h1; // @[Switch.scala 41:52:@20894.4]
  assign output_1_6 = io_outValid_6 & _T_59735; // @[Switch.scala 41:38:@20895.4]
  assign _T_59738 = select_7 == 6'h1; // @[Switch.scala 41:52:@20897.4]
  assign output_1_7 = io_outValid_7 & _T_59738; // @[Switch.scala 41:38:@20898.4]
  assign _T_59741 = select_8 == 6'h1; // @[Switch.scala 41:52:@20900.4]
  assign output_1_8 = io_outValid_8 & _T_59741; // @[Switch.scala 41:38:@20901.4]
  assign _T_59744 = select_9 == 6'h1; // @[Switch.scala 41:52:@20903.4]
  assign output_1_9 = io_outValid_9 & _T_59744; // @[Switch.scala 41:38:@20904.4]
  assign _T_59747 = select_10 == 6'h1; // @[Switch.scala 41:52:@20906.4]
  assign output_1_10 = io_outValid_10 & _T_59747; // @[Switch.scala 41:38:@20907.4]
  assign _T_59750 = select_11 == 6'h1; // @[Switch.scala 41:52:@20909.4]
  assign output_1_11 = io_outValid_11 & _T_59750; // @[Switch.scala 41:38:@20910.4]
  assign _T_59753 = select_12 == 6'h1; // @[Switch.scala 41:52:@20912.4]
  assign output_1_12 = io_outValid_12 & _T_59753; // @[Switch.scala 41:38:@20913.4]
  assign _T_59756 = select_13 == 6'h1; // @[Switch.scala 41:52:@20915.4]
  assign output_1_13 = io_outValid_13 & _T_59756; // @[Switch.scala 41:38:@20916.4]
  assign _T_59759 = select_14 == 6'h1; // @[Switch.scala 41:52:@20918.4]
  assign output_1_14 = io_outValid_14 & _T_59759; // @[Switch.scala 41:38:@20919.4]
  assign _T_59762 = select_15 == 6'h1; // @[Switch.scala 41:52:@20921.4]
  assign output_1_15 = io_outValid_15 & _T_59762; // @[Switch.scala 41:38:@20922.4]
  assign _T_59765 = select_16 == 6'h1; // @[Switch.scala 41:52:@20924.4]
  assign output_1_16 = io_outValid_16 & _T_59765; // @[Switch.scala 41:38:@20925.4]
  assign _T_59768 = select_17 == 6'h1; // @[Switch.scala 41:52:@20927.4]
  assign output_1_17 = io_outValid_17 & _T_59768; // @[Switch.scala 41:38:@20928.4]
  assign _T_59771 = select_18 == 6'h1; // @[Switch.scala 41:52:@20930.4]
  assign output_1_18 = io_outValid_18 & _T_59771; // @[Switch.scala 41:38:@20931.4]
  assign _T_59774 = select_19 == 6'h1; // @[Switch.scala 41:52:@20933.4]
  assign output_1_19 = io_outValid_19 & _T_59774; // @[Switch.scala 41:38:@20934.4]
  assign _T_59777 = select_20 == 6'h1; // @[Switch.scala 41:52:@20936.4]
  assign output_1_20 = io_outValid_20 & _T_59777; // @[Switch.scala 41:38:@20937.4]
  assign _T_59780 = select_21 == 6'h1; // @[Switch.scala 41:52:@20939.4]
  assign output_1_21 = io_outValid_21 & _T_59780; // @[Switch.scala 41:38:@20940.4]
  assign _T_59783 = select_22 == 6'h1; // @[Switch.scala 41:52:@20942.4]
  assign output_1_22 = io_outValid_22 & _T_59783; // @[Switch.scala 41:38:@20943.4]
  assign _T_59786 = select_23 == 6'h1; // @[Switch.scala 41:52:@20945.4]
  assign output_1_23 = io_outValid_23 & _T_59786; // @[Switch.scala 41:38:@20946.4]
  assign _T_59789 = select_24 == 6'h1; // @[Switch.scala 41:52:@20948.4]
  assign output_1_24 = io_outValid_24 & _T_59789; // @[Switch.scala 41:38:@20949.4]
  assign _T_59792 = select_25 == 6'h1; // @[Switch.scala 41:52:@20951.4]
  assign output_1_25 = io_outValid_25 & _T_59792; // @[Switch.scala 41:38:@20952.4]
  assign _T_59795 = select_26 == 6'h1; // @[Switch.scala 41:52:@20954.4]
  assign output_1_26 = io_outValid_26 & _T_59795; // @[Switch.scala 41:38:@20955.4]
  assign _T_59798 = select_27 == 6'h1; // @[Switch.scala 41:52:@20957.4]
  assign output_1_27 = io_outValid_27 & _T_59798; // @[Switch.scala 41:38:@20958.4]
  assign _T_59801 = select_28 == 6'h1; // @[Switch.scala 41:52:@20960.4]
  assign output_1_28 = io_outValid_28 & _T_59801; // @[Switch.scala 41:38:@20961.4]
  assign _T_59804 = select_29 == 6'h1; // @[Switch.scala 41:52:@20963.4]
  assign output_1_29 = io_outValid_29 & _T_59804; // @[Switch.scala 41:38:@20964.4]
  assign _T_59807 = select_30 == 6'h1; // @[Switch.scala 41:52:@20966.4]
  assign output_1_30 = io_outValid_30 & _T_59807; // @[Switch.scala 41:38:@20967.4]
  assign _T_59810 = select_31 == 6'h1; // @[Switch.scala 41:52:@20969.4]
  assign output_1_31 = io_outValid_31 & _T_59810; // @[Switch.scala 41:38:@20970.4]
  assign _T_59813 = select_32 == 6'h1; // @[Switch.scala 41:52:@20972.4]
  assign output_1_32 = io_outValid_32 & _T_59813; // @[Switch.scala 41:38:@20973.4]
  assign _T_59816 = select_33 == 6'h1; // @[Switch.scala 41:52:@20975.4]
  assign output_1_33 = io_outValid_33 & _T_59816; // @[Switch.scala 41:38:@20976.4]
  assign _T_59819 = select_34 == 6'h1; // @[Switch.scala 41:52:@20978.4]
  assign output_1_34 = io_outValid_34 & _T_59819; // @[Switch.scala 41:38:@20979.4]
  assign _T_59822 = select_35 == 6'h1; // @[Switch.scala 41:52:@20981.4]
  assign output_1_35 = io_outValid_35 & _T_59822; // @[Switch.scala 41:38:@20982.4]
  assign _T_59825 = select_36 == 6'h1; // @[Switch.scala 41:52:@20984.4]
  assign output_1_36 = io_outValid_36 & _T_59825; // @[Switch.scala 41:38:@20985.4]
  assign _T_59828 = select_37 == 6'h1; // @[Switch.scala 41:52:@20987.4]
  assign output_1_37 = io_outValid_37 & _T_59828; // @[Switch.scala 41:38:@20988.4]
  assign _T_59831 = select_38 == 6'h1; // @[Switch.scala 41:52:@20990.4]
  assign output_1_38 = io_outValid_38 & _T_59831; // @[Switch.scala 41:38:@20991.4]
  assign _T_59834 = select_39 == 6'h1; // @[Switch.scala 41:52:@20993.4]
  assign output_1_39 = io_outValid_39 & _T_59834; // @[Switch.scala 41:38:@20994.4]
  assign _T_59837 = select_40 == 6'h1; // @[Switch.scala 41:52:@20996.4]
  assign output_1_40 = io_outValid_40 & _T_59837; // @[Switch.scala 41:38:@20997.4]
  assign _T_59840 = select_41 == 6'h1; // @[Switch.scala 41:52:@20999.4]
  assign output_1_41 = io_outValid_41 & _T_59840; // @[Switch.scala 41:38:@21000.4]
  assign _T_59843 = select_42 == 6'h1; // @[Switch.scala 41:52:@21002.4]
  assign output_1_42 = io_outValid_42 & _T_59843; // @[Switch.scala 41:38:@21003.4]
  assign _T_59846 = select_43 == 6'h1; // @[Switch.scala 41:52:@21005.4]
  assign output_1_43 = io_outValid_43 & _T_59846; // @[Switch.scala 41:38:@21006.4]
  assign _T_59849 = select_44 == 6'h1; // @[Switch.scala 41:52:@21008.4]
  assign output_1_44 = io_outValid_44 & _T_59849; // @[Switch.scala 41:38:@21009.4]
  assign _T_59852 = select_45 == 6'h1; // @[Switch.scala 41:52:@21011.4]
  assign output_1_45 = io_outValid_45 & _T_59852; // @[Switch.scala 41:38:@21012.4]
  assign _T_59855 = select_46 == 6'h1; // @[Switch.scala 41:52:@21014.4]
  assign output_1_46 = io_outValid_46 & _T_59855; // @[Switch.scala 41:38:@21015.4]
  assign _T_59858 = select_47 == 6'h1; // @[Switch.scala 41:52:@21017.4]
  assign output_1_47 = io_outValid_47 & _T_59858; // @[Switch.scala 41:38:@21018.4]
  assign _T_59861 = select_48 == 6'h1; // @[Switch.scala 41:52:@21020.4]
  assign output_1_48 = io_outValid_48 & _T_59861; // @[Switch.scala 41:38:@21021.4]
  assign _T_59864 = select_49 == 6'h1; // @[Switch.scala 41:52:@21023.4]
  assign output_1_49 = io_outValid_49 & _T_59864; // @[Switch.scala 41:38:@21024.4]
  assign _T_59867 = select_50 == 6'h1; // @[Switch.scala 41:52:@21026.4]
  assign output_1_50 = io_outValid_50 & _T_59867; // @[Switch.scala 41:38:@21027.4]
  assign _T_59870 = select_51 == 6'h1; // @[Switch.scala 41:52:@21029.4]
  assign output_1_51 = io_outValid_51 & _T_59870; // @[Switch.scala 41:38:@21030.4]
  assign _T_59873 = select_52 == 6'h1; // @[Switch.scala 41:52:@21032.4]
  assign output_1_52 = io_outValid_52 & _T_59873; // @[Switch.scala 41:38:@21033.4]
  assign _T_59876 = select_53 == 6'h1; // @[Switch.scala 41:52:@21035.4]
  assign output_1_53 = io_outValid_53 & _T_59876; // @[Switch.scala 41:38:@21036.4]
  assign _T_59879 = select_54 == 6'h1; // @[Switch.scala 41:52:@21038.4]
  assign output_1_54 = io_outValid_54 & _T_59879; // @[Switch.scala 41:38:@21039.4]
  assign _T_59882 = select_55 == 6'h1; // @[Switch.scala 41:52:@21041.4]
  assign output_1_55 = io_outValid_55 & _T_59882; // @[Switch.scala 41:38:@21042.4]
  assign _T_59885 = select_56 == 6'h1; // @[Switch.scala 41:52:@21044.4]
  assign output_1_56 = io_outValid_56 & _T_59885; // @[Switch.scala 41:38:@21045.4]
  assign _T_59888 = select_57 == 6'h1; // @[Switch.scala 41:52:@21047.4]
  assign output_1_57 = io_outValid_57 & _T_59888; // @[Switch.scala 41:38:@21048.4]
  assign _T_59891 = select_58 == 6'h1; // @[Switch.scala 41:52:@21050.4]
  assign output_1_58 = io_outValid_58 & _T_59891; // @[Switch.scala 41:38:@21051.4]
  assign _T_59894 = select_59 == 6'h1; // @[Switch.scala 41:52:@21053.4]
  assign output_1_59 = io_outValid_59 & _T_59894; // @[Switch.scala 41:38:@21054.4]
  assign _T_59897 = select_60 == 6'h1; // @[Switch.scala 41:52:@21056.4]
  assign output_1_60 = io_outValid_60 & _T_59897; // @[Switch.scala 41:38:@21057.4]
  assign _T_59900 = select_61 == 6'h1; // @[Switch.scala 41:52:@21059.4]
  assign output_1_61 = io_outValid_61 & _T_59900; // @[Switch.scala 41:38:@21060.4]
  assign _T_59903 = select_62 == 6'h1; // @[Switch.scala 41:52:@21062.4]
  assign output_1_62 = io_outValid_62 & _T_59903; // @[Switch.scala 41:38:@21063.4]
  assign _T_59906 = select_63 == 6'h1; // @[Switch.scala 41:52:@21065.4]
  assign output_1_63 = io_outValid_63 & _T_59906; // @[Switch.scala 41:38:@21066.4]
  assign _T_59914 = {output_1_7,output_1_6,output_1_5,output_1_4,output_1_3,output_1_2,output_1_1,output_1_0}; // @[Switch.scala 43:31:@21074.4]
  assign _T_59922 = {output_1_15,output_1_14,output_1_13,output_1_12,output_1_11,output_1_10,output_1_9,output_1_8,_T_59914}; // @[Switch.scala 43:31:@21082.4]
  assign _T_59929 = {output_1_23,output_1_22,output_1_21,output_1_20,output_1_19,output_1_18,output_1_17,output_1_16}; // @[Switch.scala 43:31:@21089.4]
  assign _T_59938 = {output_1_31,output_1_30,output_1_29,output_1_28,output_1_27,output_1_26,output_1_25,output_1_24,_T_59929,_T_59922}; // @[Switch.scala 43:31:@21098.4]
  assign _T_59945 = {output_1_39,output_1_38,output_1_37,output_1_36,output_1_35,output_1_34,output_1_33,output_1_32}; // @[Switch.scala 43:31:@21105.4]
  assign _T_59953 = {output_1_47,output_1_46,output_1_45,output_1_44,output_1_43,output_1_42,output_1_41,output_1_40,_T_59945}; // @[Switch.scala 43:31:@21113.4]
  assign _T_59960 = {output_1_55,output_1_54,output_1_53,output_1_52,output_1_51,output_1_50,output_1_49,output_1_48}; // @[Switch.scala 43:31:@21120.4]
  assign _T_59969 = {output_1_63,output_1_62,output_1_61,output_1_60,output_1_59,output_1_58,output_1_57,output_1_56,_T_59960,_T_59953}; // @[Switch.scala 43:31:@21129.4]
  assign _T_59970 = {_T_59969,_T_59938}; // @[Switch.scala 43:31:@21130.4]
  assign _T_59974 = select_0 == 6'h2; // @[Switch.scala 41:52:@21133.4]
  assign output_2_0 = io_outValid_0 & _T_59974; // @[Switch.scala 41:38:@21134.4]
  assign _T_59977 = select_1 == 6'h2; // @[Switch.scala 41:52:@21136.4]
  assign output_2_1 = io_outValid_1 & _T_59977; // @[Switch.scala 41:38:@21137.4]
  assign _T_59980 = select_2 == 6'h2; // @[Switch.scala 41:52:@21139.4]
  assign output_2_2 = io_outValid_2 & _T_59980; // @[Switch.scala 41:38:@21140.4]
  assign _T_59983 = select_3 == 6'h2; // @[Switch.scala 41:52:@21142.4]
  assign output_2_3 = io_outValid_3 & _T_59983; // @[Switch.scala 41:38:@21143.4]
  assign _T_59986 = select_4 == 6'h2; // @[Switch.scala 41:52:@21145.4]
  assign output_2_4 = io_outValid_4 & _T_59986; // @[Switch.scala 41:38:@21146.4]
  assign _T_59989 = select_5 == 6'h2; // @[Switch.scala 41:52:@21148.4]
  assign output_2_5 = io_outValid_5 & _T_59989; // @[Switch.scala 41:38:@21149.4]
  assign _T_59992 = select_6 == 6'h2; // @[Switch.scala 41:52:@21151.4]
  assign output_2_6 = io_outValid_6 & _T_59992; // @[Switch.scala 41:38:@21152.4]
  assign _T_59995 = select_7 == 6'h2; // @[Switch.scala 41:52:@21154.4]
  assign output_2_7 = io_outValid_7 & _T_59995; // @[Switch.scala 41:38:@21155.4]
  assign _T_59998 = select_8 == 6'h2; // @[Switch.scala 41:52:@21157.4]
  assign output_2_8 = io_outValid_8 & _T_59998; // @[Switch.scala 41:38:@21158.4]
  assign _T_60001 = select_9 == 6'h2; // @[Switch.scala 41:52:@21160.4]
  assign output_2_9 = io_outValid_9 & _T_60001; // @[Switch.scala 41:38:@21161.4]
  assign _T_60004 = select_10 == 6'h2; // @[Switch.scala 41:52:@21163.4]
  assign output_2_10 = io_outValid_10 & _T_60004; // @[Switch.scala 41:38:@21164.4]
  assign _T_60007 = select_11 == 6'h2; // @[Switch.scala 41:52:@21166.4]
  assign output_2_11 = io_outValid_11 & _T_60007; // @[Switch.scala 41:38:@21167.4]
  assign _T_60010 = select_12 == 6'h2; // @[Switch.scala 41:52:@21169.4]
  assign output_2_12 = io_outValid_12 & _T_60010; // @[Switch.scala 41:38:@21170.4]
  assign _T_60013 = select_13 == 6'h2; // @[Switch.scala 41:52:@21172.4]
  assign output_2_13 = io_outValid_13 & _T_60013; // @[Switch.scala 41:38:@21173.4]
  assign _T_60016 = select_14 == 6'h2; // @[Switch.scala 41:52:@21175.4]
  assign output_2_14 = io_outValid_14 & _T_60016; // @[Switch.scala 41:38:@21176.4]
  assign _T_60019 = select_15 == 6'h2; // @[Switch.scala 41:52:@21178.4]
  assign output_2_15 = io_outValid_15 & _T_60019; // @[Switch.scala 41:38:@21179.4]
  assign _T_60022 = select_16 == 6'h2; // @[Switch.scala 41:52:@21181.4]
  assign output_2_16 = io_outValid_16 & _T_60022; // @[Switch.scala 41:38:@21182.4]
  assign _T_60025 = select_17 == 6'h2; // @[Switch.scala 41:52:@21184.4]
  assign output_2_17 = io_outValid_17 & _T_60025; // @[Switch.scala 41:38:@21185.4]
  assign _T_60028 = select_18 == 6'h2; // @[Switch.scala 41:52:@21187.4]
  assign output_2_18 = io_outValid_18 & _T_60028; // @[Switch.scala 41:38:@21188.4]
  assign _T_60031 = select_19 == 6'h2; // @[Switch.scala 41:52:@21190.4]
  assign output_2_19 = io_outValid_19 & _T_60031; // @[Switch.scala 41:38:@21191.4]
  assign _T_60034 = select_20 == 6'h2; // @[Switch.scala 41:52:@21193.4]
  assign output_2_20 = io_outValid_20 & _T_60034; // @[Switch.scala 41:38:@21194.4]
  assign _T_60037 = select_21 == 6'h2; // @[Switch.scala 41:52:@21196.4]
  assign output_2_21 = io_outValid_21 & _T_60037; // @[Switch.scala 41:38:@21197.4]
  assign _T_60040 = select_22 == 6'h2; // @[Switch.scala 41:52:@21199.4]
  assign output_2_22 = io_outValid_22 & _T_60040; // @[Switch.scala 41:38:@21200.4]
  assign _T_60043 = select_23 == 6'h2; // @[Switch.scala 41:52:@21202.4]
  assign output_2_23 = io_outValid_23 & _T_60043; // @[Switch.scala 41:38:@21203.4]
  assign _T_60046 = select_24 == 6'h2; // @[Switch.scala 41:52:@21205.4]
  assign output_2_24 = io_outValid_24 & _T_60046; // @[Switch.scala 41:38:@21206.4]
  assign _T_60049 = select_25 == 6'h2; // @[Switch.scala 41:52:@21208.4]
  assign output_2_25 = io_outValid_25 & _T_60049; // @[Switch.scala 41:38:@21209.4]
  assign _T_60052 = select_26 == 6'h2; // @[Switch.scala 41:52:@21211.4]
  assign output_2_26 = io_outValid_26 & _T_60052; // @[Switch.scala 41:38:@21212.4]
  assign _T_60055 = select_27 == 6'h2; // @[Switch.scala 41:52:@21214.4]
  assign output_2_27 = io_outValid_27 & _T_60055; // @[Switch.scala 41:38:@21215.4]
  assign _T_60058 = select_28 == 6'h2; // @[Switch.scala 41:52:@21217.4]
  assign output_2_28 = io_outValid_28 & _T_60058; // @[Switch.scala 41:38:@21218.4]
  assign _T_60061 = select_29 == 6'h2; // @[Switch.scala 41:52:@21220.4]
  assign output_2_29 = io_outValid_29 & _T_60061; // @[Switch.scala 41:38:@21221.4]
  assign _T_60064 = select_30 == 6'h2; // @[Switch.scala 41:52:@21223.4]
  assign output_2_30 = io_outValid_30 & _T_60064; // @[Switch.scala 41:38:@21224.4]
  assign _T_60067 = select_31 == 6'h2; // @[Switch.scala 41:52:@21226.4]
  assign output_2_31 = io_outValid_31 & _T_60067; // @[Switch.scala 41:38:@21227.4]
  assign _T_60070 = select_32 == 6'h2; // @[Switch.scala 41:52:@21229.4]
  assign output_2_32 = io_outValid_32 & _T_60070; // @[Switch.scala 41:38:@21230.4]
  assign _T_60073 = select_33 == 6'h2; // @[Switch.scala 41:52:@21232.4]
  assign output_2_33 = io_outValid_33 & _T_60073; // @[Switch.scala 41:38:@21233.4]
  assign _T_60076 = select_34 == 6'h2; // @[Switch.scala 41:52:@21235.4]
  assign output_2_34 = io_outValid_34 & _T_60076; // @[Switch.scala 41:38:@21236.4]
  assign _T_60079 = select_35 == 6'h2; // @[Switch.scala 41:52:@21238.4]
  assign output_2_35 = io_outValid_35 & _T_60079; // @[Switch.scala 41:38:@21239.4]
  assign _T_60082 = select_36 == 6'h2; // @[Switch.scala 41:52:@21241.4]
  assign output_2_36 = io_outValid_36 & _T_60082; // @[Switch.scala 41:38:@21242.4]
  assign _T_60085 = select_37 == 6'h2; // @[Switch.scala 41:52:@21244.4]
  assign output_2_37 = io_outValid_37 & _T_60085; // @[Switch.scala 41:38:@21245.4]
  assign _T_60088 = select_38 == 6'h2; // @[Switch.scala 41:52:@21247.4]
  assign output_2_38 = io_outValid_38 & _T_60088; // @[Switch.scala 41:38:@21248.4]
  assign _T_60091 = select_39 == 6'h2; // @[Switch.scala 41:52:@21250.4]
  assign output_2_39 = io_outValid_39 & _T_60091; // @[Switch.scala 41:38:@21251.4]
  assign _T_60094 = select_40 == 6'h2; // @[Switch.scala 41:52:@21253.4]
  assign output_2_40 = io_outValid_40 & _T_60094; // @[Switch.scala 41:38:@21254.4]
  assign _T_60097 = select_41 == 6'h2; // @[Switch.scala 41:52:@21256.4]
  assign output_2_41 = io_outValid_41 & _T_60097; // @[Switch.scala 41:38:@21257.4]
  assign _T_60100 = select_42 == 6'h2; // @[Switch.scala 41:52:@21259.4]
  assign output_2_42 = io_outValid_42 & _T_60100; // @[Switch.scala 41:38:@21260.4]
  assign _T_60103 = select_43 == 6'h2; // @[Switch.scala 41:52:@21262.4]
  assign output_2_43 = io_outValid_43 & _T_60103; // @[Switch.scala 41:38:@21263.4]
  assign _T_60106 = select_44 == 6'h2; // @[Switch.scala 41:52:@21265.4]
  assign output_2_44 = io_outValid_44 & _T_60106; // @[Switch.scala 41:38:@21266.4]
  assign _T_60109 = select_45 == 6'h2; // @[Switch.scala 41:52:@21268.4]
  assign output_2_45 = io_outValid_45 & _T_60109; // @[Switch.scala 41:38:@21269.4]
  assign _T_60112 = select_46 == 6'h2; // @[Switch.scala 41:52:@21271.4]
  assign output_2_46 = io_outValid_46 & _T_60112; // @[Switch.scala 41:38:@21272.4]
  assign _T_60115 = select_47 == 6'h2; // @[Switch.scala 41:52:@21274.4]
  assign output_2_47 = io_outValid_47 & _T_60115; // @[Switch.scala 41:38:@21275.4]
  assign _T_60118 = select_48 == 6'h2; // @[Switch.scala 41:52:@21277.4]
  assign output_2_48 = io_outValid_48 & _T_60118; // @[Switch.scala 41:38:@21278.4]
  assign _T_60121 = select_49 == 6'h2; // @[Switch.scala 41:52:@21280.4]
  assign output_2_49 = io_outValid_49 & _T_60121; // @[Switch.scala 41:38:@21281.4]
  assign _T_60124 = select_50 == 6'h2; // @[Switch.scala 41:52:@21283.4]
  assign output_2_50 = io_outValid_50 & _T_60124; // @[Switch.scala 41:38:@21284.4]
  assign _T_60127 = select_51 == 6'h2; // @[Switch.scala 41:52:@21286.4]
  assign output_2_51 = io_outValid_51 & _T_60127; // @[Switch.scala 41:38:@21287.4]
  assign _T_60130 = select_52 == 6'h2; // @[Switch.scala 41:52:@21289.4]
  assign output_2_52 = io_outValid_52 & _T_60130; // @[Switch.scala 41:38:@21290.4]
  assign _T_60133 = select_53 == 6'h2; // @[Switch.scala 41:52:@21292.4]
  assign output_2_53 = io_outValid_53 & _T_60133; // @[Switch.scala 41:38:@21293.4]
  assign _T_60136 = select_54 == 6'h2; // @[Switch.scala 41:52:@21295.4]
  assign output_2_54 = io_outValid_54 & _T_60136; // @[Switch.scala 41:38:@21296.4]
  assign _T_60139 = select_55 == 6'h2; // @[Switch.scala 41:52:@21298.4]
  assign output_2_55 = io_outValid_55 & _T_60139; // @[Switch.scala 41:38:@21299.4]
  assign _T_60142 = select_56 == 6'h2; // @[Switch.scala 41:52:@21301.4]
  assign output_2_56 = io_outValid_56 & _T_60142; // @[Switch.scala 41:38:@21302.4]
  assign _T_60145 = select_57 == 6'h2; // @[Switch.scala 41:52:@21304.4]
  assign output_2_57 = io_outValid_57 & _T_60145; // @[Switch.scala 41:38:@21305.4]
  assign _T_60148 = select_58 == 6'h2; // @[Switch.scala 41:52:@21307.4]
  assign output_2_58 = io_outValid_58 & _T_60148; // @[Switch.scala 41:38:@21308.4]
  assign _T_60151 = select_59 == 6'h2; // @[Switch.scala 41:52:@21310.4]
  assign output_2_59 = io_outValid_59 & _T_60151; // @[Switch.scala 41:38:@21311.4]
  assign _T_60154 = select_60 == 6'h2; // @[Switch.scala 41:52:@21313.4]
  assign output_2_60 = io_outValid_60 & _T_60154; // @[Switch.scala 41:38:@21314.4]
  assign _T_60157 = select_61 == 6'h2; // @[Switch.scala 41:52:@21316.4]
  assign output_2_61 = io_outValid_61 & _T_60157; // @[Switch.scala 41:38:@21317.4]
  assign _T_60160 = select_62 == 6'h2; // @[Switch.scala 41:52:@21319.4]
  assign output_2_62 = io_outValid_62 & _T_60160; // @[Switch.scala 41:38:@21320.4]
  assign _T_60163 = select_63 == 6'h2; // @[Switch.scala 41:52:@21322.4]
  assign output_2_63 = io_outValid_63 & _T_60163; // @[Switch.scala 41:38:@21323.4]
  assign _T_60171 = {output_2_7,output_2_6,output_2_5,output_2_4,output_2_3,output_2_2,output_2_1,output_2_0}; // @[Switch.scala 43:31:@21331.4]
  assign _T_60179 = {output_2_15,output_2_14,output_2_13,output_2_12,output_2_11,output_2_10,output_2_9,output_2_8,_T_60171}; // @[Switch.scala 43:31:@21339.4]
  assign _T_60186 = {output_2_23,output_2_22,output_2_21,output_2_20,output_2_19,output_2_18,output_2_17,output_2_16}; // @[Switch.scala 43:31:@21346.4]
  assign _T_60195 = {output_2_31,output_2_30,output_2_29,output_2_28,output_2_27,output_2_26,output_2_25,output_2_24,_T_60186,_T_60179}; // @[Switch.scala 43:31:@21355.4]
  assign _T_60202 = {output_2_39,output_2_38,output_2_37,output_2_36,output_2_35,output_2_34,output_2_33,output_2_32}; // @[Switch.scala 43:31:@21362.4]
  assign _T_60210 = {output_2_47,output_2_46,output_2_45,output_2_44,output_2_43,output_2_42,output_2_41,output_2_40,_T_60202}; // @[Switch.scala 43:31:@21370.4]
  assign _T_60217 = {output_2_55,output_2_54,output_2_53,output_2_52,output_2_51,output_2_50,output_2_49,output_2_48}; // @[Switch.scala 43:31:@21377.4]
  assign _T_60226 = {output_2_63,output_2_62,output_2_61,output_2_60,output_2_59,output_2_58,output_2_57,output_2_56,_T_60217,_T_60210}; // @[Switch.scala 43:31:@21386.4]
  assign _T_60227 = {_T_60226,_T_60195}; // @[Switch.scala 43:31:@21387.4]
  assign _T_60231 = select_0 == 6'h3; // @[Switch.scala 41:52:@21390.4]
  assign output_3_0 = io_outValid_0 & _T_60231; // @[Switch.scala 41:38:@21391.4]
  assign _T_60234 = select_1 == 6'h3; // @[Switch.scala 41:52:@21393.4]
  assign output_3_1 = io_outValid_1 & _T_60234; // @[Switch.scala 41:38:@21394.4]
  assign _T_60237 = select_2 == 6'h3; // @[Switch.scala 41:52:@21396.4]
  assign output_3_2 = io_outValid_2 & _T_60237; // @[Switch.scala 41:38:@21397.4]
  assign _T_60240 = select_3 == 6'h3; // @[Switch.scala 41:52:@21399.4]
  assign output_3_3 = io_outValid_3 & _T_60240; // @[Switch.scala 41:38:@21400.4]
  assign _T_60243 = select_4 == 6'h3; // @[Switch.scala 41:52:@21402.4]
  assign output_3_4 = io_outValid_4 & _T_60243; // @[Switch.scala 41:38:@21403.4]
  assign _T_60246 = select_5 == 6'h3; // @[Switch.scala 41:52:@21405.4]
  assign output_3_5 = io_outValid_5 & _T_60246; // @[Switch.scala 41:38:@21406.4]
  assign _T_60249 = select_6 == 6'h3; // @[Switch.scala 41:52:@21408.4]
  assign output_3_6 = io_outValid_6 & _T_60249; // @[Switch.scala 41:38:@21409.4]
  assign _T_60252 = select_7 == 6'h3; // @[Switch.scala 41:52:@21411.4]
  assign output_3_7 = io_outValid_7 & _T_60252; // @[Switch.scala 41:38:@21412.4]
  assign _T_60255 = select_8 == 6'h3; // @[Switch.scala 41:52:@21414.4]
  assign output_3_8 = io_outValid_8 & _T_60255; // @[Switch.scala 41:38:@21415.4]
  assign _T_60258 = select_9 == 6'h3; // @[Switch.scala 41:52:@21417.4]
  assign output_3_9 = io_outValid_9 & _T_60258; // @[Switch.scala 41:38:@21418.4]
  assign _T_60261 = select_10 == 6'h3; // @[Switch.scala 41:52:@21420.4]
  assign output_3_10 = io_outValid_10 & _T_60261; // @[Switch.scala 41:38:@21421.4]
  assign _T_60264 = select_11 == 6'h3; // @[Switch.scala 41:52:@21423.4]
  assign output_3_11 = io_outValid_11 & _T_60264; // @[Switch.scala 41:38:@21424.4]
  assign _T_60267 = select_12 == 6'h3; // @[Switch.scala 41:52:@21426.4]
  assign output_3_12 = io_outValid_12 & _T_60267; // @[Switch.scala 41:38:@21427.4]
  assign _T_60270 = select_13 == 6'h3; // @[Switch.scala 41:52:@21429.4]
  assign output_3_13 = io_outValid_13 & _T_60270; // @[Switch.scala 41:38:@21430.4]
  assign _T_60273 = select_14 == 6'h3; // @[Switch.scala 41:52:@21432.4]
  assign output_3_14 = io_outValid_14 & _T_60273; // @[Switch.scala 41:38:@21433.4]
  assign _T_60276 = select_15 == 6'h3; // @[Switch.scala 41:52:@21435.4]
  assign output_3_15 = io_outValid_15 & _T_60276; // @[Switch.scala 41:38:@21436.4]
  assign _T_60279 = select_16 == 6'h3; // @[Switch.scala 41:52:@21438.4]
  assign output_3_16 = io_outValid_16 & _T_60279; // @[Switch.scala 41:38:@21439.4]
  assign _T_60282 = select_17 == 6'h3; // @[Switch.scala 41:52:@21441.4]
  assign output_3_17 = io_outValid_17 & _T_60282; // @[Switch.scala 41:38:@21442.4]
  assign _T_60285 = select_18 == 6'h3; // @[Switch.scala 41:52:@21444.4]
  assign output_3_18 = io_outValid_18 & _T_60285; // @[Switch.scala 41:38:@21445.4]
  assign _T_60288 = select_19 == 6'h3; // @[Switch.scala 41:52:@21447.4]
  assign output_3_19 = io_outValid_19 & _T_60288; // @[Switch.scala 41:38:@21448.4]
  assign _T_60291 = select_20 == 6'h3; // @[Switch.scala 41:52:@21450.4]
  assign output_3_20 = io_outValid_20 & _T_60291; // @[Switch.scala 41:38:@21451.4]
  assign _T_60294 = select_21 == 6'h3; // @[Switch.scala 41:52:@21453.4]
  assign output_3_21 = io_outValid_21 & _T_60294; // @[Switch.scala 41:38:@21454.4]
  assign _T_60297 = select_22 == 6'h3; // @[Switch.scala 41:52:@21456.4]
  assign output_3_22 = io_outValid_22 & _T_60297; // @[Switch.scala 41:38:@21457.4]
  assign _T_60300 = select_23 == 6'h3; // @[Switch.scala 41:52:@21459.4]
  assign output_3_23 = io_outValid_23 & _T_60300; // @[Switch.scala 41:38:@21460.4]
  assign _T_60303 = select_24 == 6'h3; // @[Switch.scala 41:52:@21462.4]
  assign output_3_24 = io_outValid_24 & _T_60303; // @[Switch.scala 41:38:@21463.4]
  assign _T_60306 = select_25 == 6'h3; // @[Switch.scala 41:52:@21465.4]
  assign output_3_25 = io_outValid_25 & _T_60306; // @[Switch.scala 41:38:@21466.4]
  assign _T_60309 = select_26 == 6'h3; // @[Switch.scala 41:52:@21468.4]
  assign output_3_26 = io_outValid_26 & _T_60309; // @[Switch.scala 41:38:@21469.4]
  assign _T_60312 = select_27 == 6'h3; // @[Switch.scala 41:52:@21471.4]
  assign output_3_27 = io_outValid_27 & _T_60312; // @[Switch.scala 41:38:@21472.4]
  assign _T_60315 = select_28 == 6'h3; // @[Switch.scala 41:52:@21474.4]
  assign output_3_28 = io_outValid_28 & _T_60315; // @[Switch.scala 41:38:@21475.4]
  assign _T_60318 = select_29 == 6'h3; // @[Switch.scala 41:52:@21477.4]
  assign output_3_29 = io_outValid_29 & _T_60318; // @[Switch.scala 41:38:@21478.4]
  assign _T_60321 = select_30 == 6'h3; // @[Switch.scala 41:52:@21480.4]
  assign output_3_30 = io_outValid_30 & _T_60321; // @[Switch.scala 41:38:@21481.4]
  assign _T_60324 = select_31 == 6'h3; // @[Switch.scala 41:52:@21483.4]
  assign output_3_31 = io_outValid_31 & _T_60324; // @[Switch.scala 41:38:@21484.4]
  assign _T_60327 = select_32 == 6'h3; // @[Switch.scala 41:52:@21486.4]
  assign output_3_32 = io_outValid_32 & _T_60327; // @[Switch.scala 41:38:@21487.4]
  assign _T_60330 = select_33 == 6'h3; // @[Switch.scala 41:52:@21489.4]
  assign output_3_33 = io_outValid_33 & _T_60330; // @[Switch.scala 41:38:@21490.4]
  assign _T_60333 = select_34 == 6'h3; // @[Switch.scala 41:52:@21492.4]
  assign output_3_34 = io_outValid_34 & _T_60333; // @[Switch.scala 41:38:@21493.4]
  assign _T_60336 = select_35 == 6'h3; // @[Switch.scala 41:52:@21495.4]
  assign output_3_35 = io_outValid_35 & _T_60336; // @[Switch.scala 41:38:@21496.4]
  assign _T_60339 = select_36 == 6'h3; // @[Switch.scala 41:52:@21498.4]
  assign output_3_36 = io_outValid_36 & _T_60339; // @[Switch.scala 41:38:@21499.4]
  assign _T_60342 = select_37 == 6'h3; // @[Switch.scala 41:52:@21501.4]
  assign output_3_37 = io_outValid_37 & _T_60342; // @[Switch.scala 41:38:@21502.4]
  assign _T_60345 = select_38 == 6'h3; // @[Switch.scala 41:52:@21504.4]
  assign output_3_38 = io_outValid_38 & _T_60345; // @[Switch.scala 41:38:@21505.4]
  assign _T_60348 = select_39 == 6'h3; // @[Switch.scala 41:52:@21507.4]
  assign output_3_39 = io_outValid_39 & _T_60348; // @[Switch.scala 41:38:@21508.4]
  assign _T_60351 = select_40 == 6'h3; // @[Switch.scala 41:52:@21510.4]
  assign output_3_40 = io_outValid_40 & _T_60351; // @[Switch.scala 41:38:@21511.4]
  assign _T_60354 = select_41 == 6'h3; // @[Switch.scala 41:52:@21513.4]
  assign output_3_41 = io_outValid_41 & _T_60354; // @[Switch.scala 41:38:@21514.4]
  assign _T_60357 = select_42 == 6'h3; // @[Switch.scala 41:52:@21516.4]
  assign output_3_42 = io_outValid_42 & _T_60357; // @[Switch.scala 41:38:@21517.4]
  assign _T_60360 = select_43 == 6'h3; // @[Switch.scala 41:52:@21519.4]
  assign output_3_43 = io_outValid_43 & _T_60360; // @[Switch.scala 41:38:@21520.4]
  assign _T_60363 = select_44 == 6'h3; // @[Switch.scala 41:52:@21522.4]
  assign output_3_44 = io_outValid_44 & _T_60363; // @[Switch.scala 41:38:@21523.4]
  assign _T_60366 = select_45 == 6'h3; // @[Switch.scala 41:52:@21525.4]
  assign output_3_45 = io_outValid_45 & _T_60366; // @[Switch.scala 41:38:@21526.4]
  assign _T_60369 = select_46 == 6'h3; // @[Switch.scala 41:52:@21528.4]
  assign output_3_46 = io_outValid_46 & _T_60369; // @[Switch.scala 41:38:@21529.4]
  assign _T_60372 = select_47 == 6'h3; // @[Switch.scala 41:52:@21531.4]
  assign output_3_47 = io_outValid_47 & _T_60372; // @[Switch.scala 41:38:@21532.4]
  assign _T_60375 = select_48 == 6'h3; // @[Switch.scala 41:52:@21534.4]
  assign output_3_48 = io_outValid_48 & _T_60375; // @[Switch.scala 41:38:@21535.4]
  assign _T_60378 = select_49 == 6'h3; // @[Switch.scala 41:52:@21537.4]
  assign output_3_49 = io_outValid_49 & _T_60378; // @[Switch.scala 41:38:@21538.4]
  assign _T_60381 = select_50 == 6'h3; // @[Switch.scala 41:52:@21540.4]
  assign output_3_50 = io_outValid_50 & _T_60381; // @[Switch.scala 41:38:@21541.4]
  assign _T_60384 = select_51 == 6'h3; // @[Switch.scala 41:52:@21543.4]
  assign output_3_51 = io_outValid_51 & _T_60384; // @[Switch.scala 41:38:@21544.4]
  assign _T_60387 = select_52 == 6'h3; // @[Switch.scala 41:52:@21546.4]
  assign output_3_52 = io_outValid_52 & _T_60387; // @[Switch.scala 41:38:@21547.4]
  assign _T_60390 = select_53 == 6'h3; // @[Switch.scala 41:52:@21549.4]
  assign output_3_53 = io_outValid_53 & _T_60390; // @[Switch.scala 41:38:@21550.4]
  assign _T_60393 = select_54 == 6'h3; // @[Switch.scala 41:52:@21552.4]
  assign output_3_54 = io_outValid_54 & _T_60393; // @[Switch.scala 41:38:@21553.4]
  assign _T_60396 = select_55 == 6'h3; // @[Switch.scala 41:52:@21555.4]
  assign output_3_55 = io_outValid_55 & _T_60396; // @[Switch.scala 41:38:@21556.4]
  assign _T_60399 = select_56 == 6'h3; // @[Switch.scala 41:52:@21558.4]
  assign output_3_56 = io_outValid_56 & _T_60399; // @[Switch.scala 41:38:@21559.4]
  assign _T_60402 = select_57 == 6'h3; // @[Switch.scala 41:52:@21561.4]
  assign output_3_57 = io_outValid_57 & _T_60402; // @[Switch.scala 41:38:@21562.4]
  assign _T_60405 = select_58 == 6'h3; // @[Switch.scala 41:52:@21564.4]
  assign output_3_58 = io_outValid_58 & _T_60405; // @[Switch.scala 41:38:@21565.4]
  assign _T_60408 = select_59 == 6'h3; // @[Switch.scala 41:52:@21567.4]
  assign output_3_59 = io_outValid_59 & _T_60408; // @[Switch.scala 41:38:@21568.4]
  assign _T_60411 = select_60 == 6'h3; // @[Switch.scala 41:52:@21570.4]
  assign output_3_60 = io_outValid_60 & _T_60411; // @[Switch.scala 41:38:@21571.4]
  assign _T_60414 = select_61 == 6'h3; // @[Switch.scala 41:52:@21573.4]
  assign output_3_61 = io_outValid_61 & _T_60414; // @[Switch.scala 41:38:@21574.4]
  assign _T_60417 = select_62 == 6'h3; // @[Switch.scala 41:52:@21576.4]
  assign output_3_62 = io_outValid_62 & _T_60417; // @[Switch.scala 41:38:@21577.4]
  assign _T_60420 = select_63 == 6'h3; // @[Switch.scala 41:52:@21579.4]
  assign output_3_63 = io_outValid_63 & _T_60420; // @[Switch.scala 41:38:@21580.4]
  assign _T_60428 = {output_3_7,output_3_6,output_3_5,output_3_4,output_3_3,output_3_2,output_3_1,output_3_0}; // @[Switch.scala 43:31:@21588.4]
  assign _T_60436 = {output_3_15,output_3_14,output_3_13,output_3_12,output_3_11,output_3_10,output_3_9,output_3_8,_T_60428}; // @[Switch.scala 43:31:@21596.4]
  assign _T_60443 = {output_3_23,output_3_22,output_3_21,output_3_20,output_3_19,output_3_18,output_3_17,output_3_16}; // @[Switch.scala 43:31:@21603.4]
  assign _T_60452 = {output_3_31,output_3_30,output_3_29,output_3_28,output_3_27,output_3_26,output_3_25,output_3_24,_T_60443,_T_60436}; // @[Switch.scala 43:31:@21612.4]
  assign _T_60459 = {output_3_39,output_3_38,output_3_37,output_3_36,output_3_35,output_3_34,output_3_33,output_3_32}; // @[Switch.scala 43:31:@21619.4]
  assign _T_60467 = {output_3_47,output_3_46,output_3_45,output_3_44,output_3_43,output_3_42,output_3_41,output_3_40,_T_60459}; // @[Switch.scala 43:31:@21627.4]
  assign _T_60474 = {output_3_55,output_3_54,output_3_53,output_3_52,output_3_51,output_3_50,output_3_49,output_3_48}; // @[Switch.scala 43:31:@21634.4]
  assign _T_60483 = {output_3_63,output_3_62,output_3_61,output_3_60,output_3_59,output_3_58,output_3_57,output_3_56,_T_60474,_T_60467}; // @[Switch.scala 43:31:@21643.4]
  assign _T_60484 = {_T_60483,_T_60452}; // @[Switch.scala 43:31:@21644.4]
  assign _T_60488 = select_0 == 6'h4; // @[Switch.scala 41:52:@21647.4]
  assign output_4_0 = io_outValid_0 & _T_60488; // @[Switch.scala 41:38:@21648.4]
  assign _T_60491 = select_1 == 6'h4; // @[Switch.scala 41:52:@21650.4]
  assign output_4_1 = io_outValid_1 & _T_60491; // @[Switch.scala 41:38:@21651.4]
  assign _T_60494 = select_2 == 6'h4; // @[Switch.scala 41:52:@21653.4]
  assign output_4_2 = io_outValid_2 & _T_60494; // @[Switch.scala 41:38:@21654.4]
  assign _T_60497 = select_3 == 6'h4; // @[Switch.scala 41:52:@21656.4]
  assign output_4_3 = io_outValid_3 & _T_60497; // @[Switch.scala 41:38:@21657.4]
  assign _T_60500 = select_4 == 6'h4; // @[Switch.scala 41:52:@21659.4]
  assign output_4_4 = io_outValid_4 & _T_60500; // @[Switch.scala 41:38:@21660.4]
  assign _T_60503 = select_5 == 6'h4; // @[Switch.scala 41:52:@21662.4]
  assign output_4_5 = io_outValid_5 & _T_60503; // @[Switch.scala 41:38:@21663.4]
  assign _T_60506 = select_6 == 6'h4; // @[Switch.scala 41:52:@21665.4]
  assign output_4_6 = io_outValid_6 & _T_60506; // @[Switch.scala 41:38:@21666.4]
  assign _T_60509 = select_7 == 6'h4; // @[Switch.scala 41:52:@21668.4]
  assign output_4_7 = io_outValid_7 & _T_60509; // @[Switch.scala 41:38:@21669.4]
  assign _T_60512 = select_8 == 6'h4; // @[Switch.scala 41:52:@21671.4]
  assign output_4_8 = io_outValid_8 & _T_60512; // @[Switch.scala 41:38:@21672.4]
  assign _T_60515 = select_9 == 6'h4; // @[Switch.scala 41:52:@21674.4]
  assign output_4_9 = io_outValid_9 & _T_60515; // @[Switch.scala 41:38:@21675.4]
  assign _T_60518 = select_10 == 6'h4; // @[Switch.scala 41:52:@21677.4]
  assign output_4_10 = io_outValid_10 & _T_60518; // @[Switch.scala 41:38:@21678.4]
  assign _T_60521 = select_11 == 6'h4; // @[Switch.scala 41:52:@21680.4]
  assign output_4_11 = io_outValid_11 & _T_60521; // @[Switch.scala 41:38:@21681.4]
  assign _T_60524 = select_12 == 6'h4; // @[Switch.scala 41:52:@21683.4]
  assign output_4_12 = io_outValid_12 & _T_60524; // @[Switch.scala 41:38:@21684.4]
  assign _T_60527 = select_13 == 6'h4; // @[Switch.scala 41:52:@21686.4]
  assign output_4_13 = io_outValid_13 & _T_60527; // @[Switch.scala 41:38:@21687.4]
  assign _T_60530 = select_14 == 6'h4; // @[Switch.scala 41:52:@21689.4]
  assign output_4_14 = io_outValid_14 & _T_60530; // @[Switch.scala 41:38:@21690.4]
  assign _T_60533 = select_15 == 6'h4; // @[Switch.scala 41:52:@21692.4]
  assign output_4_15 = io_outValid_15 & _T_60533; // @[Switch.scala 41:38:@21693.4]
  assign _T_60536 = select_16 == 6'h4; // @[Switch.scala 41:52:@21695.4]
  assign output_4_16 = io_outValid_16 & _T_60536; // @[Switch.scala 41:38:@21696.4]
  assign _T_60539 = select_17 == 6'h4; // @[Switch.scala 41:52:@21698.4]
  assign output_4_17 = io_outValid_17 & _T_60539; // @[Switch.scala 41:38:@21699.4]
  assign _T_60542 = select_18 == 6'h4; // @[Switch.scala 41:52:@21701.4]
  assign output_4_18 = io_outValid_18 & _T_60542; // @[Switch.scala 41:38:@21702.4]
  assign _T_60545 = select_19 == 6'h4; // @[Switch.scala 41:52:@21704.4]
  assign output_4_19 = io_outValid_19 & _T_60545; // @[Switch.scala 41:38:@21705.4]
  assign _T_60548 = select_20 == 6'h4; // @[Switch.scala 41:52:@21707.4]
  assign output_4_20 = io_outValid_20 & _T_60548; // @[Switch.scala 41:38:@21708.4]
  assign _T_60551 = select_21 == 6'h4; // @[Switch.scala 41:52:@21710.4]
  assign output_4_21 = io_outValid_21 & _T_60551; // @[Switch.scala 41:38:@21711.4]
  assign _T_60554 = select_22 == 6'h4; // @[Switch.scala 41:52:@21713.4]
  assign output_4_22 = io_outValid_22 & _T_60554; // @[Switch.scala 41:38:@21714.4]
  assign _T_60557 = select_23 == 6'h4; // @[Switch.scala 41:52:@21716.4]
  assign output_4_23 = io_outValid_23 & _T_60557; // @[Switch.scala 41:38:@21717.4]
  assign _T_60560 = select_24 == 6'h4; // @[Switch.scala 41:52:@21719.4]
  assign output_4_24 = io_outValid_24 & _T_60560; // @[Switch.scala 41:38:@21720.4]
  assign _T_60563 = select_25 == 6'h4; // @[Switch.scala 41:52:@21722.4]
  assign output_4_25 = io_outValid_25 & _T_60563; // @[Switch.scala 41:38:@21723.4]
  assign _T_60566 = select_26 == 6'h4; // @[Switch.scala 41:52:@21725.4]
  assign output_4_26 = io_outValid_26 & _T_60566; // @[Switch.scala 41:38:@21726.4]
  assign _T_60569 = select_27 == 6'h4; // @[Switch.scala 41:52:@21728.4]
  assign output_4_27 = io_outValid_27 & _T_60569; // @[Switch.scala 41:38:@21729.4]
  assign _T_60572 = select_28 == 6'h4; // @[Switch.scala 41:52:@21731.4]
  assign output_4_28 = io_outValid_28 & _T_60572; // @[Switch.scala 41:38:@21732.4]
  assign _T_60575 = select_29 == 6'h4; // @[Switch.scala 41:52:@21734.4]
  assign output_4_29 = io_outValid_29 & _T_60575; // @[Switch.scala 41:38:@21735.4]
  assign _T_60578 = select_30 == 6'h4; // @[Switch.scala 41:52:@21737.4]
  assign output_4_30 = io_outValid_30 & _T_60578; // @[Switch.scala 41:38:@21738.4]
  assign _T_60581 = select_31 == 6'h4; // @[Switch.scala 41:52:@21740.4]
  assign output_4_31 = io_outValid_31 & _T_60581; // @[Switch.scala 41:38:@21741.4]
  assign _T_60584 = select_32 == 6'h4; // @[Switch.scala 41:52:@21743.4]
  assign output_4_32 = io_outValid_32 & _T_60584; // @[Switch.scala 41:38:@21744.4]
  assign _T_60587 = select_33 == 6'h4; // @[Switch.scala 41:52:@21746.4]
  assign output_4_33 = io_outValid_33 & _T_60587; // @[Switch.scala 41:38:@21747.4]
  assign _T_60590 = select_34 == 6'h4; // @[Switch.scala 41:52:@21749.4]
  assign output_4_34 = io_outValid_34 & _T_60590; // @[Switch.scala 41:38:@21750.4]
  assign _T_60593 = select_35 == 6'h4; // @[Switch.scala 41:52:@21752.4]
  assign output_4_35 = io_outValid_35 & _T_60593; // @[Switch.scala 41:38:@21753.4]
  assign _T_60596 = select_36 == 6'h4; // @[Switch.scala 41:52:@21755.4]
  assign output_4_36 = io_outValid_36 & _T_60596; // @[Switch.scala 41:38:@21756.4]
  assign _T_60599 = select_37 == 6'h4; // @[Switch.scala 41:52:@21758.4]
  assign output_4_37 = io_outValid_37 & _T_60599; // @[Switch.scala 41:38:@21759.4]
  assign _T_60602 = select_38 == 6'h4; // @[Switch.scala 41:52:@21761.4]
  assign output_4_38 = io_outValid_38 & _T_60602; // @[Switch.scala 41:38:@21762.4]
  assign _T_60605 = select_39 == 6'h4; // @[Switch.scala 41:52:@21764.4]
  assign output_4_39 = io_outValid_39 & _T_60605; // @[Switch.scala 41:38:@21765.4]
  assign _T_60608 = select_40 == 6'h4; // @[Switch.scala 41:52:@21767.4]
  assign output_4_40 = io_outValid_40 & _T_60608; // @[Switch.scala 41:38:@21768.4]
  assign _T_60611 = select_41 == 6'h4; // @[Switch.scala 41:52:@21770.4]
  assign output_4_41 = io_outValid_41 & _T_60611; // @[Switch.scala 41:38:@21771.4]
  assign _T_60614 = select_42 == 6'h4; // @[Switch.scala 41:52:@21773.4]
  assign output_4_42 = io_outValid_42 & _T_60614; // @[Switch.scala 41:38:@21774.4]
  assign _T_60617 = select_43 == 6'h4; // @[Switch.scala 41:52:@21776.4]
  assign output_4_43 = io_outValid_43 & _T_60617; // @[Switch.scala 41:38:@21777.4]
  assign _T_60620 = select_44 == 6'h4; // @[Switch.scala 41:52:@21779.4]
  assign output_4_44 = io_outValid_44 & _T_60620; // @[Switch.scala 41:38:@21780.4]
  assign _T_60623 = select_45 == 6'h4; // @[Switch.scala 41:52:@21782.4]
  assign output_4_45 = io_outValid_45 & _T_60623; // @[Switch.scala 41:38:@21783.4]
  assign _T_60626 = select_46 == 6'h4; // @[Switch.scala 41:52:@21785.4]
  assign output_4_46 = io_outValid_46 & _T_60626; // @[Switch.scala 41:38:@21786.4]
  assign _T_60629 = select_47 == 6'h4; // @[Switch.scala 41:52:@21788.4]
  assign output_4_47 = io_outValid_47 & _T_60629; // @[Switch.scala 41:38:@21789.4]
  assign _T_60632 = select_48 == 6'h4; // @[Switch.scala 41:52:@21791.4]
  assign output_4_48 = io_outValid_48 & _T_60632; // @[Switch.scala 41:38:@21792.4]
  assign _T_60635 = select_49 == 6'h4; // @[Switch.scala 41:52:@21794.4]
  assign output_4_49 = io_outValid_49 & _T_60635; // @[Switch.scala 41:38:@21795.4]
  assign _T_60638 = select_50 == 6'h4; // @[Switch.scala 41:52:@21797.4]
  assign output_4_50 = io_outValid_50 & _T_60638; // @[Switch.scala 41:38:@21798.4]
  assign _T_60641 = select_51 == 6'h4; // @[Switch.scala 41:52:@21800.4]
  assign output_4_51 = io_outValid_51 & _T_60641; // @[Switch.scala 41:38:@21801.4]
  assign _T_60644 = select_52 == 6'h4; // @[Switch.scala 41:52:@21803.4]
  assign output_4_52 = io_outValid_52 & _T_60644; // @[Switch.scala 41:38:@21804.4]
  assign _T_60647 = select_53 == 6'h4; // @[Switch.scala 41:52:@21806.4]
  assign output_4_53 = io_outValid_53 & _T_60647; // @[Switch.scala 41:38:@21807.4]
  assign _T_60650 = select_54 == 6'h4; // @[Switch.scala 41:52:@21809.4]
  assign output_4_54 = io_outValid_54 & _T_60650; // @[Switch.scala 41:38:@21810.4]
  assign _T_60653 = select_55 == 6'h4; // @[Switch.scala 41:52:@21812.4]
  assign output_4_55 = io_outValid_55 & _T_60653; // @[Switch.scala 41:38:@21813.4]
  assign _T_60656 = select_56 == 6'h4; // @[Switch.scala 41:52:@21815.4]
  assign output_4_56 = io_outValid_56 & _T_60656; // @[Switch.scala 41:38:@21816.4]
  assign _T_60659 = select_57 == 6'h4; // @[Switch.scala 41:52:@21818.4]
  assign output_4_57 = io_outValid_57 & _T_60659; // @[Switch.scala 41:38:@21819.4]
  assign _T_60662 = select_58 == 6'h4; // @[Switch.scala 41:52:@21821.4]
  assign output_4_58 = io_outValid_58 & _T_60662; // @[Switch.scala 41:38:@21822.4]
  assign _T_60665 = select_59 == 6'h4; // @[Switch.scala 41:52:@21824.4]
  assign output_4_59 = io_outValid_59 & _T_60665; // @[Switch.scala 41:38:@21825.4]
  assign _T_60668 = select_60 == 6'h4; // @[Switch.scala 41:52:@21827.4]
  assign output_4_60 = io_outValid_60 & _T_60668; // @[Switch.scala 41:38:@21828.4]
  assign _T_60671 = select_61 == 6'h4; // @[Switch.scala 41:52:@21830.4]
  assign output_4_61 = io_outValid_61 & _T_60671; // @[Switch.scala 41:38:@21831.4]
  assign _T_60674 = select_62 == 6'h4; // @[Switch.scala 41:52:@21833.4]
  assign output_4_62 = io_outValid_62 & _T_60674; // @[Switch.scala 41:38:@21834.4]
  assign _T_60677 = select_63 == 6'h4; // @[Switch.scala 41:52:@21836.4]
  assign output_4_63 = io_outValid_63 & _T_60677; // @[Switch.scala 41:38:@21837.4]
  assign _T_60685 = {output_4_7,output_4_6,output_4_5,output_4_4,output_4_3,output_4_2,output_4_1,output_4_0}; // @[Switch.scala 43:31:@21845.4]
  assign _T_60693 = {output_4_15,output_4_14,output_4_13,output_4_12,output_4_11,output_4_10,output_4_9,output_4_8,_T_60685}; // @[Switch.scala 43:31:@21853.4]
  assign _T_60700 = {output_4_23,output_4_22,output_4_21,output_4_20,output_4_19,output_4_18,output_4_17,output_4_16}; // @[Switch.scala 43:31:@21860.4]
  assign _T_60709 = {output_4_31,output_4_30,output_4_29,output_4_28,output_4_27,output_4_26,output_4_25,output_4_24,_T_60700,_T_60693}; // @[Switch.scala 43:31:@21869.4]
  assign _T_60716 = {output_4_39,output_4_38,output_4_37,output_4_36,output_4_35,output_4_34,output_4_33,output_4_32}; // @[Switch.scala 43:31:@21876.4]
  assign _T_60724 = {output_4_47,output_4_46,output_4_45,output_4_44,output_4_43,output_4_42,output_4_41,output_4_40,_T_60716}; // @[Switch.scala 43:31:@21884.4]
  assign _T_60731 = {output_4_55,output_4_54,output_4_53,output_4_52,output_4_51,output_4_50,output_4_49,output_4_48}; // @[Switch.scala 43:31:@21891.4]
  assign _T_60740 = {output_4_63,output_4_62,output_4_61,output_4_60,output_4_59,output_4_58,output_4_57,output_4_56,_T_60731,_T_60724}; // @[Switch.scala 43:31:@21900.4]
  assign _T_60741 = {_T_60740,_T_60709}; // @[Switch.scala 43:31:@21901.4]
  assign _T_60745 = select_0 == 6'h5; // @[Switch.scala 41:52:@21904.4]
  assign output_5_0 = io_outValid_0 & _T_60745; // @[Switch.scala 41:38:@21905.4]
  assign _T_60748 = select_1 == 6'h5; // @[Switch.scala 41:52:@21907.4]
  assign output_5_1 = io_outValid_1 & _T_60748; // @[Switch.scala 41:38:@21908.4]
  assign _T_60751 = select_2 == 6'h5; // @[Switch.scala 41:52:@21910.4]
  assign output_5_2 = io_outValid_2 & _T_60751; // @[Switch.scala 41:38:@21911.4]
  assign _T_60754 = select_3 == 6'h5; // @[Switch.scala 41:52:@21913.4]
  assign output_5_3 = io_outValid_3 & _T_60754; // @[Switch.scala 41:38:@21914.4]
  assign _T_60757 = select_4 == 6'h5; // @[Switch.scala 41:52:@21916.4]
  assign output_5_4 = io_outValid_4 & _T_60757; // @[Switch.scala 41:38:@21917.4]
  assign _T_60760 = select_5 == 6'h5; // @[Switch.scala 41:52:@21919.4]
  assign output_5_5 = io_outValid_5 & _T_60760; // @[Switch.scala 41:38:@21920.4]
  assign _T_60763 = select_6 == 6'h5; // @[Switch.scala 41:52:@21922.4]
  assign output_5_6 = io_outValid_6 & _T_60763; // @[Switch.scala 41:38:@21923.4]
  assign _T_60766 = select_7 == 6'h5; // @[Switch.scala 41:52:@21925.4]
  assign output_5_7 = io_outValid_7 & _T_60766; // @[Switch.scala 41:38:@21926.4]
  assign _T_60769 = select_8 == 6'h5; // @[Switch.scala 41:52:@21928.4]
  assign output_5_8 = io_outValid_8 & _T_60769; // @[Switch.scala 41:38:@21929.4]
  assign _T_60772 = select_9 == 6'h5; // @[Switch.scala 41:52:@21931.4]
  assign output_5_9 = io_outValid_9 & _T_60772; // @[Switch.scala 41:38:@21932.4]
  assign _T_60775 = select_10 == 6'h5; // @[Switch.scala 41:52:@21934.4]
  assign output_5_10 = io_outValid_10 & _T_60775; // @[Switch.scala 41:38:@21935.4]
  assign _T_60778 = select_11 == 6'h5; // @[Switch.scala 41:52:@21937.4]
  assign output_5_11 = io_outValid_11 & _T_60778; // @[Switch.scala 41:38:@21938.4]
  assign _T_60781 = select_12 == 6'h5; // @[Switch.scala 41:52:@21940.4]
  assign output_5_12 = io_outValid_12 & _T_60781; // @[Switch.scala 41:38:@21941.4]
  assign _T_60784 = select_13 == 6'h5; // @[Switch.scala 41:52:@21943.4]
  assign output_5_13 = io_outValid_13 & _T_60784; // @[Switch.scala 41:38:@21944.4]
  assign _T_60787 = select_14 == 6'h5; // @[Switch.scala 41:52:@21946.4]
  assign output_5_14 = io_outValid_14 & _T_60787; // @[Switch.scala 41:38:@21947.4]
  assign _T_60790 = select_15 == 6'h5; // @[Switch.scala 41:52:@21949.4]
  assign output_5_15 = io_outValid_15 & _T_60790; // @[Switch.scala 41:38:@21950.4]
  assign _T_60793 = select_16 == 6'h5; // @[Switch.scala 41:52:@21952.4]
  assign output_5_16 = io_outValid_16 & _T_60793; // @[Switch.scala 41:38:@21953.4]
  assign _T_60796 = select_17 == 6'h5; // @[Switch.scala 41:52:@21955.4]
  assign output_5_17 = io_outValid_17 & _T_60796; // @[Switch.scala 41:38:@21956.4]
  assign _T_60799 = select_18 == 6'h5; // @[Switch.scala 41:52:@21958.4]
  assign output_5_18 = io_outValid_18 & _T_60799; // @[Switch.scala 41:38:@21959.4]
  assign _T_60802 = select_19 == 6'h5; // @[Switch.scala 41:52:@21961.4]
  assign output_5_19 = io_outValid_19 & _T_60802; // @[Switch.scala 41:38:@21962.4]
  assign _T_60805 = select_20 == 6'h5; // @[Switch.scala 41:52:@21964.4]
  assign output_5_20 = io_outValid_20 & _T_60805; // @[Switch.scala 41:38:@21965.4]
  assign _T_60808 = select_21 == 6'h5; // @[Switch.scala 41:52:@21967.4]
  assign output_5_21 = io_outValid_21 & _T_60808; // @[Switch.scala 41:38:@21968.4]
  assign _T_60811 = select_22 == 6'h5; // @[Switch.scala 41:52:@21970.4]
  assign output_5_22 = io_outValid_22 & _T_60811; // @[Switch.scala 41:38:@21971.4]
  assign _T_60814 = select_23 == 6'h5; // @[Switch.scala 41:52:@21973.4]
  assign output_5_23 = io_outValid_23 & _T_60814; // @[Switch.scala 41:38:@21974.4]
  assign _T_60817 = select_24 == 6'h5; // @[Switch.scala 41:52:@21976.4]
  assign output_5_24 = io_outValid_24 & _T_60817; // @[Switch.scala 41:38:@21977.4]
  assign _T_60820 = select_25 == 6'h5; // @[Switch.scala 41:52:@21979.4]
  assign output_5_25 = io_outValid_25 & _T_60820; // @[Switch.scala 41:38:@21980.4]
  assign _T_60823 = select_26 == 6'h5; // @[Switch.scala 41:52:@21982.4]
  assign output_5_26 = io_outValid_26 & _T_60823; // @[Switch.scala 41:38:@21983.4]
  assign _T_60826 = select_27 == 6'h5; // @[Switch.scala 41:52:@21985.4]
  assign output_5_27 = io_outValid_27 & _T_60826; // @[Switch.scala 41:38:@21986.4]
  assign _T_60829 = select_28 == 6'h5; // @[Switch.scala 41:52:@21988.4]
  assign output_5_28 = io_outValid_28 & _T_60829; // @[Switch.scala 41:38:@21989.4]
  assign _T_60832 = select_29 == 6'h5; // @[Switch.scala 41:52:@21991.4]
  assign output_5_29 = io_outValid_29 & _T_60832; // @[Switch.scala 41:38:@21992.4]
  assign _T_60835 = select_30 == 6'h5; // @[Switch.scala 41:52:@21994.4]
  assign output_5_30 = io_outValid_30 & _T_60835; // @[Switch.scala 41:38:@21995.4]
  assign _T_60838 = select_31 == 6'h5; // @[Switch.scala 41:52:@21997.4]
  assign output_5_31 = io_outValid_31 & _T_60838; // @[Switch.scala 41:38:@21998.4]
  assign _T_60841 = select_32 == 6'h5; // @[Switch.scala 41:52:@22000.4]
  assign output_5_32 = io_outValid_32 & _T_60841; // @[Switch.scala 41:38:@22001.4]
  assign _T_60844 = select_33 == 6'h5; // @[Switch.scala 41:52:@22003.4]
  assign output_5_33 = io_outValid_33 & _T_60844; // @[Switch.scala 41:38:@22004.4]
  assign _T_60847 = select_34 == 6'h5; // @[Switch.scala 41:52:@22006.4]
  assign output_5_34 = io_outValid_34 & _T_60847; // @[Switch.scala 41:38:@22007.4]
  assign _T_60850 = select_35 == 6'h5; // @[Switch.scala 41:52:@22009.4]
  assign output_5_35 = io_outValid_35 & _T_60850; // @[Switch.scala 41:38:@22010.4]
  assign _T_60853 = select_36 == 6'h5; // @[Switch.scala 41:52:@22012.4]
  assign output_5_36 = io_outValid_36 & _T_60853; // @[Switch.scala 41:38:@22013.4]
  assign _T_60856 = select_37 == 6'h5; // @[Switch.scala 41:52:@22015.4]
  assign output_5_37 = io_outValid_37 & _T_60856; // @[Switch.scala 41:38:@22016.4]
  assign _T_60859 = select_38 == 6'h5; // @[Switch.scala 41:52:@22018.4]
  assign output_5_38 = io_outValid_38 & _T_60859; // @[Switch.scala 41:38:@22019.4]
  assign _T_60862 = select_39 == 6'h5; // @[Switch.scala 41:52:@22021.4]
  assign output_5_39 = io_outValid_39 & _T_60862; // @[Switch.scala 41:38:@22022.4]
  assign _T_60865 = select_40 == 6'h5; // @[Switch.scala 41:52:@22024.4]
  assign output_5_40 = io_outValid_40 & _T_60865; // @[Switch.scala 41:38:@22025.4]
  assign _T_60868 = select_41 == 6'h5; // @[Switch.scala 41:52:@22027.4]
  assign output_5_41 = io_outValid_41 & _T_60868; // @[Switch.scala 41:38:@22028.4]
  assign _T_60871 = select_42 == 6'h5; // @[Switch.scala 41:52:@22030.4]
  assign output_5_42 = io_outValid_42 & _T_60871; // @[Switch.scala 41:38:@22031.4]
  assign _T_60874 = select_43 == 6'h5; // @[Switch.scala 41:52:@22033.4]
  assign output_5_43 = io_outValid_43 & _T_60874; // @[Switch.scala 41:38:@22034.4]
  assign _T_60877 = select_44 == 6'h5; // @[Switch.scala 41:52:@22036.4]
  assign output_5_44 = io_outValid_44 & _T_60877; // @[Switch.scala 41:38:@22037.4]
  assign _T_60880 = select_45 == 6'h5; // @[Switch.scala 41:52:@22039.4]
  assign output_5_45 = io_outValid_45 & _T_60880; // @[Switch.scala 41:38:@22040.4]
  assign _T_60883 = select_46 == 6'h5; // @[Switch.scala 41:52:@22042.4]
  assign output_5_46 = io_outValid_46 & _T_60883; // @[Switch.scala 41:38:@22043.4]
  assign _T_60886 = select_47 == 6'h5; // @[Switch.scala 41:52:@22045.4]
  assign output_5_47 = io_outValid_47 & _T_60886; // @[Switch.scala 41:38:@22046.4]
  assign _T_60889 = select_48 == 6'h5; // @[Switch.scala 41:52:@22048.4]
  assign output_5_48 = io_outValid_48 & _T_60889; // @[Switch.scala 41:38:@22049.4]
  assign _T_60892 = select_49 == 6'h5; // @[Switch.scala 41:52:@22051.4]
  assign output_5_49 = io_outValid_49 & _T_60892; // @[Switch.scala 41:38:@22052.4]
  assign _T_60895 = select_50 == 6'h5; // @[Switch.scala 41:52:@22054.4]
  assign output_5_50 = io_outValid_50 & _T_60895; // @[Switch.scala 41:38:@22055.4]
  assign _T_60898 = select_51 == 6'h5; // @[Switch.scala 41:52:@22057.4]
  assign output_5_51 = io_outValid_51 & _T_60898; // @[Switch.scala 41:38:@22058.4]
  assign _T_60901 = select_52 == 6'h5; // @[Switch.scala 41:52:@22060.4]
  assign output_5_52 = io_outValid_52 & _T_60901; // @[Switch.scala 41:38:@22061.4]
  assign _T_60904 = select_53 == 6'h5; // @[Switch.scala 41:52:@22063.4]
  assign output_5_53 = io_outValid_53 & _T_60904; // @[Switch.scala 41:38:@22064.4]
  assign _T_60907 = select_54 == 6'h5; // @[Switch.scala 41:52:@22066.4]
  assign output_5_54 = io_outValid_54 & _T_60907; // @[Switch.scala 41:38:@22067.4]
  assign _T_60910 = select_55 == 6'h5; // @[Switch.scala 41:52:@22069.4]
  assign output_5_55 = io_outValid_55 & _T_60910; // @[Switch.scala 41:38:@22070.4]
  assign _T_60913 = select_56 == 6'h5; // @[Switch.scala 41:52:@22072.4]
  assign output_5_56 = io_outValid_56 & _T_60913; // @[Switch.scala 41:38:@22073.4]
  assign _T_60916 = select_57 == 6'h5; // @[Switch.scala 41:52:@22075.4]
  assign output_5_57 = io_outValid_57 & _T_60916; // @[Switch.scala 41:38:@22076.4]
  assign _T_60919 = select_58 == 6'h5; // @[Switch.scala 41:52:@22078.4]
  assign output_5_58 = io_outValid_58 & _T_60919; // @[Switch.scala 41:38:@22079.4]
  assign _T_60922 = select_59 == 6'h5; // @[Switch.scala 41:52:@22081.4]
  assign output_5_59 = io_outValid_59 & _T_60922; // @[Switch.scala 41:38:@22082.4]
  assign _T_60925 = select_60 == 6'h5; // @[Switch.scala 41:52:@22084.4]
  assign output_5_60 = io_outValid_60 & _T_60925; // @[Switch.scala 41:38:@22085.4]
  assign _T_60928 = select_61 == 6'h5; // @[Switch.scala 41:52:@22087.4]
  assign output_5_61 = io_outValid_61 & _T_60928; // @[Switch.scala 41:38:@22088.4]
  assign _T_60931 = select_62 == 6'h5; // @[Switch.scala 41:52:@22090.4]
  assign output_5_62 = io_outValid_62 & _T_60931; // @[Switch.scala 41:38:@22091.4]
  assign _T_60934 = select_63 == 6'h5; // @[Switch.scala 41:52:@22093.4]
  assign output_5_63 = io_outValid_63 & _T_60934; // @[Switch.scala 41:38:@22094.4]
  assign _T_60942 = {output_5_7,output_5_6,output_5_5,output_5_4,output_5_3,output_5_2,output_5_1,output_5_0}; // @[Switch.scala 43:31:@22102.4]
  assign _T_60950 = {output_5_15,output_5_14,output_5_13,output_5_12,output_5_11,output_5_10,output_5_9,output_5_8,_T_60942}; // @[Switch.scala 43:31:@22110.4]
  assign _T_60957 = {output_5_23,output_5_22,output_5_21,output_5_20,output_5_19,output_5_18,output_5_17,output_5_16}; // @[Switch.scala 43:31:@22117.4]
  assign _T_60966 = {output_5_31,output_5_30,output_5_29,output_5_28,output_5_27,output_5_26,output_5_25,output_5_24,_T_60957,_T_60950}; // @[Switch.scala 43:31:@22126.4]
  assign _T_60973 = {output_5_39,output_5_38,output_5_37,output_5_36,output_5_35,output_5_34,output_5_33,output_5_32}; // @[Switch.scala 43:31:@22133.4]
  assign _T_60981 = {output_5_47,output_5_46,output_5_45,output_5_44,output_5_43,output_5_42,output_5_41,output_5_40,_T_60973}; // @[Switch.scala 43:31:@22141.4]
  assign _T_60988 = {output_5_55,output_5_54,output_5_53,output_5_52,output_5_51,output_5_50,output_5_49,output_5_48}; // @[Switch.scala 43:31:@22148.4]
  assign _T_60997 = {output_5_63,output_5_62,output_5_61,output_5_60,output_5_59,output_5_58,output_5_57,output_5_56,_T_60988,_T_60981}; // @[Switch.scala 43:31:@22157.4]
  assign _T_60998 = {_T_60997,_T_60966}; // @[Switch.scala 43:31:@22158.4]
  assign _T_61002 = select_0 == 6'h6; // @[Switch.scala 41:52:@22161.4]
  assign output_6_0 = io_outValid_0 & _T_61002; // @[Switch.scala 41:38:@22162.4]
  assign _T_61005 = select_1 == 6'h6; // @[Switch.scala 41:52:@22164.4]
  assign output_6_1 = io_outValid_1 & _T_61005; // @[Switch.scala 41:38:@22165.4]
  assign _T_61008 = select_2 == 6'h6; // @[Switch.scala 41:52:@22167.4]
  assign output_6_2 = io_outValid_2 & _T_61008; // @[Switch.scala 41:38:@22168.4]
  assign _T_61011 = select_3 == 6'h6; // @[Switch.scala 41:52:@22170.4]
  assign output_6_3 = io_outValid_3 & _T_61011; // @[Switch.scala 41:38:@22171.4]
  assign _T_61014 = select_4 == 6'h6; // @[Switch.scala 41:52:@22173.4]
  assign output_6_4 = io_outValid_4 & _T_61014; // @[Switch.scala 41:38:@22174.4]
  assign _T_61017 = select_5 == 6'h6; // @[Switch.scala 41:52:@22176.4]
  assign output_6_5 = io_outValid_5 & _T_61017; // @[Switch.scala 41:38:@22177.4]
  assign _T_61020 = select_6 == 6'h6; // @[Switch.scala 41:52:@22179.4]
  assign output_6_6 = io_outValid_6 & _T_61020; // @[Switch.scala 41:38:@22180.4]
  assign _T_61023 = select_7 == 6'h6; // @[Switch.scala 41:52:@22182.4]
  assign output_6_7 = io_outValid_7 & _T_61023; // @[Switch.scala 41:38:@22183.4]
  assign _T_61026 = select_8 == 6'h6; // @[Switch.scala 41:52:@22185.4]
  assign output_6_8 = io_outValid_8 & _T_61026; // @[Switch.scala 41:38:@22186.4]
  assign _T_61029 = select_9 == 6'h6; // @[Switch.scala 41:52:@22188.4]
  assign output_6_9 = io_outValid_9 & _T_61029; // @[Switch.scala 41:38:@22189.4]
  assign _T_61032 = select_10 == 6'h6; // @[Switch.scala 41:52:@22191.4]
  assign output_6_10 = io_outValid_10 & _T_61032; // @[Switch.scala 41:38:@22192.4]
  assign _T_61035 = select_11 == 6'h6; // @[Switch.scala 41:52:@22194.4]
  assign output_6_11 = io_outValid_11 & _T_61035; // @[Switch.scala 41:38:@22195.4]
  assign _T_61038 = select_12 == 6'h6; // @[Switch.scala 41:52:@22197.4]
  assign output_6_12 = io_outValid_12 & _T_61038; // @[Switch.scala 41:38:@22198.4]
  assign _T_61041 = select_13 == 6'h6; // @[Switch.scala 41:52:@22200.4]
  assign output_6_13 = io_outValid_13 & _T_61041; // @[Switch.scala 41:38:@22201.4]
  assign _T_61044 = select_14 == 6'h6; // @[Switch.scala 41:52:@22203.4]
  assign output_6_14 = io_outValid_14 & _T_61044; // @[Switch.scala 41:38:@22204.4]
  assign _T_61047 = select_15 == 6'h6; // @[Switch.scala 41:52:@22206.4]
  assign output_6_15 = io_outValid_15 & _T_61047; // @[Switch.scala 41:38:@22207.4]
  assign _T_61050 = select_16 == 6'h6; // @[Switch.scala 41:52:@22209.4]
  assign output_6_16 = io_outValid_16 & _T_61050; // @[Switch.scala 41:38:@22210.4]
  assign _T_61053 = select_17 == 6'h6; // @[Switch.scala 41:52:@22212.4]
  assign output_6_17 = io_outValid_17 & _T_61053; // @[Switch.scala 41:38:@22213.4]
  assign _T_61056 = select_18 == 6'h6; // @[Switch.scala 41:52:@22215.4]
  assign output_6_18 = io_outValid_18 & _T_61056; // @[Switch.scala 41:38:@22216.4]
  assign _T_61059 = select_19 == 6'h6; // @[Switch.scala 41:52:@22218.4]
  assign output_6_19 = io_outValid_19 & _T_61059; // @[Switch.scala 41:38:@22219.4]
  assign _T_61062 = select_20 == 6'h6; // @[Switch.scala 41:52:@22221.4]
  assign output_6_20 = io_outValid_20 & _T_61062; // @[Switch.scala 41:38:@22222.4]
  assign _T_61065 = select_21 == 6'h6; // @[Switch.scala 41:52:@22224.4]
  assign output_6_21 = io_outValid_21 & _T_61065; // @[Switch.scala 41:38:@22225.4]
  assign _T_61068 = select_22 == 6'h6; // @[Switch.scala 41:52:@22227.4]
  assign output_6_22 = io_outValid_22 & _T_61068; // @[Switch.scala 41:38:@22228.4]
  assign _T_61071 = select_23 == 6'h6; // @[Switch.scala 41:52:@22230.4]
  assign output_6_23 = io_outValid_23 & _T_61071; // @[Switch.scala 41:38:@22231.4]
  assign _T_61074 = select_24 == 6'h6; // @[Switch.scala 41:52:@22233.4]
  assign output_6_24 = io_outValid_24 & _T_61074; // @[Switch.scala 41:38:@22234.4]
  assign _T_61077 = select_25 == 6'h6; // @[Switch.scala 41:52:@22236.4]
  assign output_6_25 = io_outValid_25 & _T_61077; // @[Switch.scala 41:38:@22237.4]
  assign _T_61080 = select_26 == 6'h6; // @[Switch.scala 41:52:@22239.4]
  assign output_6_26 = io_outValid_26 & _T_61080; // @[Switch.scala 41:38:@22240.4]
  assign _T_61083 = select_27 == 6'h6; // @[Switch.scala 41:52:@22242.4]
  assign output_6_27 = io_outValid_27 & _T_61083; // @[Switch.scala 41:38:@22243.4]
  assign _T_61086 = select_28 == 6'h6; // @[Switch.scala 41:52:@22245.4]
  assign output_6_28 = io_outValid_28 & _T_61086; // @[Switch.scala 41:38:@22246.4]
  assign _T_61089 = select_29 == 6'h6; // @[Switch.scala 41:52:@22248.4]
  assign output_6_29 = io_outValid_29 & _T_61089; // @[Switch.scala 41:38:@22249.4]
  assign _T_61092 = select_30 == 6'h6; // @[Switch.scala 41:52:@22251.4]
  assign output_6_30 = io_outValid_30 & _T_61092; // @[Switch.scala 41:38:@22252.4]
  assign _T_61095 = select_31 == 6'h6; // @[Switch.scala 41:52:@22254.4]
  assign output_6_31 = io_outValid_31 & _T_61095; // @[Switch.scala 41:38:@22255.4]
  assign _T_61098 = select_32 == 6'h6; // @[Switch.scala 41:52:@22257.4]
  assign output_6_32 = io_outValid_32 & _T_61098; // @[Switch.scala 41:38:@22258.4]
  assign _T_61101 = select_33 == 6'h6; // @[Switch.scala 41:52:@22260.4]
  assign output_6_33 = io_outValid_33 & _T_61101; // @[Switch.scala 41:38:@22261.4]
  assign _T_61104 = select_34 == 6'h6; // @[Switch.scala 41:52:@22263.4]
  assign output_6_34 = io_outValid_34 & _T_61104; // @[Switch.scala 41:38:@22264.4]
  assign _T_61107 = select_35 == 6'h6; // @[Switch.scala 41:52:@22266.4]
  assign output_6_35 = io_outValid_35 & _T_61107; // @[Switch.scala 41:38:@22267.4]
  assign _T_61110 = select_36 == 6'h6; // @[Switch.scala 41:52:@22269.4]
  assign output_6_36 = io_outValid_36 & _T_61110; // @[Switch.scala 41:38:@22270.4]
  assign _T_61113 = select_37 == 6'h6; // @[Switch.scala 41:52:@22272.4]
  assign output_6_37 = io_outValid_37 & _T_61113; // @[Switch.scala 41:38:@22273.4]
  assign _T_61116 = select_38 == 6'h6; // @[Switch.scala 41:52:@22275.4]
  assign output_6_38 = io_outValid_38 & _T_61116; // @[Switch.scala 41:38:@22276.4]
  assign _T_61119 = select_39 == 6'h6; // @[Switch.scala 41:52:@22278.4]
  assign output_6_39 = io_outValid_39 & _T_61119; // @[Switch.scala 41:38:@22279.4]
  assign _T_61122 = select_40 == 6'h6; // @[Switch.scala 41:52:@22281.4]
  assign output_6_40 = io_outValid_40 & _T_61122; // @[Switch.scala 41:38:@22282.4]
  assign _T_61125 = select_41 == 6'h6; // @[Switch.scala 41:52:@22284.4]
  assign output_6_41 = io_outValid_41 & _T_61125; // @[Switch.scala 41:38:@22285.4]
  assign _T_61128 = select_42 == 6'h6; // @[Switch.scala 41:52:@22287.4]
  assign output_6_42 = io_outValid_42 & _T_61128; // @[Switch.scala 41:38:@22288.4]
  assign _T_61131 = select_43 == 6'h6; // @[Switch.scala 41:52:@22290.4]
  assign output_6_43 = io_outValid_43 & _T_61131; // @[Switch.scala 41:38:@22291.4]
  assign _T_61134 = select_44 == 6'h6; // @[Switch.scala 41:52:@22293.4]
  assign output_6_44 = io_outValid_44 & _T_61134; // @[Switch.scala 41:38:@22294.4]
  assign _T_61137 = select_45 == 6'h6; // @[Switch.scala 41:52:@22296.4]
  assign output_6_45 = io_outValid_45 & _T_61137; // @[Switch.scala 41:38:@22297.4]
  assign _T_61140 = select_46 == 6'h6; // @[Switch.scala 41:52:@22299.4]
  assign output_6_46 = io_outValid_46 & _T_61140; // @[Switch.scala 41:38:@22300.4]
  assign _T_61143 = select_47 == 6'h6; // @[Switch.scala 41:52:@22302.4]
  assign output_6_47 = io_outValid_47 & _T_61143; // @[Switch.scala 41:38:@22303.4]
  assign _T_61146 = select_48 == 6'h6; // @[Switch.scala 41:52:@22305.4]
  assign output_6_48 = io_outValid_48 & _T_61146; // @[Switch.scala 41:38:@22306.4]
  assign _T_61149 = select_49 == 6'h6; // @[Switch.scala 41:52:@22308.4]
  assign output_6_49 = io_outValid_49 & _T_61149; // @[Switch.scala 41:38:@22309.4]
  assign _T_61152 = select_50 == 6'h6; // @[Switch.scala 41:52:@22311.4]
  assign output_6_50 = io_outValid_50 & _T_61152; // @[Switch.scala 41:38:@22312.4]
  assign _T_61155 = select_51 == 6'h6; // @[Switch.scala 41:52:@22314.4]
  assign output_6_51 = io_outValid_51 & _T_61155; // @[Switch.scala 41:38:@22315.4]
  assign _T_61158 = select_52 == 6'h6; // @[Switch.scala 41:52:@22317.4]
  assign output_6_52 = io_outValid_52 & _T_61158; // @[Switch.scala 41:38:@22318.4]
  assign _T_61161 = select_53 == 6'h6; // @[Switch.scala 41:52:@22320.4]
  assign output_6_53 = io_outValid_53 & _T_61161; // @[Switch.scala 41:38:@22321.4]
  assign _T_61164 = select_54 == 6'h6; // @[Switch.scala 41:52:@22323.4]
  assign output_6_54 = io_outValid_54 & _T_61164; // @[Switch.scala 41:38:@22324.4]
  assign _T_61167 = select_55 == 6'h6; // @[Switch.scala 41:52:@22326.4]
  assign output_6_55 = io_outValid_55 & _T_61167; // @[Switch.scala 41:38:@22327.4]
  assign _T_61170 = select_56 == 6'h6; // @[Switch.scala 41:52:@22329.4]
  assign output_6_56 = io_outValid_56 & _T_61170; // @[Switch.scala 41:38:@22330.4]
  assign _T_61173 = select_57 == 6'h6; // @[Switch.scala 41:52:@22332.4]
  assign output_6_57 = io_outValid_57 & _T_61173; // @[Switch.scala 41:38:@22333.4]
  assign _T_61176 = select_58 == 6'h6; // @[Switch.scala 41:52:@22335.4]
  assign output_6_58 = io_outValid_58 & _T_61176; // @[Switch.scala 41:38:@22336.4]
  assign _T_61179 = select_59 == 6'h6; // @[Switch.scala 41:52:@22338.4]
  assign output_6_59 = io_outValid_59 & _T_61179; // @[Switch.scala 41:38:@22339.4]
  assign _T_61182 = select_60 == 6'h6; // @[Switch.scala 41:52:@22341.4]
  assign output_6_60 = io_outValid_60 & _T_61182; // @[Switch.scala 41:38:@22342.4]
  assign _T_61185 = select_61 == 6'h6; // @[Switch.scala 41:52:@22344.4]
  assign output_6_61 = io_outValid_61 & _T_61185; // @[Switch.scala 41:38:@22345.4]
  assign _T_61188 = select_62 == 6'h6; // @[Switch.scala 41:52:@22347.4]
  assign output_6_62 = io_outValid_62 & _T_61188; // @[Switch.scala 41:38:@22348.4]
  assign _T_61191 = select_63 == 6'h6; // @[Switch.scala 41:52:@22350.4]
  assign output_6_63 = io_outValid_63 & _T_61191; // @[Switch.scala 41:38:@22351.4]
  assign _T_61199 = {output_6_7,output_6_6,output_6_5,output_6_4,output_6_3,output_6_2,output_6_1,output_6_0}; // @[Switch.scala 43:31:@22359.4]
  assign _T_61207 = {output_6_15,output_6_14,output_6_13,output_6_12,output_6_11,output_6_10,output_6_9,output_6_8,_T_61199}; // @[Switch.scala 43:31:@22367.4]
  assign _T_61214 = {output_6_23,output_6_22,output_6_21,output_6_20,output_6_19,output_6_18,output_6_17,output_6_16}; // @[Switch.scala 43:31:@22374.4]
  assign _T_61223 = {output_6_31,output_6_30,output_6_29,output_6_28,output_6_27,output_6_26,output_6_25,output_6_24,_T_61214,_T_61207}; // @[Switch.scala 43:31:@22383.4]
  assign _T_61230 = {output_6_39,output_6_38,output_6_37,output_6_36,output_6_35,output_6_34,output_6_33,output_6_32}; // @[Switch.scala 43:31:@22390.4]
  assign _T_61238 = {output_6_47,output_6_46,output_6_45,output_6_44,output_6_43,output_6_42,output_6_41,output_6_40,_T_61230}; // @[Switch.scala 43:31:@22398.4]
  assign _T_61245 = {output_6_55,output_6_54,output_6_53,output_6_52,output_6_51,output_6_50,output_6_49,output_6_48}; // @[Switch.scala 43:31:@22405.4]
  assign _T_61254 = {output_6_63,output_6_62,output_6_61,output_6_60,output_6_59,output_6_58,output_6_57,output_6_56,_T_61245,_T_61238}; // @[Switch.scala 43:31:@22414.4]
  assign _T_61255 = {_T_61254,_T_61223}; // @[Switch.scala 43:31:@22415.4]
  assign _T_61259 = select_0 == 6'h7; // @[Switch.scala 41:52:@22418.4]
  assign output_7_0 = io_outValid_0 & _T_61259; // @[Switch.scala 41:38:@22419.4]
  assign _T_61262 = select_1 == 6'h7; // @[Switch.scala 41:52:@22421.4]
  assign output_7_1 = io_outValid_1 & _T_61262; // @[Switch.scala 41:38:@22422.4]
  assign _T_61265 = select_2 == 6'h7; // @[Switch.scala 41:52:@22424.4]
  assign output_7_2 = io_outValid_2 & _T_61265; // @[Switch.scala 41:38:@22425.4]
  assign _T_61268 = select_3 == 6'h7; // @[Switch.scala 41:52:@22427.4]
  assign output_7_3 = io_outValid_3 & _T_61268; // @[Switch.scala 41:38:@22428.4]
  assign _T_61271 = select_4 == 6'h7; // @[Switch.scala 41:52:@22430.4]
  assign output_7_4 = io_outValid_4 & _T_61271; // @[Switch.scala 41:38:@22431.4]
  assign _T_61274 = select_5 == 6'h7; // @[Switch.scala 41:52:@22433.4]
  assign output_7_5 = io_outValid_5 & _T_61274; // @[Switch.scala 41:38:@22434.4]
  assign _T_61277 = select_6 == 6'h7; // @[Switch.scala 41:52:@22436.4]
  assign output_7_6 = io_outValid_6 & _T_61277; // @[Switch.scala 41:38:@22437.4]
  assign _T_61280 = select_7 == 6'h7; // @[Switch.scala 41:52:@22439.4]
  assign output_7_7 = io_outValid_7 & _T_61280; // @[Switch.scala 41:38:@22440.4]
  assign _T_61283 = select_8 == 6'h7; // @[Switch.scala 41:52:@22442.4]
  assign output_7_8 = io_outValid_8 & _T_61283; // @[Switch.scala 41:38:@22443.4]
  assign _T_61286 = select_9 == 6'h7; // @[Switch.scala 41:52:@22445.4]
  assign output_7_9 = io_outValid_9 & _T_61286; // @[Switch.scala 41:38:@22446.4]
  assign _T_61289 = select_10 == 6'h7; // @[Switch.scala 41:52:@22448.4]
  assign output_7_10 = io_outValid_10 & _T_61289; // @[Switch.scala 41:38:@22449.4]
  assign _T_61292 = select_11 == 6'h7; // @[Switch.scala 41:52:@22451.4]
  assign output_7_11 = io_outValid_11 & _T_61292; // @[Switch.scala 41:38:@22452.4]
  assign _T_61295 = select_12 == 6'h7; // @[Switch.scala 41:52:@22454.4]
  assign output_7_12 = io_outValid_12 & _T_61295; // @[Switch.scala 41:38:@22455.4]
  assign _T_61298 = select_13 == 6'h7; // @[Switch.scala 41:52:@22457.4]
  assign output_7_13 = io_outValid_13 & _T_61298; // @[Switch.scala 41:38:@22458.4]
  assign _T_61301 = select_14 == 6'h7; // @[Switch.scala 41:52:@22460.4]
  assign output_7_14 = io_outValid_14 & _T_61301; // @[Switch.scala 41:38:@22461.4]
  assign _T_61304 = select_15 == 6'h7; // @[Switch.scala 41:52:@22463.4]
  assign output_7_15 = io_outValid_15 & _T_61304; // @[Switch.scala 41:38:@22464.4]
  assign _T_61307 = select_16 == 6'h7; // @[Switch.scala 41:52:@22466.4]
  assign output_7_16 = io_outValid_16 & _T_61307; // @[Switch.scala 41:38:@22467.4]
  assign _T_61310 = select_17 == 6'h7; // @[Switch.scala 41:52:@22469.4]
  assign output_7_17 = io_outValid_17 & _T_61310; // @[Switch.scala 41:38:@22470.4]
  assign _T_61313 = select_18 == 6'h7; // @[Switch.scala 41:52:@22472.4]
  assign output_7_18 = io_outValid_18 & _T_61313; // @[Switch.scala 41:38:@22473.4]
  assign _T_61316 = select_19 == 6'h7; // @[Switch.scala 41:52:@22475.4]
  assign output_7_19 = io_outValid_19 & _T_61316; // @[Switch.scala 41:38:@22476.4]
  assign _T_61319 = select_20 == 6'h7; // @[Switch.scala 41:52:@22478.4]
  assign output_7_20 = io_outValid_20 & _T_61319; // @[Switch.scala 41:38:@22479.4]
  assign _T_61322 = select_21 == 6'h7; // @[Switch.scala 41:52:@22481.4]
  assign output_7_21 = io_outValid_21 & _T_61322; // @[Switch.scala 41:38:@22482.4]
  assign _T_61325 = select_22 == 6'h7; // @[Switch.scala 41:52:@22484.4]
  assign output_7_22 = io_outValid_22 & _T_61325; // @[Switch.scala 41:38:@22485.4]
  assign _T_61328 = select_23 == 6'h7; // @[Switch.scala 41:52:@22487.4]
  assign output_7_23 = io_outValid_23 & _T_61328; // @[Switch.scala 41:38:@22488.4]
  assign _T_61331 = select_24 == 6'h7; // @[Switch.scala 41:52:@22490.4]
  assign output_7_24 = io_outValid_24 & _T_61331; // @[Switch.scala 41:38:@22491.4]
  assign _T_61334 = select_25 == 6'h7; // @[Switch.scala 41:52:@22493.4]
  assign output_7_25 = io_outValid_25 & _T_61334; // @[Switch.scala 41:38:@22494.4]
  assign _T_61337 = select_26 == 6'h7; // @[Switch.scala 41:52:@22496.4]
  assign output_7_26 = io_outValid_26 & _T_61337; // @[Switch.scala 41:38:@22497.4]
  assign _T_61340 = select_27 == 6'h7; // @[Switch.scala 41:52:@22499.4]
  assign output_7_27 = io_outValid_27 & _T_61340; // @[Switch.scala 41:38:@22500.4]
  assign _T_61343 = select_28 == 6'h7; // @[Switch.scala 41:52:@22502.4]
  assign output_7_28 = io_outValid_28 & _T_61343; // @[Switch.scala 41:38:@22503.4]
  assign _T_61346 = select_29 == 6'h7; // @[Switch.scala 41:52:@22505.4]
  assign output_7_29 = io_outValid_29 & _T_61346; // @[Switch.scala 41:38:@22506.4]
  assign _T_61349 = select_30 == 6'h7; // @[Switch.scala 41:52:@22508.4]
  assign output_7_30 = io_outValid_30 & _T_61349; // @[Switch.scala 41:38:@22509.4]
  assign _T_61352 = select_31 == 6'h7; // @[Switch.scala 41:52:@22511.4]
  assign output_7_31 = io_outValid_31 & _T_61352; // @[Switch.scala 41:38:@22512.4]
  assign _T_61355 = select_32 == 6'h7; // @[Switch.scala 41:52:@22514.4]
  assign output_7_32 = io_outValid_32 & _T_61355; // @[Switch.scala 41:38:@22515.4]
  assign _T_61358 = select_33 == 6'h7; // @[Switch.scala 41:52:@22517.4]
  assign output_7_33 = io_outValid_33 & _T_61358; // @[Switch.scala 41:38:@22518.4]
  assign _T_61361 = select_34 == 6'h7; // @[Switch.scala 41:52:@22520.4]
  assign output_7_34 = io_outValid_34 & _T_61361; // @[Switch.scala 41:38:@22521.4]
  assign _T_61364 = select_35 == 6'h7; // @[Switch.scala 41:52:@22523.4]
  assign output_7_35 = io_outValid_35 & _T_61364; // @[Switch.scala 41:38:@22524.4]
  assign _T_61367 = select_36 == 6'h7; // @[Switch.scala 41:52:@22526.4]
  assign output_7_36 = io_outValid_36 & _T_61367; // @[Switch.scala 41:38:@22527.4]
  assign _T_61370 = select_37 == 6'h7; // @[Switch.scala 41:52:@22529.4]
  assign output_7_37 = io_outValid_37 & _T_61370; // @[Switch.scala 41:38:@22530.4]
  assign _T_61373 = select_38 == 6'h7; // @[Switch.scala 41:52:@22532.4]
  assign output_7_38 = io_outValid_38 & _T_61373; // @[Switch.scala 41:38:@22533.4]
  assign _T_61376 = select_39 == 6'h7; // @[Switch.scala 41:52:@22535.4]
  assign output_7_39 = io_outValid_39 & _T_61376; // @[Switch.scala 41:38:@22536.4]
  assign _T_61379 = select_40 == 6'h7; // @[Switch.scala 41:52:@22538.4]
  assign output_7_40 = io_outValid_40 & _T_61379; // @[Switch.scala 41:38:@22539.4]
  assign _T_61382 = select_41 == 6'h7; // @[Switch.scala 41:52:@22541.4]
  assign output_7_41 = io_outValid_41 & _T_61382; // @[Switch.scala 41:38:@22542.4]
  assign _T_61385 = select_42 == 6'h7; // @[Switch.scala 41:52:@22544.4]
  assign output_7_42 = io_outValid_42 & _T_61385; // @[Switch.scala 41:38:@22545.4]
  assign _T_61388 = select_43 == 6'h7; // @[Switch.scala 41:52:@22547.4]
  assign output_7_43 = io_outValid_43 & _T_61388; // @[Switch.scala 41:38:@22548.4]
  assign _T_61391 = select_44 == 6'h7; // @[Switch.scala 41:52:@22550.4]
  assign output_7_44 = io_outValid_44 & _T_61391; // @[Switch.scala 41:38:@22551.4]
  assign _T_61394 = select_45 == 6'h7; // @[Switch.scala 41:52:@22553.4]
  assign output_7_45 = io_outValid_45 & _T_61394; // @[Switch.scala 41:38:@22554.4]
  assign _T_61397 = select_46 == 6'h7; // @[Switch.scala 41:52:@22556.4]
  assign output_7_46 = io_outValid_46 & _T_61397; // @[Switch.scala 41:38:@22557.4]
  assign _T_61400 = select_47 == 6'h7; // @[Switch.scala 41:52:@22559.4]
  assign output_7_47 = io_outValid_47 & _T_61400; // @[Switch.scala 41:38:@22560.4]
  assign _T_61403 = select_48 == 6'h7; // @[Switch.scala 41:52:@22562.4]
  assign output_7_48 = io_outValid_48 & _T_61403; // @[Switch.scala 41:38:@22563.4]
  assign _T_61406 = select_49 == 6'h7; // @[Switch.scala 41:52:@22565.4]
  assign output_7_49 = io_outValid_49 & _T_61406; // @[Switch.scala 41:38:@22566.4]
  assign _T_61409 = select_50 == 6'h7; // @[Switch.scala 41:52:@22568.4]
  assign output_7_50 = io_outValid_50 & _T_61409; // @[Switch.scala 41:38:@22569.4]
  assign _T_61412 = select_51 == 6'h7; // @[Switch.scala 41:52:@22571.4]
  assign output_7_51 = io_outValid_51 & _T_61412; // @[Switch.scala 41:38:@22572.4]
  assign _T_61415 = select_52 == 6'h7; // @[Switch.scala 41:52:@22574.4]
  assign output_7_52 = io_outValid_52 & _T_61415; // @[Switch.scala 41:38:@22575.4]
  assign _T_61418 = select_53 == 6'h7; // @[Switch.scala 41:52:@22577.4]
  assign output_7_53 = io_outValid_53 & _T_61418; // @[Switch.scala 41:38:@22578.4]
  assign _T_61421 = select_54 == 6'h7; // @[Switch.scala 41:52:@22580.4]
  assign output_7_54 = io_outValid_54 & _T_61421; // @[Switch.scala 41:38:@22581.4]
  assign _T_61424 = select_55 == 6'h7; // @[Switch.scala 41:52:@22583.4]
  assign output_7_55 = io_outValid_55 & _T_61424; // @[Switch.scala 41:38:@22584.4]
  assign _T_61427 = select_56 == 6'h7; // @[Switch.scala 41:52:@22586.4]
  assign output_7_56 = io_outValid_56 & _T_61427; // @[Switch.scala 41:38:@22587.4]
  assign _T_61430 = select_57 == 6'h7; // @[Switch.scala 41:52:@22589.4]
  assign output_7_57 = io_outValid_57 & _T_61430; // @[Switch.scala 41:38:@22590.4]
  assign _T_61433 = select_58 == 6'h7; // @[Switch.scala 41:52:@22592.4]
  assign output_7_58 = io_outValid_58 & _T_61433; // @[Switch.scala 41:38:@22593.4]
  assign _T_61436 = select_59 == 6'h7; // @[Switch.scala 41:52:@22595.4]
  assign output_7_59 = io_outValid_59 & _T_61436; // @[Switch.scala 41:38:@22596.4]
  assign _T_61439 = select_60 == 6'h7; // @[Switch.scala 41:52:@22598.4]
  assign output_7_60 = io_outValid_60 & _T_61439; // @[Switch.scala 41:38:@22599.4]
  assign _T_61442 = select_61 == 6'h7; // @[Switch.scala 41:52:@22601.4]
  assign output_7_61 = io_outValid_61 & _T_61442; // @[Switch.scala 41:38:@22602.4]
  assign _T_61445 = select_62 == 6'h7; // @[Switch.scala 41:52:@22604.4]
  assign output_7_62 = io_outValid_62 & _T_61445; // @[Switch.scala 41:38:@22605.4]
  assign _T_61448 = select_63 == 6'h7; // @[Switch.scala 41:52:@22607.4]
  assign output_7_63 = io_outValid_63 & _T_61448; // @[Switch.scala 41:38:@22608.4]
  assign _T_61456 = {output_7_7,output_7_6,output_7_5,output_7_4,output_7_3,output_7_2,output_7_1,output_7_0}; // @[Switch.scala 43:31:@22616.4]
  assign _T_61464 = {output_7_15,output_7_14,output_7_13,output_7_12,output_7_11,output_7_10,output_7_9,output_7_8,_T_61456}; // @[Switch.scala 43:31:@22624.4]
  assign _T_61471 = {output_7_23,output_7_22,output_7_21,output_7_20,output_7_19,output_7_18,output_7_17,output_7_16}; // @[Switch.scala 43:31:@22631.4]
  assign _T_61480 = {output_7_31,output_7_30,output_7_29,output_7_28,output_7_27,output_7_26,output_7_25,output_7_24,_T_61471,_T_61464}; // @[Switch.scala 43:31:@22640.4]
  assign _T_61487 = {output_7_39,output_7_38,output_7_37,output_7_36,output_7_35,output_7_34,output_7_33,output_7_32}; // @[Switch.scala 43:31:@22647.4]
  assign _T_61495 = {output_7_47,output_7_46,output_7_45,output_7_44,output_7_43,output_7_42,output_7_41,output_7_40,_T_61487}; // @[Switch.scala 43:31:@22655.4]
  assign _T_61502 = {output_7_55,output_7_54,output_7_53,output_7_52,output_7_51,output_7_50,output_7_49,output_7_48}; // @[Switch.scala 43:31:@22662.4]
  assign _T_61511 = {output_7_63,output_7_62,output_7_61,output_7_60,output_7_59,output_7_58,output_7_57,output_7_56,_T_61502,_T_61495}; // @[Switch.scala 43:31:@22671.4]
  assign _T_61512 = {_T_61511,_T_61480}; // @[Switch.scala 43:31:@22672.4]
  assign _T_61516 = select_0 == 6'h8; // @[Switch.scala 41:52:@22675.4]
  assign output_8_0 = io_outValid_0 & _T_61516; // @[Switch.scala 41:38:@22676.4]
  assign _T_61519 = select_1 == 6'h8; // @[Switch.scala 41:52:@22678.4]
  assign output_8_1 = io_outValid_1 & _T_61519; // @[Switch.scala 41:38:@22679.4]
  assign _T_61522 = select_2 == 6'h8; // @[Switch.scala 41:52:@22681.4]
  assign output_8_2 = io_outValid_2 & _T_61522; // @[Switch.scala 41:38:@22682.4]
  assign _T_61525 = select_3 == 6'h8; // @[Switch.scala 41:52:@22684.4]
  assign output_8_3 = io_outValid_3 & _T_61525; // @[Switch.scala 41:38:@22685.4]
  assign _T_61528 = select_4 == 6'h8; // @[Switch.scala 41:52:@22687.4]
  assign output_8_4 = io_outValid_4 & _T_61528; // @[Switch.scala 41:38:@22688.4]
  assign _T_61531 = select_5 == 6'h8; // @[Switch.scala 41:52:@22690.4]
  assign output_8_5 = io_outValid_5 & _T_61531; // @[Switch.scala 41:38:@22691.4]
  assign _T_61534 = select_6 == 6'h8; // @[Switch.scala 41:52:@22693.4]
  assign output_8_6 = io_outValid_6 & _T_61534; // @[Switch.scala 41:38:@22694.4]
  assign _T_61537 = select_7 == 6'h8; // @[Switch.scala 41:52:@22696.4]
  assign output_8_7 = io_outValid_7 & _T_61537; // @[Switch.scala 41:38:@22697.4]
  assign _T_61540 = select_8 == 6'h8; // @[Switch.scala 41:52:@22699.4]
  assign output_8_8 = io_outValid_8 & _T_61540; // @[Switch.scala 41:38:@22700.4]
  assign _T_61543 = select_9 == 6'h8; // @[Switch.scala 41:52:@22702.4]
  assign output_8_9 = io_outValid_9 & _T_61543; // @[Switch.scala 41:38:@22703.4]
  assign _T_61546 = select_10 == 6'h8; // @[Switch.scala 41:52:@22705.4]
  assign output_8_10 = io_outValid_10 & _T_61546; // @[Switch.scala 41:38:@22706.4]
  assign _T_61549 = select_11 == 6'h8; // @[Switch.scala 41:52:@22708.4]
  assign output_8_11 = io_outValid_11 & _T_61549; // @[Switch.scala 41:38:@22709.4]
  assign _T_61552 = select_12 == 6'h8; // @[Switch.scala 41:52:@22711.4]
  assign output_8_12 = io_outValid_12 & _T_61552; // @[Switch.scala 41:38:@22712.4]
  assign _T_61555 = select_13 == 6'h8; // @[Switch.scala 41:52:@22714.4]
  assign output_8_13 = io_outValid_13 & _T_61555; // @[Switch.scala 41:38:@22715.4]
  assign _T_61558 = select_14 == 6'h8; // @[Switch.scala 41:52:@22717.4]
  assign output_8_14 = io_outValid_14 & _T_61558; // @[Switch.scala 41:38:@22718.4]
  assign _T_61561 = select_15 == 6'h8; // @[Switch.scala 41:52:@22720.4]
  assign output_8_15 = io_outValid_15 & _T_61561; // @[Switch.scala 41:38:@22721.4]
  assign _T_61564 = select_16 == 6'h8; // @[Switch.scala 41:52:@22723.4]
  assign output_8_16 = io_outValid_16 & _T_61564; // @[Switch.scala 41:38:@22724.4]
  assign _T_61567 = select_17 == 6'h8; // @[Switch.scala 41:52:@22726.4]
  assign output_8_17 = io_outValid_17 & _T_61567; // @[Switch.scala 41:38:@22727.4]
  assign _T_61570 = select_18 == 6'h8; // @[Switch.scala 41:52:@22729.4]
  assign output_8_18 = io_outValid_18 & _T_61570; // @[Switch.scala 41:38:@22730.4]
  assign _T_61573 = select_19 == 6'h8; // @[Switch.scala 41:52:@22732.4]
  assign output_8_19 = io_outValid_19 & _T_61573; // @[Switch.scala 41:38:@22733.4]
  assign _T_61576 = select_20 == 6'h8; // @[Switch.scala 41:52:@22735.4]
  assign output_8_20 = io_outValid_20 & _T_61576; // @[Switch.scala 41:38:@22736.4]
  assign _T_61579 = select_21 == 6'h8; // @[Switch.scala 41:52:@22738.4]
  assign output_8_21 = io_outValid_21 & _T_61579; // @[Switch.scala 41:38:@22739.4]
  assign _T_61582 = select_22 == 6'h8; // @[Switch.scala 41:52:@22741.4]
  assign output_8_22 = io_outValid_22 & _T_61582; // @[Switch.scala 41:38:@22742.4]
  assign _T_61585 = select_23 == 6'h8; // @[Switch.scala 41:52:@22744.4]
  assign output_8_23 = io_outValid_23 & _T_61585; // @[Switch.scala 41:38:@22745.4]
  assign _T_61588 = select_24 == 6'h8; // @[Switch.scala 41:52:@22747.4]
  assign output_8_24 = io_outValid_24 & _T_61588; // @[Switch.scala 41:38:@22748.4]
  assign _T_61591 = select_25 == 6'h8; // @[Switch.scala 41:52:@22750.4]
  assign output_8_25 = io_outValid_25 & _T_61591; // @[Switch.scala 41:38:@22751.4]
  assign _T_61594 = select_26 == 6'h8; // @[Switch.scala 41:52:@22753.4]
  assign output_8_26 = io_outValid_26 & _T_61594; // @[Switch.scala 41:38:@22754.4]
  assign _T_61597 = select_27 == 6'h8; // @[Switch.scala 41:52:@22756.4]
  assign output_8_27 = io_outValid_27 & _T_61597; // @[Switch.scala 41:38:@22757.4]
  assign _T_61600 = select_28 == 6'h8; // @[Switch.scala 41:52:@22759.4]
  assign output_8_28 = io_outValid_28 & _T_61600; // @[Switch.scala 41:38:@22760.4]
  assign _T_61603 = select_29 == 6'h8; // @[Switch.scala 41:52:@22762.4]
  assign output_8_29 = io_outValid_29 & _T_61603; // @[Switch.scala 41:38:@22763.4]
  assign _T_61606 = select_30 == 6'h8; // @[Switch.scala 41:52:@22765.4]
  assign output_8_30 = io_outValid_30 & _T_61606; // @[Switch.scala 41:38:@22766.4]
  assign _T_61609 = select_31 == 6'h8; // @[Switch.scala 41:52:@22768.4]
  assign output_8_31 = io_outValid_31 & _T_61609; // @[Switch.scala 41:38:@22769.4]
  assign _T_61612 = select_32 == 6'h8; // @[Switch.scala 41:52:@22771.4]
  assign output_8_32 = io_outValid_32 & _T_61612; // @[Switch.scala 41:38:@22772.4]
  assign _T_61615 = select_33 == 6'h8; // @[Switch.scala 41:52:@22774.4]
  assign output_8_33 = io_outValid_33 & _T_61615; // @[Switch.scala 41:38:@22775.4]
  assign _T_61618 = select_34 == 6'h8; // @[Switch.scala 41:52:@22777.4]
  assign output_8_34 = io_outValid_34 & _T_61618; // @[Switch.scala 41:38:@22778.4]
  assign _T_61621 = select_35 == 6'h8; // @[Switch.scala 41:52:@22780.4]
  assign output_8_35 = io_outValid_35 & _T_61621; // @[Switch.scala 41:38:@22781.4]
  assign _T_61624 = select_36 == 6'h8; // @[Switch.scala 41:52:@22783.4]
  assign output_8_36 = io_outValid_36 & _T_61624; // @[Switch.scala 41:38:@22784.4]
  assign _T_61627 = select_37 == 6'h8; // @[Switch.scala 41:52:@22786.4]
  assign output_8_37 = io_outValid_37 & _T_61627; // @[Switch.scala 41:38:@22787.4]
  assign _T_61630 = select_38 == 6'h8; // @[Switch.scala 41:52:@22789.4]
  assign output_8_38 = io_outValid_38 & _T_61630; // @[Switch.scala 41:38:@22790.4]
  assign _T_61633 = select_39 == 6'h8; // @[Switch.scala 41:52:@22792.4]
  assign output_8_39 = io_outValid_39 & _T_61633; // @[Switch.scala 41:38:@22793.4]
  assign _T_61636 = select_40 == 6'h8; // @[Switch.scala 41:52:@22795.4]
  assign output_8_40 = io_outValid_40 & _T_61636; // @[Switch.scala 41:38:@22796.4]
  assign _T_61639 = select_41 == 6'h8; // @[Switch.scala 41:52:@22798.4]
  assign output_8_41 = io_outValid_41 & _T_61639; // @[Switch.scala 41:38:@22799.4]
  assign _T_61642 = select_42 == 6'h8; // @[Switch.scala 41:52:@22801.4]
  assign output_8_42 = io_outValid_42 & _T_61642; // @[Switch.scala 41:38:@22802.4]
  assign _T_61645 = select_43 == 6'h8; // @[Switch.scala 41:52:@22804.4]
  assign output_8_43 = io_outValid_43 & _T_61645; // @[Switch.scala 41:38:@22805.4]
  assign _T_61648 = select_44 == 6'h8; // @[Switch.scala 41:52:@22807.4]
  assign output_8_44 = io_outValid_44 & _T_61648; // @[Switch.scala 41:38:@22808.4]
  assign _T_61651 = select_45 == 6'h8; // @[Switch.scala 41:52:@22810.4]
  assign output_8_45 = io_outValid_45 & _T_61651; // @[Switch.scala 41:38:@22811.4]
  assign _T_61654 = select_46 == 6'h8; // @[Switch.scala 41:52:@22813.4]
  assign output_8_46 = io_outValid_46 & _T_61654; // @[Switch.scala 41:38:@22814.4]
  assign _T_61657 = select_47 == 6'h8; // @[Switch.scala 41:52:@22816.4]
  assign output_8_47 = io_outValid_47 & _T_61657; // @[Switch.scala 41:38:@22817.4]
  assign _T_61660 = select_48 == 6'h8; // @[Switch.scala 41:52:@22819.4]
  assign output_8_48 = io_outValid_48 & _T_61660; // @[Switch.scala 41:38:@22820.4]
  assign _T_61663 = select_49 == 6'h8; // @[Switch.scala 41:52:@22822.4]
  assign output_8_49 = io_outValid_49 & _T_61663; // @[Switch.scala 41:38:@22823.4]
  assign _T_61666 = select_50 == 6'h8; // @[Switch.scala 41:52:@22825.4]
  assign output_8_50 = io_outValid_50 & _T_61666; // @[Switch.scala 41:38:@22826.4]
  assign _T_61669 = select_51 == 6'h8; // @[Switch.scala 41:52:@22828.4]
  assign output_8_51 = io_outValid_51 & _T_61669; // @[Switch.scala 41:38:@22829.4]
  assign _T_61672 = select_52 == 6'h8; // @[Switch.scala 41:52:@22831.4]
  assign output_8_52 = io_outValid_52 & _T_61672; // @[Switch.scala 41:38:@22832.4]
  assign _T_61675 = select_53 == 6'h8; // @[Switch.scala 41:52:@22834.4]
  assign output_8_53 = io_outValid_53 & _T_61675; // @[Switch.scala 41:38:@22835.4]
  assign _T_61678 = select_54 == 6'h8; // @[Switch.scala 41:52:@22837.4]
  assign output_8_54 = io_outValid_54 & _T_61678; // @[Switch.scala 41:38:@22838.4]
  assign _T_61681 = select_55 == 6'h8; // @[Switch.scala 41:52:@22840.4]
  assign output_8_55 = io_outValid_55 & _T_61681; // @[Switch.scala 41:38:@22841.4]
  assign _T_61684 = select_56 == 6'h8; // @[Switch.scala 41:52:@22843.4]
  assign output_8_56 = io_outValid_56 & _T_61684; // @[Switch.scala 41:38:@22844.4]
  assign _T_61687 = select_57 == 6'h8; // @[Switch.scala 41:52:@22846.4]
  assign output_8_57 = io_outValid_57 & _T_61687; // @[Switch.scala 41:38:@22847.4]
  assign _T_61690 = select_58 == 6'h8; // @[Switch.scala 41:52:@22849.4]
  assign output_8_58 = io_outValid_58 & _T_61690; // @[Switch.scala 41:38:@22850.4]
  assign _T_61693 = select_59 == 6'h8; // @[Switch.scala 41:52:@22852.4]
  assign output_8_59 = io_outValid_59 & _T_61693; // @[Switch.scala 41:38:@22853.4]
  assign _T_61696 = select_60 == 6'h8; // @[Switch.scala 41:52:@22855.4]
  assign output_8_60 = io_outValid_60 & _T_61696; // @[Switch.scala 41:38:@22856.4]
  assign _T_61699 = select_61 == 6'h8; // @[Switch.scala 41:52:@22858.4]
  assign output_8_61 = io_outValid_61 & _T_61699; // @[Switch.scala 41:38:@22859.4]
  assign _T_61702 = select_62 == 6'h8; // @[Switch.scala 41:52:@22861.4]
  assign output_8_62 = io_outValid_62 & _T_61702; // @[Switch.scala 41:38:@22862.4]
  assign _T_61705 = select_63 == 6'h8; // @[Switch.scala 41:52:@22864.4]
  assign output_8_63 = io_outValid_63 & _T_61705; // @[Switch.scala 41:38:@22865.4]
  assign _T_61713 = {output_8_7,output_8_6,output_8_5,output_8_4,output_8_3,output_8_2,output_8_1,output_8_0}; // @[Switch.scala 43:31:@22873.4]
  assign _T_61721 = {output_8_15,output_8_14,output_8_13,output_8_12,output_8_11,output_8_10,output_8_9,output_8_8,_T_61713}; // @[Switch.scala 43:31:@22881.4]
  assign _T_61728 = {output_8_23,output_8_22,output_8_21,output_8_20,output_8_19,output_8_18,output_8_17,output_8_16}; // @[Switch.scala 43:31:@22888.4]
  assign _T_61737 = {output_8_31,output_8_30,output_8_29,output_8_28,output_8_27,output_8_26,output_8_25,output_8_24,_T_61728,_T_61721}; // @[Switch.scala 43:31:@22897.4]
  assign _T_61744 = {output_8_39,output_8_38,output_8_37,output_8_36,output_8_35,output_8_34,output_8_33,output_8_32}; // @[Switch.scala 43:31:@22904.4]
  assign _T_61752 = {output_8_47,output_8_46,output_8_45,output_8_44,output_8_43,output_8_42,output_8_41,output_8_40,_T_61744}; // @[Switch.scala 43:31:@22912.4]
  assign _T_61759 = {output_8_55,output_8_54,output_8_53,output_8_52,output_8_51,output_8_50,output_8_49,output_8_48}; // @[Switch.scala 43:31:@22919.4]
  assign _T_61768 = {output_8_63,output_8_62,output_8_61,output_8_60,output_8_59,output_8_58,output_8_57,output_8_56,_T_61759,_T_61752}; // @[Switch.scala 43:31:@22928.4]
  assign _T_61769 = {_T_61768,_T_61737}; // @[Switch.scala 43:31:@22929.4]
  assign _T_61773 = select_0 == 6'h9; // @[Switch.scala 41:52:@22932.4]
  assign output_9_0 = io_outValid_0 & _T_61773; // @[Switch.scala 41:38:@22933.4]
  assign _T_61776 = select_1 == 6'h9; // @[Switch.scala 41:52:@22935.4]
  assign output_9_1 = io_outValid_1 & _T_61776; // @[Switch.scala 41:38:@22936.4]
  assign _T_61779 = select_2 == 6'h9; // @[Switch.scala 41:52:@22938.4]
  assign output_9_2 = io_outValid_2 & _T_61779; // @[Switch.scala 41:38:@22939.4]
  assign _T_61782 = select_3 == 6'h9; // @[Switch.scala 41:52:@22941.4]
  assign output_9_3 = io_outValid_3 & _T_61782; // @[Switch.scala 41:38:@22942.4]
  assign _T_61785 = select_4 == 6'h9; // @[Switch.scala 41:52:@22944.4]
  assign output_9_4 = io_outValid_4 & _T_61785; // @[Switch.scala 41:38:@22945.4]
  assign _T_61788 = select_5 == 6'h9; // @[Switch.scala 41:52:@22947.4]
  assign output_9_5 = io_outValid_5 & _T_61788; // @[Switch.scala 41:38:@22948.4]
  assign _T_61791 = select_6 == 6'h9; // @[Switch.scala 41:52:@22950.4]
  assign output_9_6 = io_outValid_6 & _T_61791; // @[Switch.scala 41:38:@22951.4]
  assign _T_61794 = select_7 == 6'h9; // @[Switch.scala 41:52:@22953.4]
  assign output_9_7 = io_outValid_7 & _T_61794; // @[Switch.scala 41:38:@22954.4]
  assign _T_61797 = select_8 == 6'h9; // @[Switch.scala 41:52:@22956.4]
  assign output_9_8 = io_outValid_8 & _T_61797; // @[Switch.scala 41:38:@22957.4]
  assign _T_61800 = select_9 == 6'h9; // @[Switch.scala 41:52:@22959.4]
  assign output_9_9 = io_outValid_9 & _T_61800; // @[Switch.scala 41:38:@22960.4]
  assign _T_61803 = select_10 == 6'h9; // @[Switch.scala 41:52:@22962.4]
  assign output_9_10 = io_outValid_10 & _T_61803; // @[Switch.scala 41:38:@22963.4]
  assign _T_61806 = select_11 == 6'h9; // @[Switch.scala 41:52:@22965.4]
  assign output_9_11 = io_outValid_11 & _T_61806; // @[Switch.scala 41:38:@22966.4]
  assign _T_61809 = select_12 == 6'h9; // @[Switch.scala 41:52:@22968.4]
  assign output_9_12 = io_outValid_12 & _T_61809; // @[Switch.scala 41:38:@22969.4]
  assign _T_61812 = select_13 == 6'h9; // @[Switch.scala 41:52:@22971.4]
  assign output_9_13 = io_outValid_13 & _T_61812; // @[Switch.scala 41:38:@22972.4]
  assign _T_61815 = select_14 == 6'h9; // @[Switch.scala 41:52:@22974.4]
  assign output_9_14 = io_outValid_14 & _T_61815; // @[Switch.scala 41:38:@22975.4]
  assign _T_61818 = select_15 == 6'h9; // @[Switch.scala 41:52:@22977.4]
  assign output_9_15 = io_outValid_15 & _T_61818; // @[Switch.scala 41:38:@22978.4]
  assign _T_61821 = select_16 == 6'h9; // @[Switch.scala 41:52:@22980.4]
  assign output_9_16 = io_outValid_16 & _T_61821; // @[Switch.scala 41:38:@22981.4]
  assign _T_61824 = select_17 == 6'h9; // @[Switch.scala 41:52:@22983.4]
  assign output_9_17 = io_outValid_17 & _T_61824; // @[Switch.scala 41:38:@22984.4]
  assign _T_61827 = select_18 == 6'h9; // @[Switch.scala 41:52:@22986.4]
  assign output_9_18 = io_outValid_18 & _T_61827; // @[Switch.scala 41:38:@22987.4]
  assign _T_61830 = select_19 == 6'h9; // @[Switch.scala 41:52:@22989.4]
  assign output_9_19 = io_outValid_19 & _T_61830; // @[Switch.scala 41:38:@22990.4]
  assign _T_61833 = select_20 == 6'h9; // @[Switch.scala 41:52:@22992.4]
  assign output_9_20 = io_outValid_20 & _T_61833; // @[Switch.scala 41:38:@22993.4]
  assign _T_61836 = select_21 == 6'h9; // @[Switch.scala 41:52:@22995.4]
  assign output_9_21 = io_outValid_21 & _T_61836; // @[Switch.scala 41:38:@22996.4]
  assign _T_61839 = select_22 == 6'h9; // @[Switch.scala 41:52:@22998.4]
  assign output_9_22 = io_outValid_22 & _T_61839; // @[Switch.scala 41:38:@22999.4]
  assign _T_61842 = select_23 == 6'h9; // @[Switch.scala 41:52:@23001.4]
  assign output_9_23 = io_outValid_23 & _T_61842; // @[Switch.scala 41:38:@23002.4]
  assign _T_61845 = select_24 == 6'h9; // @[Switch.scala 41:52:@23004.4]
  assign output_9_24 = io_outValid_24 & _T_61845; // @[Switch.scala 41:38:@23005.4]
  assign _T_61848 = select_25 == 6'h9; // @[Switch.scala 41:52:@23007.4]
  assign output_9_25 = io_outValid_25 & _T_61848; // @[Switch.scala 41:38:@23008.4]
  assign _T_61851 = select_26 == 6'h9; // @[Switch.scala 41:52:@23010.4]
  assign output_9_26 = io_outValid_26 & _T_61851; // @[Switch.scala 41:38:@23011.4]
  assign _T_61854 = select_27 == 6'h9; // @[Switch.scala 41:52:@23013.4]
  assign output_9_27 = io_outValid_27 & _T_61854; // @[Switch.scala 41:38:@23014.4]
  assign _T_61857 = select_28 == 6'h9; // @[Switch.scala 41:52:@23016.4]
  assign output_9_28 = io_outValid_28 & _T_61857; // @[Switch.scala 41:38:@23017.4]
  assign _T_61860 = select_29 == 6'h9; // @[Switch.scala 41:52:@23019.4]
  assign output_9_29 = io_outValid_29 & _T_61860; // @[Switch.scala 41:38:@23020.4]
  assign _T_61863 = select_30 == 6'h9; // @[Switch.scala 41:52:@23022.4]
  assign output_9_30 = io_outValid_30 & _T_61863; // @[Switch.scala 41:38:@23023.4]
  assign _T_61866 = select_31 == 6'h9; // @[Switch.scala 41:52:@23025.4]
  assign output_9_31 = io_outValid_31 & _T_61866; // @[Switch.scala 41:38:@23026.4]
  assign _T_61869 = select_32 == 6'h9; // @[Switch.scala 41:52:@23028.4]
  assign output_9_32 = io_outValid_32 & _T_61869; // @[Switch.scala 41:38:@23029.4]
  assign _T_61872 = select_33 == 6'h9; // @[Switch.scala 41:52:@23031.4]
  assign output_9_33 = io_outValid_33 & _T_61872; // @[Switch.scala 41:38:@23032.4]
  assign _T_61875 = select_34 == 6'h9; // @[Switch.scala 41:52:@23034.4]
  assign output_9_34 = io_outValid_34 & _T_61875; // @[Switch.scala 41:38:@23035.4]
  assign _T_61878 = select_35 == 6'h9; // @[Switch.scala 41:52:@23037.4]
  assign output_9_35 = io_outValid_35 & _T_61878; // @[Switch.scala 41:38:@23038.4]
  assign _T_61881 = select_36 == 6'h9; // @[Switch.scala 41:52:@23040.4]
  assign output_9_36 = io_outValid_36 & _T_61881; // @[Switch.scala 41:38:@23041.4]
  assign _T_61884 = select_37 == 6'h9; // @[Switch.scala 41:52:@23043.4]
  assign output_9_37 = io_outValid_37 & _T_61884; // @[Switch.scala 41:38:@23044.4]
  assign _T_61887 = select_38 == 6'h9; // @[Switch.scala 41:52:@23046.4]
  assign output_9_38 = io_outValid_38 & _T_61887; // @[Switch.scala 41:38:@23047.4]
  assign _T_61890 = select_39 == 6'h9; // @[Switch.scala 41:52:@23049.4]
  assign output_9_39 = io_outValid_39 & _T_61890; // @[Switch.scala 41:38:@23050.4]
  assign _T_61893 = select_40 == 6'h9; // @[Switch.scala 41:52:@23052.4]
  assign output_9_40 = io_outValid_40 & _T_61893; // @[Switch.scala 41:38:@23053.4]
  assign _T_61896 = select_41 == 6'h9; // @[Switch.scala 41:52:@23055.4]
  assign output_9_41 = io_outValid_41 & _T_61896; // @[Switch.scala 41:38:@23056.4]
  assign _T_61899 = select_42 == 6'h9; // @[Switch.scala 41:52:@23058.4]
  assign output_9_42 = io_outValid_42 & _T_61899; // @[Switch.scala 41:38:@23059.4]
  assign _T_61902 = select_43 == 6'h9; // @[Switch.scala 41:52:@23061.4]
  assign output_9_43 = io_outValid_43 & _T_61902; // @[Switch.scala 41:38:@23062.4]
  assign _T_61905 = select_44 == 6'h9; // @[Switch.scala 41:52:@23064.4]
  assign output_9_44 = io_outValid_44 & _T_61905; // @[Switch.scala 41:38:@23065.4]
  assign _T_61908 = select_45 == 6'h9; // @[Switch.scala 41:52:@23067.4]
  assign output_9_45 = io_outValid_45 & _T_61908; // @[Switch.scala 41:38:@23068.4]
  assign _T_61911 = select_46 == 6'h9; // @[Switch.scala 41:52:@23070.4]
  assign output_9_46 = io_outValid_46 & _T_61911; // @[Switch.scala 41:38:@23071.4]
  assign _T_61914 = select_47 == 6'h9; // @[Switch.scala 41:52:@23073.4]
  assign output_9_47 = io_outValid_47 & _T_61914; // @[Switch.scala 41:38:@23074.4]
  assign _T_61917 = select_48 == 6'h9; // @[Switch.scala 41:52:@23076.4]
  assign output_9_48 = io_outValid_48 & _T_61917; // @[Switch.scala 41:38:@23077.4]
  assign _T_61920 = select_49 == 6'h9; // @[Switch.scala 41:52:@23079.4]
  assign output_9_49 = io_outValid_49 & _T_61920; // @[Switch.scala 41:38:@23080.4]
  assign _T_61923 = select_50 == 6'h9; // @[Switch.scala 41:52:@23082.4]
  assign output_9_50 = io_outValid_50 & _T_61923; // @[Switch.scala 41:38:@23083.4]
  assign _T_61926 = select_51 == 6'h9; // @[Switch.scala 41:52:@23085.4]
  assign output_9_51 = io_outValid_51 & _T_61926; // @[Switch.scala 41:38:@23086.4]
  assign _T_61929 = select_52 == 6'h9; // @[Switch.scala 41:52:@23088.4]
  assign output_9_52 = io_outValid_52 & _T_61929; // @[Switch.scala 41:38:@23089.4]
  assign _T_61932 = select_53 == 6'h9; // @[Switch.scala 41:52:@23091.4]
  assign output_9_53 = io_outValid_53 & _T_61932; // @[Switch.scala 41:38:@23092.4]
  assign _T_61935 = select_54 == 6'h9; // @[Switch.scala 41:52:@23094.4]
  assign output_9_54 = io_outValid_54 & _T_61935; // @[Switch.scala 41:38:@23095.4]
  assign _T_61938 = select_55 == 6'h9; // @[Switch.scala 41:52:@23097.4]
  assign output_9_55 = io_outValid_55 & _T_61938; // @[Switch.scala 41:38:@23098.4]
  assign _T_61941 = select_56 == 6'h9; // @[Switch.scala 41:52:@23100.4]
  assign output_9_56 = io_outValid_56 & _T_61941; // @[Switch.scala 41:38:@23101.4]
  assign _T_61944 = select_57 == 6'h9; // @[Switch.scala 41:52:@23103.4]
  assign output_9_57 = io_outValid_57 & _T_61944; // @[Switch.scala 41:38:@23104.4]
  assign _T_61947 = select_58 == 6'h9; // @[Switch.scala 41:52:@23106.4]
  assign output_9_58 = io_outValid_58 & _T_61947; // @[Switch.scala 41:38:@23107.4]
  assign _T_61950 = select_59 == 6'h9; // @[Switch.scala 41:52:@23109.4]
  assign output_9_59 = io_outValid_59 & _T_61950; // @[Switch.scala 41:38:@23110.4]
  assign _T_61953 = select_60 == 6'h9; // @[Switch.scala 41:52:@23112.4]
  assign output_9_60 = io_outValid_60 & _T_61953; // @[Switch.scala 41:38:@23113.4]
  assign _T_61956 = select_61 == 6'h9; // @[Switch.scala 41:52:@23115.4]
  assign output_9_61 = io_outValid_61 & _T_61956; // @[Switch.scala 41:38:@23116.4]
  assign _T_61959 = select_62 == 6'h9; // @[Switch.scala 41:52:@23118.4]
  assign output_9_62 = io_outValid_62 & _T_61959; // @[Switch.scala 41:38:@23119.4]
  assign _T_61962 = select_63 == 6'h9; // @[Switch.scala 41:52:@23121.4]
  assign output_9_63 = io_outValid_63 & _T_61962; // @[Switch.scala 41:38:@23122.4]
  assign _T_61970 = {output_9_7,output_9_6,output_9_5,output_9_4,output_9_3,output_9_2,output_9_1,output_9_0}; // @[Switch.scala 43:31:@23130.4]
  assign _T_61978 = {output_9_15,output_9_14,output_9_13,output_9_12,output_9_11,output_9_10,output_9_9,output_9_8,_T_61970}; // @[Switch.scala 43:31:@23138.4]
  assign _T_61985 = {output_9_23,output_9_22,output_9_21,output_9_20,output_9_19,output_9_18,output_9_17,output_9_16}; // @[Switch.scala 43:31:@23145.4]
  assign _T_61994 = {output_9_31,output_9_30,output_9_29,output_9_28,output_9_27,output_9_26,output_9_25,output_9_24,_T_61985,_T_61978}; // @[Switch.scala 43:31:@23154.4]
  assign _T_62001 = {output_9_39,output_9_38,output_9_37,output_9_36,output_9_35,output_9_34,output_9_33,output_9_32}; // @[Switch.scala 43:31:@23161.4]
  assign _T_62009 = {output_9_47,output_9_46,output_9_45,output_9_44,output_9_43,output_9_42,output_9_41,output_9_40,_T_62001}; // @[Switch.scala 43:31:@23169.4]
  assign _T_62016 = {output_9_55,output_9_54,output_9_53,output_9_52,output_9_51,output_9_50,output_9_49,output_9_48}; // @[Switch.scala 43:31:@23176.4]
  assign _T_62025 = {output_9_63,output_9_62,output_9_61,output_9_60,output_9_59,output_9_58,output_9_57,output_9_56,_T_62016,_T_62009}; // @[Switch.scala 43:31:@23185.4]
  assign _T_62026 = {_T_62025,_T_61994}; // @[Switch.scala 43:31:@23186.4]
  assign _T_62030 = select_0 == 6'ha; // @[Switch.scala 41:52:@23189.4]
  assign output_10_0 = io_outValid_0 & _T_62030; // @[Switch.scala 41:38:@23190.4]
  assign _T_62033 = select_1 == 6'ha; // @[Switch.scala 41:52:@23192.4]
  assign output_10_1 = io_outValid_1 & _T_62033; // @[Switch.scala 41:38:@23193.4]
  assign _T_62036 = select_2 == 6'ha; // @[Switch.scala 41:52:@23195.4]
  assign output_10_2 = io_outValid_2 & _T_62036; // @[Switch.scala 41:38:@23196.4]
  assign _T_62039 = select_3 == 6'ha; // @[Switch.scala 41:52:@23198.4]
  assign output_10_3 = io_outValid_3 & _T_62039; // @[Switch.scala 41:38:@23199.4]
  assign _T_62042 = select_4 == 6'ha; // @[Switch.scala 41:52:@23201.4]
  assign output_10_4 = io_outValid_4 & _T_62042; // @[Switch.scala 41:38:@23202.4]
  assign _T_62045 = select_5 == 6'ha; // @[Switch.scala 41:52:@23204.4]
  assign output_10_5 = io_outValid_5 & _T_62045; // @[Switch.scala 41:38:@23205.4]
  assign _T_62048 = select_6 == 6'ha; // @[Switch.scala 41:52:@23207.4]
  assign output_10_6 = io_outValid_6 & _T_62048; // @[Switch.scala 41:38:@23208.4]
  assign _T_62051 = select_7 == 6'ha; // @[Switch.scala 41:52:@23210.4]
  assign output_10_7 = io_outValid_7 & _T_62051; // @[Switch.scala 41:38:@23211.4]
  assign _T_62054 = select_8 == 6'ha; // @[Switch.scala 41:52:@23213.4]
  assign output_10_8 = io_outValid_8 & _T_62054; // @[Switch.scala 41:38:@23214.4]
  assign _T_62057 = select_9 == 6'ha; // @[Switch.scala 41:52:@23216.4]
  assign output_10_9 = io_outValid_9 & _T_62057; // @[Switch.scala 41:38:@23217.4]
  assign _T_62060 = select_10 == 6'ha; // @[Switch.scala 41:52:@23219.4]
  assign output_10_10 = io_outValid_10 & _T_62060; // @[Switch.scala 41:38:@23220.4]
  assign _T_62063 = select_11 == 6'ha; // @[Switch.scala 41:52:@23222.4]
  assign output_10_11 = io_outValid_11 & _T_62063; // @[Switch.scala 41:38:@23223.4]
  assign _T_62066 = select_12 == 6'ha; // @[Switch.scala 41:52:@23225.4]
  assign output_10_12 = io_outValid_12 & _T_62066; // @[Switch.scala 41:38:@23226.4]
  assign _T_62069 = select_13 == 6'ha; // @[Switch.scala 41:52:@23228.4]
  assign output_10_13 = io_outValid_13 & _T_62069; // @[Switch.scala 41:38:@23229.4]
  assign _T_62072 = select_14 == 6'ha; // @[Switch.scala 41:52:@23231.4]
  assign output_10_14 = io_outValid_14 & _T_62072; // @[Switch.scala 41:38:@23232.4]
  assign _T_62075 = select_15 == 6'ha; // @[Switch.scala 41:52:@23234.4]
  assign output_10_15 = io_outValid_15 & _T_62075; // @[Switch.scala 41:38:@23235.4]
  assign _T_62078 = select_16 == 6'ha; // @[Switch.scala 41:52:@23237.4]
  assign output_10_16 = io_outValid_16 & _T_62078; // @[Switch.scala 41:38:@23238.4]
  assign _T_62081 = select_17 == 6'ha; // @[Switch.scala 41:52:@23240.4]
  assign output_10_17 = io_outValid_17 & _T_62081; // @[Switch.scala 41:38:@23241.4]
  assign _T_62084 = select_18 == 6'ha; // @[Switch.scala 41:52:@23243.4]
  assign output_10_18 = io_outValid_18 & _T_62084; // @[Switch.scala 41:38:@23244.4]
  assign _T_62087 = select_19 == 6'ha; // @[Switch.scala 41:52:@23246.4]
  assign output_10_19 = io_outValid_19 & _T_62087; // @[Switch.scala 41:38:@23247.4]
  assign _T_62090 = select_20 == 6'ha; // @[Switch.scala 41:52:@23249.4]
  assign output_10_20 = io_outValid_20 & _T_62090; // @[Switch.scala 41:38:@23250.4]
  assign _T_62093 = select_21 == 6'ha; // @[Switch.scala 41:52:@23252.4]
  assign output_10_21 = io_outValid_21 & _T_62093; // @[Switch.scala 41:38:@23253.4]
  assign _T_62096 = select_22 == 6'ha; // @[Switch.scala 41:52:@23255.4]
  assign output_10_22 = io_outValid_22 & _T_62096; // @[Switch.scala 41:38:@23256.4]
  assign _T_62099 = select_23 == 6'ha; // @[Switch.scala 41:52:@23258.4]
  assign output_10_23 = io_outValid_23 & _T_62099; // @[Switch.scala 41:38:@23259.4]
  assign _T_62102 = select_24 == 6'ha; // @[Switch.scala 41:52:@23261.4]
  assign output_10_24 = io_outValid_24 & _T_62102; // @[Switch.scala 41:38:@23262.4]
  assign _T_62105 = select_25 == 6'ha; // @[Switch.scala 41:52:@23264.4]
  assign output_10_25 = io_outValid_25 & _T_62105; // @[Switch.scala 41:38:@23265.4]
  assign _T_62108 = select_26 == 6'ha; // @[Switch.scala 41:52:@23267.4]
  assign output_10_26 = io_outValid_26 & _T_62108; // @[Switch.scala 41:38:@23268.4]
  assign _T_62111 = select_27 == 6'ha; // @[Switch.scala 41:52:@23270.4]
  assign output_10_27 = io_outValid_27 & _T_62111; // @[Switch.scala 41:38:@23271.4]
  assign _T_62114 = select_28 == 6'ha; // @[Switch.scala 41:52:@23273.4]
  assign output_10_28 = io_outValid_28 & _T_62114; // @[Switch.scala 41:38:@23274.4]
  assign _T_62117 = select_29 == 6'ha; // @[Switch.scala 41:52:@23276.4]
  assign output_10_29 = io_outValid_29 & _T_62117; // @[Switch.scala 41:38:@23277.4]
  assign _T_62120 = select_30 == 6'ha; // @[Switch.scala 41:52:@23279.4]
  assign output_10_30 = io_outValid_30 & _T_62120; // @[Switch.scala 41:38:@23280.4]
  assign _T_62123 = select_31 == 6'ha; // @[Switch.scala 41:52:@23282.4]
  assign output_10_31 = io_outValid_31 & _T_62123; // @[Switch.scala 41:38:@23283.4]
  assign _T_62126 = select_32 == 6'ha; // @[Switch.scala 41:52:@23285.4]
  assign output_10_32 = io_outValid_32 & _T_62126; // @[Switch.scala 41:38:@23286.4]
  assign _T_62129 = select_33 == 6'ha; // @[Switch.scala 41:52:@23288.4]
  assign output_10_33 = io_outValid_33 & _T_62129; // @[Switch.scala 41:38:@23289.4]
  assign _T_62132 = select_34 == 6'ha; // @[Switch.scala 41:52:@23291.4]
  assign output_10_34 = io_outValid_34 & _T_62132; // @[Switch.scala 41:38:@23292.4]
  assign _T_62135 = select_35 == 6'ha; // @[Switch.scala 41:52:@23294.4]
  assign output_10_35 = io_outValid_35 & _T_62135; // @[Switch.scala 41:38:@23295.4]
  assign _T_62138 = select_36 == 6'ha; // @[Switch.scala 41:52:@23297.4]
  assign output_10_36 = io_outValid_36 & _T_62138; // @[Switch.scala 41:38:@23298.4]
  assign _T_62141 = select_37 == 6'ha; // @[Switch.scala 41:52:@23300.4]
  assign output_10_37 = io_outValid_37 & _T_62141; // @[Switch.scala 41:38:@23301.4]
  assign _T_62144 = select_38 == 6'ha; // @[Switch.scala 41:52:@23303.4]
  assign output_10_38 = io_outValid_38 & _T_62144; // @[Switch.scala 41:38:@23304.4]
  assign _T_62147 = select_39 == 6'ha; // @[Switch.scala 41:52:@23306.4]
  assign output_10_39 = io_outValid_39 & _T_62147; // @[Switch.scala 41:38:@23307.4]
  assign _T_62150 = select_40 == 6'ha; // @[Switch.scala 41:52:@23309.4]
  assign output_10_40 = io_outValid_40 & _T_62150; // @[Switch.scala 41:38:@23310.4]
  assign _T_62153 = select_41 == 6'ha; // @[Switch.scala 41:52:@23312.4]
  assign output_10_41 = io_outValid_41 & _T_62153; // @[Switch.scala 41:38:@23313.4]
  assign _T_62156 = select_42 == 6'ha; // @[Switch.scala 41:52:@23315.4]
  assign output_10_42 = io_outValid_42 & _T_62156; // @[Switch.scala 41:38:@23316.4]
  assign _T_62159 = select_43 == 6'ha; // @[Switch.scala 41:52:@23318.4]
  assign output_10_43 = io_outValid_43 & _T_62159; // @[Switch.scala 41:38:@23319.4]
  assign _T_62162 = select_44 == 6'ha; // @[Switch.scala 41:52:@23321.4]
  assign output_10_44 = io_outValid_44 & _T_62162; // @[Switch.scala 41:38:@23322.4]
  assign _T_62165 = select_45 == 6'ha; // @[Switch.scala 41:52:@23324.4]
  assign output_10_45 = io_outValid_45 & _T_62165; // @[Switch.scala 41:38:@23325.4]
  assign _T_62168 = select_46 == 6'ha; // @[Switch.scala 41:52:@23327.4]
  assign output_10_46 = io_outValid_46 & _T_62168; // @[Switch.scala 41:38:@23328.4]
  assign _T_62171 = select_47 == 6'ha; // @[Switch.scala 41:52:@23330.4]
  assign output_10_47 = io_outValid_47 & _T_62171; // @[Switch.scala 41:38:@23331.4]
  assign _T_62174 = select_48 == 6'ha; // @[Switch.scala 41:52:@23333.4]
  assign output_10_48 = io_outValid_48 & _T_62174; // @[Switch.scala 41:38:@23334.4]
  assign _T_62177 = select_49 == 6'ha; // @[Switch.scala 41:52:@23336.4]
  assign output_10_49 = io_outValid_49 & _T_62177; // @[Switch.scala 41:38:@23337.4]
  assign _T_62180 = select_50 == 6'ha; // @[Switch.scala 41:52:@23339.4]
  assign output_10_50 = io_outValid_50 & _T_62180; // @[Switch.scala 41:38:@23340.4]
  assign _T_62183 = select_51 == 6'ha; // @[Switch.scala 41:52:@23342.4]
  assign output_10_51 = io_outValid_51 & _T_62183; // @[Switch.scala 41:38:@23343.4]
  assign _T_62186 = select_52 == 6'ha; // @[Switch.scala 41:52:@23345.4]
  assign output_10_52 = io_outValid_52 & _T_62186; // @[Switch.scala 41:38:@23346.4]
  assign _T_62189 = select_53 == 6'ha; // @[Switch.scala 41:52:@23348.4]
  assign output_10_53 = io_outValid_53 & _T_62189; // @[Switch.scala 41:38:@23349.4]
  assign _T_62192 = select_54 == 6'ha; // @[Switch.scala 41:52:@23351.4]
  assign output_10_54 = io_outValid_54 & _T_62192; // @[Switch.scala 41:38:@23352.4]
  assign _T_62195 = select_55 == 6'ha; // @[Switch.scala 41:52:@23354.4]
  assign output_10_55 = io_outValid_55 & _T_62195; // @[Switch.scala 41:38:@23355.4]
  assign _T_62198 = select_56 == 6'ha; // @[Switch.scala 41:52:@23357.4]
  assign output_10_56 = io_outValid_56 & _T_62198; // @[Switch.scala 41:38:@23358.4]
  assign _T_62201 = select_57 == 6'ha; // @[Switch.scala 41:52:@23360.4]
  assign output_10_57 = io_outValid_57 & _T_62201; // @[Switch.scala 41:38:@23361.4]
  assign _T_62204 = select_58 == 6'ha; // @[Switch.scala 41:52:@23363.4]
  assign output_10_58 = io_outValid_58 & _T_62204; // @[Switch.scala 41:38:@23364.4]
  assign _T_62207 = select_59 == 6'ha; // @[Switch.scala 41:52:@23366.4]
  assign output_10_59 = io_outValid_59 & _T_62207; // @[Switch.scala 41:38:@23367.4]
  assign _T_62210 = select_60 == 6'ha; // @[Switch.scala 41:52:@23369.4]
  assign output_10_60 = io_outValid_60 & _T_62210; // @[Switch.scala 41:38:@23370.4]
  assign _T_62213 = select_61 == 6'ha; // @[Switch.scala 41:52:@23372.4]
  assign output_10_61 = io_outValid_61 & _T_62213; // @[Switch.scala 41:38:@23373.4]
  assign _T_62216 = select_62 == 6'ha; // @[Switch.scala 41:52:@23375.4]
  assign output_10_62 = io_outValid_62 & _T_62216; // @[Switch.scala 41:38:@23376.4]
  assign _T_62219 = select_63 == 6'ha; // @[Switch.scala 41:52:@23378.4]
  assign output_10_63 = io_outValid_63 & _T_62219; // @[Switch.scala 41:38:@23379.4]
  assign _T_62227 = {output_10_7,output_10_6,output_10_5,output_10_4,output_10_3,output_10_2,output_10_1,output_10_0}; // @[Switch.scala 43:31:@23387.4]
  assign _T_62235 = {output_10_15,output_10_14,output_10_13,output_10_12,output_10_11,output_10_10,output_10_9,output_10_8,_T_62227}; // @[Switch.scala 43:31:@23395.4]
  assign _T_62242 = {output_10_23,output_10_22,output_10_21,output_10_20,output_10_19,output_10_18,output_10_17,output_10_16}; // @[Switch.scala 43:31:@23402.4]
  assign _T_62251 = {output_10_31,output_10_30,output_10_29,output_10_28,output_10_27,output_10_26,output_10_25,output_10_24,_T_62242,_T_62235}; // @[Switch.scala 43:31:@23411.4]
  assign _T_62258 = {output_10_39,output_10_38,output_10_37,output_10_36,output_10_35,output_10_34,output_10_33,output_10_32}; // @[Switch.scala 43:31:@23418.4]
  assign _T_62266 = {output_10_47,output_10_46,output_10_45,output_10_44,output_10_43,output_10_42,output_10_41,output_10_40,_T_62258}; // @[Switch.scala 43:31:@23426.4]
  assign _T_62273 = {output_10_55,output_10_54,output_10_53,output_10_52,output_10_51,output_10_50,output_10_49,output_10_48}; // @[Switch.scala 43:31:@23433.4]
  assign _T_62282 = {output_10_63,output_10_62,output_10_61,output_10_60,output_10_59,output_10_58,output_10_57,output_10_56,_T_62273,_T_62266}; // @[Switch.scala 43:31:@23442.4]
  assign _T_62283 = {_T_62282,_T_62251}; // @[Switch.scala 43:31:@23443.4]
  assign _T_62287 = select_0 == 6'hb; // @[Switch.scala 41:52:@23446.4]
  assign output_11_0 = io_outValid_0 & _T_62287; // @[Switch.scala 41:38:@23447.4]
  assign _T_62290 = select_1 == 6'hb; // @[Switch.scala 41:52:@23449.4]
  assign output_11_1 = io_outValid_1 & _T_62290; // @[Switch.scala 41:38:@23450.4]
  assign _T_62293 = select_2 == 6'hb; // @[Switch.scala 41:52:@23452.4]
  assign output_11_2 = io_outValid_2 & _T_62293; // @[Switch.scala 41:38:@23453.4]
  assign _T_62296 = select_3 == 6'hb; // @[Switch.scala 41:52:@23455.4]
  assign output_11_3 = io_outValid_3 & _T_62296; // @[Switch.scala 41:38:@23456.4]
  assign _T_62299 = select_4 == 6'hb; // @[Switch.scala 41:52:@23458.4]
  assign output_11_4 = io_outValid_4 & _T_62299; // @[Switch.scala 41:38:@23459.4]
  assign _T_62302 = select_5 == 6'hb; // @[Switch.scala 41:52:@23461.4]
  assign output_11_5 = io_outValid_5 & _T_62302; // @[Switch.scala 41:38:@23462.4]
  assign _T_62305 = select_6 == 6'hb; // @[Switch.scala 41:52:@23464.4]
  assign output_11_6 = io_outValid_6 & _T_62305; // @[Switch.scala 41:38:@23465.4]
  assign _T_62308 = select_7 == 6'hb; // @[Switch.scala 41:52:@23467.4]
  assign output_11_7 = io_outValid_7 & _T_62308; // @[Switch.scala 41:38:@23468.4]
  assign _T_62311 = select_8 == 6'hb; // @[Switch.scala 41:52:@23470.4]
  assign output_11_8 = io_outValid_8 & _T_62311; // @[Switch.scala 41:38:@23471.4]
  assign _T_62314 = select_9 == 6'hb; // @[Switch.scala 41:52:@23473.4]
  assign output_11_9 = io_outValid_9 & _T_62314; // @[Switch.scala 41:38:@23474.4]
  assign _T_62317 = select_10 == 6'hb; // @[Switch.scala 41:52:@23476.4]
  assign output_11_10 = io_outValid_10 & _T_62317; // @[Switch.scala 41:38:@23477.4]
  assign _T_62320 = select_11 == 6'hb; // @[Switch.scala 41:52:@23479.4]
  assign output_11_11 = io_outValid_11 & _T_62320; // @[Switch.scala 41:38:@23480.4]
  assign _T_62323 = select_12 == 6'hb; // @[Switch.scala 41:52:@23482.4]
  assign output_11_12 = io_outValid_12 & _T_62323; // @[Switch.scala 41:38:@23483.4]
  assign _T_62326 = select_13 == 6'hb; // @[Switch.scala 41:52:@23485.4]
  assign output_11_13 = io_outValid_13 & _T_62326; // @[Switch.scala 41:38:@23486.4]
  assign _T_62329 = select_14 == 6'hb; // @[Switch.scala 41:52:@23488.4]
  assign output_11_14 = io_outValid_14 & _T_62329; // @[Switch.scala 41:38:@23489.4]
  assign _T_62332 = select_15 == 6'hb; // @[Switch.scala 41:52:@23491.4]
  assign output_11_15 = io_outValid_15 & _T_62332; // @[Switch.scala 41:38:@23492.4]
  assign _T_62335 = select_16 == 6'hb; // @[Switch.scala 41:52:@23494.4]
  assign output_11_16 = io_outValid_16 & _T_62335; // @[Switch.scala 41:38:@23495.4]
  assign _T_62338 = select_17 == 6'hb; // @[Switch.scala 41:52:@23497.4]
  assign output_11_17 = io_outValid_17 & _T_62338; // @[Switch.scala 41:38:@23498.4]
  assign _T_62341 = select_18 == 6'hb; // @[Switch.scala 41:52:@23500.4]
  assign output_11_18 = io_outValid_18 & _T_62341; // @[Switch.scala 41:38:@23501.4]
  assign _T_62344 = select_19 == 6'hb; // @[Switch.scala 41:52:@23503.4]
  assign output_11_19 = io_outValid_19 & _T_62344; // @[Switch.scala 41:38:@23504.4]
  assign _T_62347 = select_20 == 6'hb; // @[Switch.scala 41:52:@23506.4]
  assign output_11_20 = io_outValid_20 & _T_62347; // @[Switch.scala 41:38:@23507.4]
  assign _T_62350 = select_21 == 6'hb; // @[Switch.scala 41:52:@23509.4]
  assign output_11_21 = io_outValid_21 & _T_62350; // @[Switch.scala 41:38:@23510.4]
  assign _T_62353 = select_22 == 6'hb; // @[Switch.scala 41:52:@23512.4]
  assign output_11_22 = io_outValid_22 & _T_62353; // @[Switch.scala 41:38:@23513.4]
  assign _T_62356 = select_23 == 6'hb; // @[Switch.scala 41:52:@23515.4]
  assign output_11_23 = io_outValid_23 & _T_62356; // @[Switch.scala 41:38:@23516.4]
  assign _T_62359 = select_24 == 6'hb; // @[Switch.scala 41:52:@23518.4]
  assign output_11_24 = io_outValid_24 & _T_62359; // @[Switch.scala 41:38:@23519.4]
  assign _T_62362 = select_25 == 6'hb; // @[Switch.scala 41:52:@23521.4]
  assign output_11_25 = io_outValid_25 & _T_62362; // @[Switch.scala 41:38:@23522.4]
  assign _T_62365 = select_26 == 6'hb; // @[Switch.scala 41:52:@23524.4]
  assign output_11_26 = io_outValid_26 & _T_62365; // @[Switch.scala 41:38:@23525.4]
  assign _T_62368 = select_27 == 6'hb; // @[Switch.scala 41:52:@23527.4]
  assign output_11_27 = io_outValid_27 & _T_62368; // @[Switch.scala 41:38:@23528.4]
  assign _T_62371 = select_28 == 6'hb; // @[Switch.scala 41:52:@23530.4]
  assign output_11_28 = io_outValid_28 & _T_62371; // @[Switch.scala 41:38:@23531.4]
  assign _T_62374 = select_29 == 6'hb; // @[Switch.scala 41:52:@23533.4]
  assign output_11_29 = io_outValid_29 & _T_62374; // @[Switch.scala 41:38:@23534.4]
  assign _T_62377 = select_30 == 6'hb; // @[Switch.scala 41:52:@23536.4]
  assign output_11_30 = io_outValid_30 & _T_62377; // @[Switch.scala 41:38:@23537.4]
  assign _T_62380 = select_31 == 6'hb; // @[Switch.scala 41:52:@23539.4]
  assign output_11_31 = io_outValid_31 & _T_62380; // @[Switch.scala 41:38:@23540.4]
  assign _T_62383 = select_32 == 6'hb; // @[Switch.scala 41:52:@23542.4]
  assign output_11_32 = io_outValid_32 & _T_62383; // @[Switch.scala 41:38:@23543.4]
  assign _T_62386 = select_33 == 6'hb; // @[Switch.scala 41:52:@23545.4]
  assign output_11_33 = io_outValid_33 & _T_62386; // @[Switch.scala 41:38:@23546.4]
  assign _T_62389 = select_34 == 6'hb; // @[Switch.scala 41:52:@23548.4]
  assign output_11_34 = io_outValid_34 & _T_62389; // @[Switch.scala 41:38:@23549.4]
  assign _T_62392 = select_35 == 6'hb; // @[Switch.scala 41:52:@23551.4]
  assign output_11_35 = io_outValid_35 & _T_62392; // @[Switch.scala 41:38:@23552.4]
  assign _T_62395 = select_36 == 6'hb; // @[Switch.scala 41:52:@23554.4]
  assign output_11_36 = io_outValid_36 & _T_62395; // @[Switch.scala 41:38:@23555.4]
  assign _T_62398 = select_37 == 6'hb; // @[Switch.scala 41:52:@23557.4]
  assign output_11_37 = io_outValid_37 & _T_62398; // @[Switch.scala 41:38:@23558.4]
  assign _T_62401 = select_38 == 6'hb; // @[Switch.scala 41:52:@23560.4]
  assign output_11_38 = io_outValid_38 & _T_62401; // @[Switch.scala 41:38:@23561.4]
  assign _T_62404 = select_39 == 6'hb; // @[Switch.scala 41:52:@23563.4]
  assign output_11_39 = io_outValid_39 & _T_62404; // @[Switch.scala 41:38:@23564.4]
  assign _T_62407 = select_40 == 6'hb; // @[Switch.scala 41:52:@23566.4]
  assign output_11_40 = io_outValid_40 & _T_62407; // @[Switch.scala 41:38:@23567.4]
  assign _T_62410 = select_41 == 6'hb; // @[Switch.scala 41:52:@23569.4]
  assign output_11_41 = io_outValid_41 & _T_62410; // @[Switch.scala 41:38:@23570.4]
  assign _T_62413 = select_42 == 6'hb; // @[Switch.scala 41:52:@23572.4]
  assign output_11_42 = io_outValid_42 & _T_62413; // @[Switch.scala 41:38:@23573.4]
  assign _T_62416 = select_43 == 6'hb; // @[Switch.scala 41:52:@23575.4]
  assign output_11_43 = io_outValid_43 & _T_62416; // @[Switch.scala 41:38:@23576.4]
  assign _T_62419 = select_44 == 6'hb; // @[Switch.scala 41:52:@23578.4]
  assign output_11_44 = io_outValid_44 & _T_62419; // @[Switch.scala 41:38:@23579.4]
  assign _T_62422 = select_45 == 6'hb; // @[Switch.scala 41:52:@23581.4]
  assign output_11_45 = io_outValid_45 & _T_62422; // @[Switch.scala 41:38:@23582.4]
  assign _T_62425 = select_46 == 6'hb; // @[Switch.scala 41:52:@23584.4]
  assign output_11_46 = io_outValid_46 & _T_62425; // @[Switch.scala 41:38:@23585.4]
  assign _T_62428 = select_47 == 6'hb; // @[Switch.scala 41:52:@23587.4]
  assign output_11_47 = io_outValid_47 & _T_62428; // @[Switch.scala 41:38:@23588.4]
  assign _T_62431 = select_48 == 6'hb; // @[Switch.scala 41:52:@23590.4]
  assign output_11_48 = io_outValid_48 & _T_62431; // @[Switch.scala 41:38:@23591.4]
  assign _T_62434 = select_49 == 6'hb; // @[Switch.scala 41:52:@23593.4]
  assign output_11_49 = io_outValid_49 & _T_62434; // @[Switch.scala 41:38:@23594.4]
  assign _T_62437 = select_50 == 6'hb; // @[Switch.scala 41:52:@23596.4]
  assign output_11_50 = io_outValid_50 & _T_62437; // @[Switch.scala 41:38:@23597.4]
  assign _T_62440 = select_51 == 6'hb; // @[Switch.scala 41:52:@23599.4]
  assign output_11_51 = io_outValid_51 & _T_62440; // @[Switch.scala 41:38:@23600.4]
  assign _T_62443 = select_52 == 6'hb; // @[Switch.scala 41:52:@23602.4]
  assign output_11_52 = io_outValid_52 & _T_62443; // @[Switch.scala 41:38:@23603.4]
  assign _T_62446 = select_53 == 6'hb; // @[Switch.scala 41:52:@23605.4]
  assign output_11_53 = io_outValid_53 & _T_62446; // @[Switch.scala 41:38:@23606.4]
  assign _T_62449 = select_54 == 6'hb; // @[Switch.scala 41:52:@23608.4]
  assign output_11_54 = io_outValid_54 & _T_62449; // @[Switch.scala 41:38:@23609.4]
  assign _T_62452 = select_55 == 6'hb; // @[Switch.scala 41:52:@23611.4]
  assign output_11_55 = io_outValid_55 & _T_62452; // @[Switch.scala 41:38:@23612.4]
  assign _T_62455 = select_56 == 6'hb; // @[Switch.scala 41:52:@23614.4]
  assign output_11_56 = io_outValid_56 & _T_62455; // @[Switch.scala 41:38:@23615.4]
  assign _T_62458 = select_57 == 6'hb; // @[Switch.scala 41:52:@23617.4]
  assign output_11_57 = io_outValid_57 & _T_62458; // @[Switch.scala 41:38:@23618.4]
  assign _T_62461 = select_58 == 6'hb; // @[Switch.scala 41:52:@23620.4]
  assign output_11_58 = io_outValid_58 & _T_62461; // @[Switch.scala 41:38:@23621.4]
  assign _T_62464 = select_59 == 6'hb; // @[Switch.scala 41:52:@23623.4]
  assign output_11_59 = io_outValid_59 & _T_62464; // @[Switch.scala 41:38:@23624.4]
  assign _T_62467 = select_60 == 6'hb; // @[Switch.scala 41:52:@23626.4]
  assign output_11_60 = io_outValid_60 & _T_62467; // @[Switch.scala 41:38:@23627.4]
  assign _T_62470 = select_61 == 6'hb; // @[Switch.scala 41:52:@23629.4]
  assign output_11_61 = io_outValid_61 & _T_62470; // @[Switch.scala 41:38:@23630.4]
  assign _T_62473 = select_62 == 6'hb; // @[Switch.scala 41:52:@23632.4]
  assign output_11_62 = io_outValid_62 & _T_62473; // @[Switch.scala 41:38:@23633.4]
  assign _T_62476 = select_63 == 6'hb; // @[Switch.scala 41:52:@23635.4]
  assign output_11_63 = io_outValid_63 & _T_62476; // @[Switch.scala 41:38:@23636.4]
  assign _T_62484 = {output_11_7,output_11_6,output_11_5,output_11_4,output_11_3,output_11_2,output_11_1,output_11_0}; // @[Switch.scala 43:31:@23644.4]
  assign _T_62492 = {output_11_15,output_11_14,output_11_13,output_11_12,output_11_11,output_11_10,output_11_9,output_11_8,_T_62484}; // @[Switch.scala 43:31:@23652.4]
  assign _T_62499 = {output_11_23,output_11_22,output_11_21,output_11_20,output_11_19,output_11_18,output_11_17,output_11_16}; // @[Switch.scala 43:31:@23659.4]
  assign _T_62508 = {output_11_31,output_11_30,output_11_29,output_11_28,output_11_27,output_11_26,output_11_25,output_11_24,_T_62499,_T_62492}; // @[Switch.scala 43:31:@23668.4]
  assign _T_62515 = {output_11_39,output_11_38,output_11_37,output_11_36,output_11_35,output_11_34,output_11_33,output_11_32}; // @[Switch.scala 43:31:@23675.4]
  assign _T_62523 = {output_11_47,output_11_46,output_11_45,output_11_44,output_11_43,output_11_42,output_11_41,output_11_40,_T_62515}; // @[Switch.scala 43:31:@23683.4]
  assign _T_62530 = {output_11_55,output_11_54,output_11_53,output_11_52,output_11_51,output_11_50,output_11_49,output_11_48}; // @[Switch.scala 43:31:@23690.4]
  assign _T_62539 = {output_11_63,output_11_62,output_11_61,output_11_60,output_11_59,output_11_58,output_11_57,output_11_56,_T_62530,_T_62523}; // @[Switch.scala 43:31:@23699.4]
  assign _T_62540 = {_T_62539,_T_62508}; // @[Switch.scala 43:31:@23700.4]
  assign _T_62544 = select_0 == 6'hc; // @[Switch.scala 41:52:@23703.4]
  assign output_12_0 = io_outValid_0 & _T_62544; // @[Switch.scala 41:38:@23704.4]
  assign _T_62547 = select_1 == 6'hc; // @[Switch.scala 41:52:@23706.4]
  assign output_12_1 = io_outValid_1 & _T_62547; // @[Switch.scala 41:38:@23707.4]
  assign _T_62550 = select_2 == 6'hc; // @[Switch.scala 41:52:@23709.4]
  assign output_12_2 = io_outValid_2 & _T_62550; // @[Switch.scala 41:38:@23710.4]
  assign _T_62553 = select_3 == 6'hc; // @[Switch.scala 41:52:@23712.4]
  assign output_12_3 = io_outValid_3 & _T_62553; // @[Switch.scala 41:38:@23713.4]
  assign _T_62556 = select_4 == 6'hc; // @[Switch.scala 41:52:@23715.4]
  assign output_12_4 = io_outValid_4 & _T_62556; // @[Switch.scala 41:38:@23716.4]
  assign _T_62559 = select_5 == 6'hc; // @[Switch.scala 41:52:@23718.4]
  assign output_12_5 = io_outValid_5 & _T_62559; // @[Switch.scala 41:38:@23719.4]
  assign _T_62562 = select_6 == 6'hc; // @[Switch.scala 41:52:@23721.4]
  assign output_12_6 = io_outValid_6 & _T_62562; // @[Switch.scala 41:38:@23722.4]
  assign _T_62565 = select_7 == 6'hc; // @[Switch.scala 41:52:@23724.4]
  assign output_12_7 = io_outValid_7 & _T_62565; // @[Switch.scala 41:38:@23725.4]
  assign _T_62568 = select_8 == 6'hc; // @[Switch.scala 41:52:@23727.4]
  assign output_12_8 = io_outValid_8 & _T_62568; // @[Switch.scala 41:38:@23728.4]
  assign _T_62571 = select_9 == 6'hc; // @[Switch.scala 41:52:@23730.4]
  assign output_12_9 = io_outValid_9 & _T_62571; // @[Switch.scala 41:38:@23731.4]
  assign _T_62574 = select_10 == 6'hc; // @[Switch.scala 41:52:@23733.4]
  assign output_12_10 = io_outValid_10 & _T_62574; // @[Switch.scala 41:38:@23734.4]
  assign _T_62577 = select_11 == 6'hc; // @[Switch.scala 41:52:@23736.4]
  assign output_12_11 = io_outValid_11 & _T_62577; // @[Switch.scala 41:38:@23737.4]
  assign _T_62580 = select_12 == 6'hc; // @[Switch.scala 41:52:@23739.4]
  assign output_12_12 = io_outValid_12 & _T_62580; // @[Switch.scala 41:38:@23740.4]
  assign _T_62583 = select_13 == 6'hc; // @[Switch.scala 41:52:@23742.4]
  assign output_12_13 = io_outValid_13 & _T_62583; // @[Switch.scala 41:38:@23743.4]
  assign _T_62586 = select_14 == 6'hc; // @[Switch.scala 41:52:@23745.4]
  assign output_12_14 = io_outValid_14 & _T_62586; // @[Switch.scala 41:38:@23746.4]
  assign _T_62589 = select_15 == 6'hc; // @[Switch.scala 41:52:@23748.4]
  assign output_12_15 = io_outValid_15 & _T_62589; // @[Switch.scala 41:38:@23749.4]
  assign _T_62592 = select_16 == 6'hc; // @[Switch.scala 41:52:@23751.4]
  assign output_12_16 = io_outValid_16 & _T_62592; // @[Switch.scala 41:38:@23752.4]
  assign _T_62595 = select_17 == 6'hc; // @[Switch.scala 41:52:@23754.4]
  assign output_12_17 = io_outValid_17 & _T_62595; // @[Switch.scala 41:38:@23755.4]
  assign _T_62598 = select_18 == 6'hc; // @[Switch.scala 41:52:@23757.4]
  assign output_12_18 = io_outValid_18 & _T_62598; // @[Switch.scala 41:38:@23758.4]
  assign _T_62601 = select_19 == 6'hc; // @[Switch.scala 41:52:@23760.4]
  assign output_12_19 = io_outValid_19 & _T_62601; // @[Switch.scala 41:38:@23761.4]
  assign _T_62604 = select_20 == 6'hc; // @[Switch.scala 41:52:@23763.4]
  assign output_12_20 = io_outValid_20 & _T_62604; // @[Switch.scala 41:38:@23764.4]
  assign _T_62607 = select_21 == 6'hc; // @[Switch.scala 41:52:@23766.4]
  assign output_12_21 = io_outValid_21 & _T_62607; // @[Switch.scala 41:38:@23767.4]
  assign _T_62610 = select_22 == 6'hc; // @[Switch.scala 41:52:@23769.4]
  assign output_12_22 = io_outValid_22 & _T_62610; // @[Switch.scala 41:38:@23770.4]
  assign _T_62613 = select_23 == 6'hc; // @[Switch.scala 41:52:@23772.4]
  assign output_12_23 = io_outValid_23 & _T_62613; // @[Switch.scala 41:38:@23773.4]
  assign _T_62616 = select_24 == 6'hc; // @[Switch.scala 41:52:@23775.4]
  assign output_12_24 = io_outValid_24 & _T_62616; // @[Switch.scala 41:38:@23776.4]
  assign _T_62619 = select_25 == 6'hc; // @[Switch.scala 41:52:@23778.4]
  assign output_12_25 = io_outValid_25 & _T_62619; // @[Switch.scala 41:38:@23779.4]
  assign _T_62622 = select_26 == 6'hc; // @[Switch.scala 41:52:@23781.4]
  assign output_12_26 = io_outValid_26 & _T_62622; // @[Switch.scala 41:38:@23782.4]
  assign _T_62625 = select_27 == 6'hc; // @[Switch.scala 41:52:@23784.4]
  assign output_12_27 = io_outValid_27 & _T_62625; // @[Switch.scala 41:38:@23785.4]
  assign _T_62628 = select_28 == 6'hc; // @[Switch.scala 41:52:@23787.4]
  assign output_12_28 = io_outValid_28 & _T_62628; // @[Switch.scala 41:38:@23788.4]
  assign _T_62631 = select_29 == 6'hc; // @[Switch.scala 41:52:@23790.4]
  assign output_12_29 = io_outValid_29 & _T_62631; // @[Switch.scala 41:38:@23791.4]
  assign _T_62634 = select_30 == 6'hc; // @[Switch.scala 41:52:@23793.4]
  assign output_12_30 = io_outValid_30 & _T_62634; // @[Switch.scala 41:38:@23794.4]
  assign _T_62637 = select_31 == 6'hc; // @[Switch.scala 41:52:@23796.4]
  assign output_12_31 = io_outValid_31 & _T_62637; // @[Switch.scala 41:38:@23797.4]
  assign _T_62640 = select_32 == 6'hc; // @[Switch.scala 41:52:@23799.4]
  assign output_12_32 = io_outValid_32 & _T_62640; // @[Switch.scala 41:38:@23800.4]
  assign _T_62643 = select_33 == 6'hc; // @[Switch.scala 41:52:@23802.4]
  assign output_12_33 = io_outValid_33 & _T_62643; // @[Switch.scala 41:38:@23803.4]
  assign _T_62646 = select_34 == 6'hc; // @[Switch.scala 41:52:@23805.4]
  assign output_12_34 = io_outValid_34 & _T_62646; // @[Switch.scala 41:38:@23806.4]
  assign _T_62649 = select_35 == 6'hc; // @[Switch.scala 41:52:@23808.4]
  assign output_12_35 = io_outValid_35 & _T_62649; // @[Switch.scala 41:38:@23809.4]
  assign _T_62652 = select_36 == 6'hc; // @[Switch.scala 41:52:@23811.4]
  assign output_12_36 = io_outValid_36 & _T_62652; // @[Switch.scala 41:38:@23812.4]
  assign _T_62655 = select_37 == 6'hc; // @[Switch.scala 41:52:@23814.4]
  assign output_12_37 = io_outValid_37 & _T_62655; // @[Switch.scala 41:38:@23815.4]
  assign _T_62658 = select_38 == 6'hc; // @[Switch.scala 41:52:@23817.4]
  assign output_12_38 = io_outValid_38 & _T_62658; // @[Switch.scala 41:38:@23818.4]
  assign _T_62661 = select_39 == 6'hc; // @[Switch.scala 41:52:@23820.4]
  assign output_12_39 = io_outValid_39 & _T_62661; // @[Switch.scala 41:38:@23821.4]
  assign _T_62664 = select_40 == 6'hc; // @[Switch.scala 41:52:@23823.4]
  assign output_12_40 = io_outValid_40 & _T_62664; // @[Switch.scala 41:38:@23824.4]
  assign _T_62667 = select_41 == 6'hc; // @[Switch.scala 41:52:@23826.4]
  assign output_12_41 = io_outValid_41 & _T_62667; // @[Switch.scala 41:38:@23827.4]
  assign _T_62670 = select_42 == 6'hc; // @[Switch.scala 41:52:@23829.4]
  assign output_12_42 = io_outValid_42 & _T_62670; // @[Switch.scala 41:38:@23830.4]
  assign _T_62673 = select_43 == 6'hc; // @[Switch.scala 41:52:@23832.4]
  assign output_12_43 = io_outValid_43 & _T_62673; // @[Switch.scala 41:38:@23833.4]
  assign _T_62676 = select_44 == 6'hc; // @[Switch.scala 41:52:@23835.4]
  assign output_12_44 = io_outValid_44 & _T_62676; // @[Switch.scala 41:38:@23836.4]
  assign _T_62679 = select_45 == 6'hc; // @[Switch.scala 41:52:@23838.4]
  assign output_12_45 = io_outValid_45 & _T_62679; // @[Switch.scala 41:38:@23839.4]
  assign _T_62682 = select_46 == 6'hc; // @[Switch.scala 41:52:@23841.4]
  assign output_12_46 = io_outValid_46 & _T_62682; // @[Switch.scala 41:38:@23842.4]
  assign _T_62685 = select_47 == 6'hc; // @[Switch.scala 41:52:@23844.4]
  assign output_12_47 = io_outValid_47 & _T_62685; // @[Switch.scala 41:38:@23845.4]
  assign _T_62688 = select_48 == 6'hc; // @[Switch.scala 41:52:@23847.4]
  assign output_12_48 = io_outValid_48 & _T_62688; // @[Switch.scala 41:38:@23848.4]
  assign _T_62691 = select_49 == 6'hc; // @[Switch.scala 41:52:@23850.4]
  assign output_12_49 = io_outValid_49 & _T_62691; // @[Switch.scala 41:38:@23851.4]
  assign _T_62694 = select_50 == 6'hc; // @[Switch.scala 41:52:@23853.4]
  assign output_12_50 = io_outValid_50 & _T_62694; // @[Switch.scala 41:38:@23854.4]
  assign _T_62697 = select_51 == 6'hc; // @[Switch.scala 41:52:@23856.4]
  assign output_12_51 = io_outValid_51 & _T_62697; // @[Switch.scala 41:38:@23857.4]
  assign _T_62700 = select_52 == 6'hc; // @[Switch.scala 41:52:@23859.4]
  assign output_12_52 = io_outValid_52 & _T_62700; // @[Switch.scala 41:38:@23860.4]
  assign _T_62703 = select_53 == 6'hc; // @[Switch.scala 41:52:@23862.4]
  assign output_12_53 = io_outValid_53 & _T_62703; // @[Switch.scala 41:38:@23863.4]
  assign _T_62706 = select_54 == 6'hc; // @[Switch.scala 41:52:@23865.4]
  assign output_12_54 = io_outValid_54 & _T_62706; // @[Switch.scala 41:38:@23866.4]
  assign _T_62709 = select_55 == 6'hc; // @[Switch.scala 41:52:@23868.4]
  assign output_12_55 = io_outValid_55 & _T_62709; // @[Switch.scala 41:38:@23869.4]
  assign _T_62712 = select_56 == 6'hc; // @[Switch.scala 41:52:@23871.4]
  assign output_12_56 = io_outValid_56 & _T_62712; // @[Switch.scala 41:38:@23872.4]
  assign _T_62715 = select_57 == 6'hc; // @[Switch.scala 41:52:@23874.4]
  assign output_12_57 = io_outValid_57 & _T_62715; // @[Switch.scala 41:38:@23875.4]
  assign _T_62718 = select_58 == 6'hc; // @[Switch.scala 41:52:@23877.4]
  assign output_12_58 = io_outValid_58 & _T_62718; // @[Switch.scala 41:38:@23878.4]
  assign _T_62721 = select_59 == 6'hc; // @[Switch.scala 41:52:@23880.4]
  assign output_12_59 = io_outValid_59 & _T_62721; // @[Switch.scala 41:38:@23881.4]
  assign _T_62724 = select_60 == 6'hc; // @[Switch.scala 41:52:@23883.4]
  assign output_12_60 = io_outValid_60 & _T_62724; // @[Switch.scala 41:38:@23884.4]
  assign _T_62727 = select_61 == 6'hc; // @[Switch.scala 41:52:@23886.4]
  assign output_12_61 = io_outValid_61 & _T_62727; // @[Switch.scala 41:38:@23887.4]
  assign _T_62730 = select_62 == 6'hc; // @[Switch.scala 41:52:@23889.4]
  assign output_12_62 = io_outValid_62 & _T_62730; // @[Switch.scala 41:38:@23890.4]
  assign _T_62733 = select_63 == 6'hc; // @[Switch.scala 41:52:@23892.4]
  assign output_12_63 = io_outValid_63 & _T_62733; // @[Switch.scala 41:38:@23893.4]
  assign _T_62741 = {output_12_7,output_12_6,output_12_5,output_12_4,output_12_3,output_12_2,output_12_1,output_12_0}; // @[Switch.scala 43:31:@23901.4]
  assign _T_62749 = {output_12_15,output_12_14,output_12_13,output_12_12,output_12_11,output_12_10,output_12_9,output_12_8,_T_62741}; // @[Switch.scala 43:31:@23909.4]
  assign _T_62756 = {output_12_23,output_12_22,output_12_21,output_12_20,output_12_19,output_12_18,output_12_17,output_12_16}; // @[Switch.scala 43:31:@23916.4]
  assign _T_62765 = {output_12_31,output_12_30,output_12_29,output_12_28,output_12_27,output_12_26,output_12_25,output_12_24,_T_62756,_T_62749}; // @[Switch.scala 43:31:@23925.4]
  assign _T_62772 = {output_12_39,output_12_38,output_12_37,output_12_36,output_12_35,output_12_34,output_12_33,output_12_32}; // @[Switch.scala 43:31:@23932.4]
  assign _T_62780 = {output_12_47,output_12_46,output_12_45,output_12_44,output_12_43,output_12_42,output_12_41,output_12_40,_T_62772}; // @[Switch.scala 43:31:@23940.4]
  assign _T_62787 = {output_12_55,output_12_54,output_12_53,output_12_52,output_12_51,output_12_50,output_12_49,output_12_48}; // @[Switch.scala 43:31:@23947.4]
  assign _T_62796 = {output_12_63,output_12_62,output_12_61,output_12_60,output_12_59,output_12_58,output_12_57,output_12_56,_T_62787,_T_62780}; // @[Switch.scala 43:31:@23956.4]
  assign _T_62797 = {_T_62796,_T_62765}; // @[Switch.scala 43:31:@23957.4]
  assign _T_62801 = select_0 == 6'hd; // @[Switch.scala 41:52:@23960.4]
  assign output_13_0 = io_outValid_0 & _T_62801; // @[Switch.scala 41:38:@23961.4]
  assign _T_62804 = select_1 == 6'hd; // @[Switch.scala 41:52:@23963.4]
  assign output_13_1 = io_outValid_1 & _T_62804; // @[Switch.scala 41:38:@23964.4]
  assign _T_62807 = select_2 == 6'hd; // @[Switch.scala 41:52:@23966.4]
  assign output_13_2 = io_outValid_2 & _T_62807; // @[Switch.scala 41:38:@23967.4]
  assign _T_62810 = select_3 == 6'hd; // @[Switch.scala 41:52:@23969.4]
  assign output_13_3 = io_outValid_3 & _T_62810; // @[Switch.scala 41:38:@23970.4]
  assign _T_62813 = select_4 == 6'hd; // @[Switch.scala 41:52:@23972.4]
  assign output_13_4 = io_outValid_4 & _T_62813; // @[Switch.scala 41:38:@23973.4]
  assign _T_62816 = select_5 == 6'hd; // @[Switch.scala 41:52:@23975.4]
  assign output_13_5 = io_outValid_5 & _T_62816; // @[Switch.scala 41:38:@23976.4]
  assign _T_62819 = select_6 == 6'hd; // @[Switch.scala 41:52:@23978.4]
  assign output_13_6 = io_outValid_6 & _T_62819; // @[Switch.scala 41:38:@23979.4]
  assign _T_62822 = select_7 == 6'hd; // @[Switch.scala 41:52:@23981.4]
  assign output_13_7 = io_outValid_7 & _T_62822; // @[Switch.scala 41:38:@23982.4]
  assign _T_62825 = select_8 == 6'hd; // @[Switch.scala 41:52:@23984.4]
  assign output_13_8 = io_outValid_8 & _T_62825; // @[Switch.scala 41:38:@23985.4]
  assign _T_62828 = select_9 == 6'hd; // @[Switch.scala 41:52:@23987.4]
  assign output_13_9 = io_outValid_9 & _T_62828; // @[Switch.scala 41:38:@23988.4]
  assign _T_62831 = select_10 == 6'hd; // @[Switch.scala 41:52:@23990.4]
  assign output_13_10 = io_outValid_10 & _T_62831; // @[Switch.scala 41:38:@23991.4]
  assign _T_62834 = select_11 == 6'hd; // @[Switch.scala 41:52:@23993.4]
  assign output_13_11 = io_outValid_11 & _T_62834; // @[Switch.scala 41:38:@23994.4]
  assign _T_62837 = select_12 == 6'hd; // @[Switch.scala 41:52:@23996.4]
  assign output_13_12 = io_outValid_12 & _T_62837; // @[Switch.scala 41:38:@23997.4]
  assign _T_62840 = select_13 == 6'hd; // @[Switch.scala 41:52:@23999.4]
  assign output_13_13 = io_outValid_13 & _T_62840; // @[Switch.scala 41:38:@24000.4]
  assign _T_62843 = select_14 == 6'hd; // @[Switch.scala 41:52:@24002.4]
  assign output_13_14 = io_outValid_14 & _T_62843; // @[Switch.scala 41:38:@24003.4]
  assign _T_62846 = select_15 == 6'hd; // @[Switch.scala 41:52:@24005.4]
  assign output_13_15 = io_outValid_15 & _T_62846; // @[Switch.scala 41:38:@24006.4]
  assign _T_62849 = select_16 == 6'hd; // @[Switch.scala 41:52:@24008.4]
  assign output_13_16 = io_outValid_16 & _T_62849; // @[Switch.scala 41:38:@24009.4]
  assign _T_62852 = select_17 == 6'hd; // @[Switch.scala 41:52:@24011.4]
  assign output_13_17 = io_outValid_17 & _T_62852; // @[Switch.scala 41:38:@24012.4]
  assign _T_62855 = select_18 == 6'hd; // @[Switch.scala 41:52:@24014.4]
  assign output_13_18 = io_outValid_18 & _T_62855; // @[Switch.scala 41:38:@24015.4]
  assign _T_62858 = select_19 == 6'hd; // @[Switch.scala 41:52:@24017.4]
  assign output_13_19 = io_outValid_19 & _T_62858; // @[Switch.scala 41:38:@24018.4]
  assign _T_62861 = select_20 == 6'hd; // @[Switch.scala 41:52:@24020.4]
  assign output_13_20 = io_outValid_20 & _T_62861; // @[Switch.scala 41:38:@24021.4]
  assign _T_62864 = select_21 == 6'hd; // @[Switch.scala 41:52:@24023.4]
  assign output_13_21 = io_outValid_21 & _T_62864; // @[Switch.scala 41:38:@24024.4]
  assign _T_62867 = select_22 == 6'hd; // @[Switch.scala 41:52:@24026.4]
  assign output_13_22 = io_outValid_22 & _T_62867; // @[Switch.scala 41:38:@24027.4]
  assign _T_62870 = select_23 == 6'hd; // @[Switch.scala 41:52:@24029.4]
  assign output_13_23 = io_outValid_23 & _T_62870; // @[Switch.scala 41:38:@24030.4]
  assign _T_62873 = select_24 == 6'hd; // @[Switch.scala 41:52:@24032.4]
  assign output_13_24 = io_outValid_24 & _T_62873; // @[Switch.scala 41:38:@24033.4]
  assign _T_62876 = select_25 == 6'hd; // @[Switch.scala 41:52:@24035.4]
  assign output_13_25 = io_outValid_25 & _T_62876; // @[Switch.scala 41:38:@24036.4]
  assign _T_62879 = select_26 == 6'hd; // @[Switch.scala 41:52:@24038.4]
  assign output_13_26 = io_outValid_26 & _T_62879; // @[Switch.scala 41:38:@24039.4]
  assign _T_62882 = select_27 == 6'hd; // @[Switch.scala 41:52:@24041.4]
  assign output_13_27 = io_outValid_27 & _T_62882; // @[Switch.scala 41:38:@24042.4]
  assign _T_62885 = select_28 == 6'hd; // @[Switch.scala 41:52:@24044.4]
  assign output_13_28 = io_outValid_28 & _T_62885; // @[Switch.scala 41:38:@24045.4]
  assign _T_62888 = select_29 == 6'hd; // @[Switch.scala 41:52:@24047.4]
  assign output_13_29 = io_outValid_29 & _T_62888; // @[Switch.scala 41:38:@24048.4]
  assign _T_62891 = select_30 == 6'hd; // @[Switch.scala 41:52:@24050.4]
  assign output_13_30 = io_outValid_30 & _T_62891; // @[Switch.scala 41:38:@24051.4]
  assign _T_62894 = select_31 == 6'hd; // @[Switch.scala 41:52:@24053.4]
  assign output_13_31 = io_outValid_31 & _T_62894; // @[Switch.scala 41:38:@24054.4]
  assign _T_62897 = select_32 == 6'hd; // @[Switch.scala 41:52:@24056.4]
  assign output_13_32 = io_outValid_32 & _T_62897; // @[Switch.scala 41:38:@24057.4]
  assign _T_62900 = select_33 == 6'hd; // @[Switch.scala 41:52:@24059.4]
  assign output_13_33 = io_outValid_33 & _T_62900; // @[Switch.scala 41:38:@24060.4]
  assign _T_62903 = select_34 == 6'hd; // @[Switch.scala 41:52:@24062.4]
  assign output_13_34 = io_outValid_34 & _T_62903; // @[Switch.scala 41:38:@24063.4]
  assign _T_62906 = select_35 == 6'hd; // @[Switch.scala 41:52:@24065.4]
  assign output_13_35 = io_outValid_35 & _T_62906; // @[Switch.scala 41:38:@24066.4]
  assign _T_62909 = select_36 == 6'hd; // @[Switch.scala 41:52:@24068.4]
  assign output_13_36 = io_outValid_36 & _T_62909; // @[Switch.scala 41:38:@24069.4]
  assign _T_62912 = select_37 == 6'hd; // @[Switch.scala 41:52:@24071.4]
  assign output_13_37 = io_outValid_37 & _T_62912; // @[Switch.scala 41:38:@24072.4]
  assign _T_62915 = select_38 == 6'hd; // @[Switch.scala 41:52:@24074.4]
  assign output_13_38 = io_outValid_38 & _T_62915; // @[Switch.scala 41:38:@24075.4]
  assign _T_62918 = select_39 == 6'hd; // @[Switch.scala 41:52:@24077.4]
  assign output_13_39 = io_outValid_39 & _T_62918; // @[Switch.scala 41:38:@24078.4]
  assign _T_62921 = select_40 == 6'hd; // @[Switch.scala 41:52:@24080.4]
  assign output_13_40 = io_outValid_40 & _T_62921; // @[Switch.scala 41:38:@24081.4]
  assign _T_62924 = select_41 == 6'hd; // @[Switch.scala 41:52:@24083.4]
  assign output_13_41 = io_outValid_41 & _T_62924; // @[Switch.scala 41:38:@24084.4]
  assign _T_62927 = select_42 == 6'hd; // @[Switch.scala 41:52:@24086.4]
  assign output_13_42 = io_outValid_42 & _T_62927; // @[Switch.scala 41:38:@24087.4]
  assign _T_62930 = select_43 == 6'hd; // @[Switch.scala 41:52:@24089.4]
  assign output_13_43 = io_outValid_43 & _T_62930; // @[Switch.scala 41:38:@24090.4]
  assign _T_62933 = select_44 == 6'hd; // @[Switch.scala 41:52:@24092.4]
  assign output_13_44 = io_outValid_44 & _T_62933; // @[Switch.scala 41:38:@24093.4]
  assign _T_62936 = select_45 == 6'hd; // @[Switch.scala 41:52:@24095.4]
  assign output_13_45 = io_outValid_45 & _T_62936; // @[Switch.scala 41:38:@24096.4]
  assign _T_62939 = select_46 == 6'hd; // @[Switch.scala 41:52:@24098.4]
  assign output_13_46 = io_outValid_46 & _T_62939; // @[Switch.scala 41:38:@24099.4]
  assign _T_62942 = select_47 == 6'hd; // @[Switch.scala 41:52:@24101.4]
  assign output_13_47 = io_outValid_47 & _T_62942; // @[Switch.scala 41:38:@24102.4]
  assign _T_62945 = select_48 == 6'hd; // @[Switch.scala 41:52:@24104.4]
  assign output_13_48 = io_outValid_48 & _T_62945; // @[Switch.scala 41:38:@24105.4]
  assign _T_62948 = select_49 == 6'hd; // @[Switch.scala 41:52:@24107.4]
  assign output_13_49 = io_outValid_49 & _T_62948; // @[Switch.scala 41:38:@24108.4]
  assign _T_62951 = select_50 == 6'hd; // @[Switch.scala 41:52:@24110.4]
  assign output_13_50 = io_outValid_50 & _T_62951; // @[Switch.scala 41:38:@24111.4]
  assign _T_62954 = select_51 == 6'hd; // @[Switch.scala 41:52:@24113.4]
  assign output_13_51 = io_outValid_51 & _T_62954; // @[Switch.scala 41:38:@24114.4]
  assign _T_62957 = select_52 == 6'hd; // @[Switch.scala 41:52:@24116.4]
  assign output_13_52 = io_outValid_52 & _T_62957; // @[Switch.scala 41:38:@24117.4]
  assign _T_62960 = select_53 == 6'hd; // @[Switch.scala 41:52:@24119.4]
  assign output_13_53 = io_outValid_53 & _T_62960; // @[Switch.scala 41:38:@24120.4]
  assign _T_62963 = select_54 == 6'hd; // @[Switch.scala 41:52:@24122.4]
  assign output_13_54 = io_outValid_54 & _T_62963; // @[Switch.scala 41:38:@24123.4]
  assign _T_62966 = select_55 == 6'hd; // @[Switch.scala 41:52:@24125.4]
  assign output_13_55 = io_outValid_55 & _T_62966; // @[Switch.scala 41:38:@24126.4]
  assign _T_62969 = select_56 == 6'hd; // @[Switch.scala 41:52:@24128.4]
  assign output_13_56 = io_outValid_56 & _T_62969; // @[Switch.scala 41:38:@24129.4]
  assign _T_62972 = select_57 == 6'hd; // @[Switch.scala 41:52:@24131.4]
  assign output_13_57 = io_outValid_57 & _T_62972; // @[Switch.scala 41:38:@24132.4]
  assign _T_62975 = select_58 == 6'hd; // @[Switch.scala 41:52:@24134.4]
  assign output_13_58 = io_outValid_58 & _T_62975; // @[Switch.scala 41:38:@24135.4]
  assign _T_62978 = select_59 == 6'hd; // @[Switch.scala 41:52:@24137.4]
  assign output_13_59 = io_outValid_59 & _T_62978; // @[Switch.scala 41:38:@24138.4]
  assign _T_62981 = select_60 == 6'hd; // @[Switch.scala 41:52:@24140.4]
  assign output_13_60 = io_outValid_60 & _T_62981; // @[Switch.scala 41:38:@24141.4]
  assign _T_62984 = select_61 == 6'hd; // @[Switch.scala 41:52:@24143.4]
  assign output_13_61 = io_outValid_61 & _T_62984; // @[Switch.scala 41:38:@24144.4]
  assign _T_62987 = select_62 == 6'hd; // @[Switch.scala 41:52:@24146.4]
  assign output_13_62 = io_outValid_62 & _T_62987; // @[Switch.scala 41:38:@24147.4]
  assign _T_62990 = select_63 == 6'hd; // @[Switch.scala 41:52:@24149.4]
  assign output_13_63 = io_outValid_63 & _T_62990; // @[Switch.scala 41:38:@24150.4]
  assign _T_62998 = {output_13_7,output_13_6,output_13_5,output_13_4,output_13_3,output_13_2,output_13_1,output_13_0}; // @[Switch.scala 43:31:@24158.4]
  assign _T_63006 = {output_13_15,output_13_14,output_13_13,output_13_12,output_13_11,output_13_10,output_13_9,output_13_8,_T_62998}; // @[Switch.scala 43:31:@24166.4]
  assign _T_63013 = {output_13_23,output_13_22,output_13_21,output_13_20,output_13_19,output_13_18,output_13_17,output_13_16}; // @[Switch.scala 43:31:@24173.4]
  assign _T_63022 = {output_13_31,output_13_30,output_13_29,output_13_28,output_13_27,output_13_26,output_13_25,output_13_24,_T_63013,_T_63006}; // @[Switch.scala 43:31:@24182.4]
  assign _T_63029 = {output_13_39,output_13_38,output_13_37,output_13_36,output_13_35,output_13_34,output_13_33,output_13_32}; // @[Switch.scala 43:31:@24189.4]
  assign _T_63037 = {output_13_47,output_13_46,output_13_45,output_13_44,output_13_43,output_13_42,output_13_41,output_13_40,_T_63029}; // @[Switch.scala 43:31:@24197.4]
  assign _T_63044 = {output_13_55,output_13_54,output_13_53,output_13_52,output_13_51,output_13_50,output_13_49,output_13_48}; // @[Switch.scala 43:31:@24204.4]
  assign _T_63053 = {output_13_63,output_13_62,output_13_61,output_13_60,output_13_59,output_13_58,output_13_57,output_13_56,_T_63044,_T_63037}; // @[Switch.scala 43:31:@24213.4]
  assign _T_63054 = {_T_63053,_T_63022}; // @[Switch.scala 43:31:@24214.4]
  assign _T_63058 = select_0 == 6'he; // @[Switch.scala 41:52:@24217.4]
  assign output_14_0 = io_outValid_0 & _T_63058; // @[Switch.scala 41:38:@24218.4]
  assign _T_63061 = select_1 == 6'he; // @[Switch.scala 41:52:@24220.4]
  assign output_14_1 = io_outValid_1 & _T_63061; // @[Switch.scala 41:38:@24221.4]
  assign _T_63064 = select_2 == 6'he; // @[Switch.scala 41:52:@24223.4]
  assign output_14_2 = io_outValid_2 & _T_63064; // @[Switch.scala 41:38:@24224.4]
  assign _T_63067 = select_3 == 6'he; // @[Switch.scala 41:52:@24226.4]
  assign output_14_3 = io_outValid_3 & _T_63067; // @[Switch.scala 41:38:@24227.4]
  assign _T_63070 = select_4 == 6'he; // @[Switch.scala 41:52:@24229.4]
  assign output_14_4 = io_outValid_4 & _T_63070; // @[Switch.scala 41:38:@24230.4]
  assign _T_63073 = select_5 == 6'he; // @[Switch.scala 41:52:@24232.4]
  assign output_14_5 = io_outValid_5 & _T_63073; // @[Switch.scala 41:38:@24233.4]
  assign _T_63076 = select_6 == 6'he; // @[Switch.scala 41:52:@24235.4]
  assign output_14_6 = io_outValid_6 & _T_63076; // @[Switch.scala 41:38:@24236.4]
  assign _T_63079 = select_7 == 6'he; // @[Switch.scala 41:52:@24238.4]
  assign output_14_7 = io_outValid_7 & _T_63079; // @[Switch.scala 41:38:@24239.4]
  assign _T_63082 = select_8 == 6'he; // @[Switch.scala 41:52:@24241.4]
  assign output_14_8 = io_outValid_8 & _T_63082; // @[Switch.scala 41:38:@24242.4]
  assign _T_63085 = select_9 == 6'he; // @[Switch.scala 41:52:@24244.4]
  assign output_14_9 = io_outValid_9 & _T_63085; // @[Switch.scala 41:38:@24245.4]
  assign _T_63088 = select_10 == 6'he; // @[Switch.scala 41:52:@24247.4]
  assign output_14_10 = io_outValid_10 & _T_63088; // @[Switch.scala 41:38:@24248.4]
  assign _T_63091 = select_11 == 6'he; // @[Switch.scala 41:52:@24250.4]
  assign output_14_11 = io_outValid_11 & _T_63091; // @[Switch.scala 41:38:@24251.4]
  assign _T_63094 = select_12 == 6'he; // @[Switch.scala 41:52:@24253.4]
  assign output_14_12 = io_outValid_12 & _T_63094; // @[Switch.scala 41:38:@24254.4]
  assign _T_63097 = select_13 == 6'he; // @[Switch.scala 41:52:@24256.4]
  assign output_14_13 = io_outValid_13 & _T_63097; // @[Switch.scala 41:38:@24257.4]
  assign _T_63100 = select_14 == 6'he; // @[Switch.scala 41:52:@24259.4]
  assign output_14_14 = io_outValid_14 & _T_63100; // @[Switch.scala 41:38:@24260.4]
  assign _T_63103 = select_15 == 6'he; // @[Switch.scala 41:52:@24262.4]
  assign output_14_15 = io_outValid_15 & _T_63103; // @[Switch.scala 41:38:@24263.4]
  assign _T_63106 = select_16 == 6'he; // @[Switch.scala 41:52:@24265.4]
  assign output_14_16 = io_outValid_16 & _T_63106; // @[Switch.scala 41:38:@24266.4]
  assign _T_63109 = select_17 == 6'he; // @[Switch.scala 41:52:@24268.4]
  assign output_14_17 = io_outValid_17 & _T_63109; // @[Switch.scala 41:38:@24269.4]
  assign _T_63112 = select_18 == 6'he; // @[Switch.scala 41:52:@24271.4]
  assign output_14_18 = io_outValid_18 & _T_63112; // @[Switch.scala 41:38:@24272.4]
  assign _T_63115 = select_19 == 6'he; // @[Switch.scala 41:52:@24274.4]
  assign output_14_19 = io_outValid_19 & _T_63115; // @[Switch.scala 41:38:@24275.4]
  assign _T_63118 = select_20 == 6'he; // @[Switch.scala 41:52:@24277.4]
  assign output_14_20 = io_outValid_20 & _T_63118; // @[Switch.scala 41:38:@24278.4]
  assign _T_63121 = select_21 == 6'he; // @[Switch.scala 41:52:@24280.4]
  assign output_14_21 = io_outValid_21 & _T_63121; // @[Switch.scala 41:38:@24281.4]
  assign _T_63124 = select_22 == 6'he; // @[Switch.scala 41:52:@24283.4]
  assign output_14_22 = io_outValid_22 & _T_63124; // @[Switch.scala 41:38:@24284.4]
  assign _T_63127 = select_23 == 6'he; // @[Switch.scala 41:52:@24286.4]
  assign output_14_23 = io_outValid_23 & _T_63127; // @[Switch.scala 41:38:@24287.4]
  assign _T_63130 = select_24 == 6'he; // @[Switch.scala 41:52:@24289.4]
  assign output_14_24 = io_outValid_24 & _T_63130; // @[Switch.scala 41:38:@24290.4]
  assign _T_63133 = select_25 == 6'he; // @[Switch.scala 41:52:@24292.4]
  assign output_14_25 = io_outValid_25 & _T_63133; // @[Switch.scala 41:38:@24293.4]
  assign _T_63136 = select_26 == 6'he; // @[Switch.scala 41:52:@24295.4]
  assign output_14_26 = io_outValid_26 & _T_63136; // @[Switch.scala 41:38:@24296.4]
  assign _T_63139 = select_27 == 6'he; // @[Switch.scala 41:52:@24298.4]
  assign output_14_27 = io_outValid_27 & _T_63139; // @[Switch.scala 41:38:@24299.4]
  assign _T_63142 = select_28 == 6'he; // @[Switch.scala 41:52:@24301.4]
  assign output_14_28 = io_outValid_28 & _T_63142; // @[Switch.scala 41:38:@24302.4]
  assign _T_63145 = select_29 == 6'he; // @[Switch.scala 41:52:@24304.4]
  assign output_14_29 = io_outValid_29 & _T_63145; // @[Switch.scala 41:38:@24305.4]
  assign _T_63148 = select_30 == 6'he; // @[Switch.scala 41:52:@24307.4]
  assign output_14_30 = io_outValid_30 & _T_63148; // @[Switch.scala 41:38:@24308.4]
  assign _T_63151 = select_31 == 6'he; // @[Switch.scala 41:52:@24310.4]
  assign output_14_31 = io_outValid_31 & _T_63151; // @[Switch.scala 41:38:@24311.4]
  assign _T_63154 = select_32 == 6'he; // @[Switch.scala 41:52:@24313.4]
  assign output_14_32 = io_outValid_32 & _T_63154; // @[Switch.scala 41:38:@24314.4]
  assign _T_63157 = select_33 == 6'he; // @[Switch.scala 41:52:@24316.4]
  assign output_14_33 = io_outValid_33 & _T_63157; // @[Switch.scala 41:38:@24317.4]
  assign _T_63160 = select_34 == 6'he; // @[Switch.scala 41:52:@24319.4]
  assign output_14_34 = io_outValid_34 & _T_63160; // @[Switch.scala 41:38:@24320.4]
  assign _T_63163 = select_35 == 6'he; // @[Switch.scala 41:52:@24322.4]
  assign output_14_35 = io_outValid_35 & _T_63163; // @[Switch.scala 41:38:@24323.4]
  assign _T_63166 = select_36 == 6'he; // @[Switch.scala 41:52:@24325.4]
  assign output_14_36 = io_outValid_36 & _T_63166; // @[Switch.scala 41:38:@24326.4]
  assign _T_63169 = select_37 == 6'he; // @[Switch.scala 41:52:@24328.4]
  assign output_14_37 = io_outValid_37 & _T_63169; // @[Switch.scala 41:38:@24329.4]
  assign _T_63172 = select_38 == 6'he; // @[Switch.scala 41:52:@24331.4]
  assign output_14_38 = io_outValid_38 & _T_63172; // @[Switch.scala 41:38:@24332.4]
  assign _T_63175 = select_39 == 6'he; // @[Switch.scala 41:52:@24334.4]
  assign output_14_39 = io_outValid_39 & _T_63175; // @[Switch.scala 41:38:@24335.4]
  assign _T_63178 = select_40 == 6'he; // @[Switch.scala 41:52:@24337.4]
  assign output_14_40 = io_outValid_40 & _T_63178; // @[Switch.scala 41:38:@24338.4]
  assign _T_63181 = select_41 == 6'he; // @[Switch.scala 41:52:@24340.4]
  assign output_14_41 = io_outValid_41 & _T_63181; // @[Switch.scala 41:38:@24341.4]
  assign _T_63184 = select_42 == 6'he; // @[Switch.scala 41:52:@24343.4]
  assign output_14_42 = io_outValid_42 & _T_63184; // @[Switch.scala 41:38:@24344.4]
  assign _T_63187 = select_43 == 6'he; // @[Switch.scala 41:52:@24346.4]
  assign output_14_43 = io_outValid_43 & _T_63187; // @[Switch.scala 41:38:@24347.4]
  assign _T_63190 = select_44 == 6'he; // @[Switch.scala 41:52:@24349.4]
  assign output_14_44 = io_outValid_44 & _T_63190; // @[Switch.scala 41:38:@24350.4]
  assign _T_63193 = select_45 == 6'he; // @[Switch.scala 41:52:@24352.4]
  assign output_14_45 = io_outValid_45 & _T_63193; // @[Switch.scala 41:38:@24353.4]
  assign _T_63196 = select_46 == 6'he; // @[Switch.scala 41:52:@24355.4]
  assign output_14_46 = io_outValid_46 & _T_63196; // @[Switch.scala 41:38:@24356.4]
  assign _T_63199 = select_47 == 6'he; // @[Switch.scala 41:52:@24358.4]
  assign output_14_47 = io_outValid_47 & _T_63199; // @[Switch.scala 41:38:@24359.4]
  assign _T_63202 = select_48 == 6'he; // @[Switch.scala 41:52:@24361.4]
  assign output_14_48 = io_outValid_48 & _T_63202; // @[Switch.scala 41:38:@24362.4]
  assign _T_63205 = select_49 == 6'he; // @[Switch.scala 41:52:@24364.4]
  assign output_14_49 = io_outValid_49 & _T_63205; // @[Switch.scala 41:38:@24365.4]
  assign _T_63208 = select_50 == 6'he; // @[Switch.scala 41:52:@24367.4]
  assign output_14_50 = io_outValid_50 & _T_63208; // @[Switch.scala 41:38:@24368.4]
  assign _T_63211 = select_51 == 6'he; // @[Switch.scala 41:52:@24370.4]
  assign output_14_51 = io_outValid_51 & _T_63211; // @[Switch.scala 41:38:@24371.4]
  assign _T_63214 = select_52 == 6'he; // @[Switch.scala 41:52:@24373.4]
  assign output_14_52 = io_outValid_52 & _T_63214; // @[Switch.scala 41:38:@24374.4]
  assign _T_63217 = select_53 == 6'he; // @[Switch.scala 41:52:@24376.4]
  assign output_14_53 = io_outValid_53 & _T_63217; // @[Switch.scala 41:38:@24377.4]
  assign _T_63220 = select_54 == 6'he; // @[Switch.scala 41:52:@24379.4]
  assign output_14_54 = io_outValid_54 & _T_63220; // @[Switch.scala 41:38:@24380.4]
  assign _T_63223 = select_55 == 6'he; // @[Switch.scala 41:52:@24382.4]
  assign output_14_55 = io_outValid_55 & _T_63223; // @[Switch.scala 41:38:@24383.4]
  assign _T_63226 = select_56 == 6'he; // @[Switch.scala 41:52:@24385.4]
  assign output_14_56 = io_outValid_56 & _T_63226; // @[Switch.scala 41:38:@24386.4]
  assign _T_63229 = select_57 == 6'he; // @[Switch.scala 41:52:@24388.4]
  assign output_14_57 = io_outValid_57 & _T_63229; // @[Switch.scala 41:38:@24389.4]
  assign _T_63232 = select_58 == 6'he; // @[Switch.scala 41:52:@24391.4]
  assign output_14_58 = io_outValid_58 & _T_63232; // @[Switch.scala 41:38:@24392.4]
  assign _T_63235 = select_59 == 6'he; // @[Switch.scala 41:52:@24394.4]
  assign output_14_59 = io_outValid_59 & _T_63235; // @[Switch.scala 41:38:@24395.4]
  assign _T_63238 = select_60 == 6'he; // @[Switch.scala 41:52:@24397.4]
  assign output_14_60 = io_outValid_60 & _T_63238; // @[Switch.scala 41:38:@24398.4]
  assign _T_63241 = select_61 == 6'he; // @[Switch.scala 41:52:@24400.4]
  assign output_14_61 = io_outValid_61 & _T_63241; // @[Switch.scala 41:38:@24401.4]
  assign _T_63244 = select_62 == 6'he; // @[Switch.scala 41:52:@24403.4]
  assign output_14_62 = io_outValid_62 & _T_63244; // @[Switch.scala 41:38:@24404.4]
  assign _T_63247 = select_63 == 6'he; // @[Switch.scala 41:52:@24406.4]
  assign output_14_63 = io_outValid_63 & _T_63247; // @[Switch.scala 41:38:@24407.4]
  assign _T_63255 = {output_14_7,output_14_6,output_14_5,output_14_4,output_14_3,output_14_2,output_14_1,output_14_0}; // @[Switch.scala 43:31:@24415.4]
  assign _T_63263 = {output_14_15,output_14_14,output_14_13,output_14_12,output_14_11,output_14_10,output_14_9,output_14_8,_T_63255}; // @[Switch.scala 43:31:@24423.4]
  assign _T_63270 = {output_14_23,output_14_22,output_14_21,output_14_20,output_14_19,output_14_18,output_14_17,output_14_16}; // @[Switch.scala 43:31:@24430.4]
  assign _T_63279 = {output_14_31,output_14_30,output_14_29,output_14_28,output_14_27,output_14_26,output_14_25,output_14_24,_T_63270,_T_63263}; // @[Switch.scala 43:31:@24439.4]
  assign _T_63286 = {output_14_39,output_14_38,output_14_37,output_14_36,output_14_35,output_14_34,output_14_33,output_14_32}; // @[Switch.scala 43:31:@24446.4]
  assign _T_63294 = {output_14_47,output_14_46,output_14_45,output_14_44,output_14_43,output_14_42,output_14_41,output_14_40,_T_63286}; // @[Switch.scala 43:31:@24454.4]
  assign _T_63301 = {output_14_55,output_14_54,output_14_53,output_14_52,output_14_51,output_14_50,output_14_49,output_14_48}; // @[Switch.scala 43:31:@24461.4]
  assign _T_63310 = {output_14_63,output_14_62,output_14_61,output_14_60,output_14_59,output_14_58,output_14_57,output_14_56,_T_63301,_T_63294}; // @[Switch.scala 43:31:@24470.4]
  assign _T_63311 = {_T_63310,_T_63279}; // @[Switch.scala 43:31:@24471.4]
  assign _T_63315 = select_0 == 6'hf; // @[Switch.scala 41:52:@24474.4]
  assign output_15_0 = io_outValid_0 & _T_63315; // @[Switch.scala 41:38:@24475.4]
  assign _T_63318 = select_1 == 6'hf; // @[Switch.scala 41:52:@24477.4]
  assign output_15_1 = io_outValid_1 & _T_63318; // @[Switch.scala 41:38:@24478.4]
  assign _T_63321 = select_2 == 6'hf; // @[Switch.scala 41:52:@24480.4]
  assign output_15_2 = io_outValid_2 & _T_63321; // @[Switch.scala 41:38:@24481.4]
  assign _T_63324 = select_3 == 6'hf; // @[Switch.scala 41:52:@24483.4]
  assign output_15_3 = io_outValid_3 & _T_63324; // @[Switch.scala 41:38:@24484.4]
  assign _T_63327 = select_4 == 6'hf; // @[Switch.scala 41:52:@24486.4]
  assign output_15_4 = io_outValid_4 & _T_63327; // @[Switch.scala 41:38:@24487.4]
  assign _T_63330 = select_5 == 6'hf; // @[Switch.scala 41:52:@24489.4]
  assign output_15_5 = io_outValid_5 & _T_63330; // @[Switch.scala 41:38:@24490.4]
  assign _T_63333 = select_6 == 6'hf; // @[Switch.scala 41:52:@24492.4]
  assign output_15_6 = io_outValid_6 & _T_63333; // @[Switch.scala 41:38:@24493.4]
  assign _T_63336 = select_7 == 6'hf; // @[Switch.scala 41:52:@24495.4]
  assign output_15_7 = io_outValid_7 & _T_63336; // @[Switch.scala 41:38:@24496.4]
  assign _T_63339 = select_8 == 6'hf; // @[Switch.scala 41:52:@24498.4]
  assign output_15_8 = io_outValid_8 & _T_63339; // @[Switch.scala 41:38:@24499.4]
  assign _T_63342 = select_9 == 6'hf; // @[Switch.scala 41:52:@24501.4]
  assign output_15_9 = io_outValid_9 & _T_63342; // @[Switch.scala 41:38:@24502.4]
  assign _T_63345 = select_10 == 6'hf; // @[Switch.scala 41:52:@24504.4]
  assign output_15_10 = io_outValid_10 & _T_63345; // @[Switch.scala 41:38:@24505.4]
  assign _T_63348 = select_11 == 6'hf; // @[Switch.scala 41:52:@24507.4]
  assign output_15_11 = io_outValid_11 & _T_63348; // @[Switch.scala 41:38:@24508.4]
  assign _T_63351 = select_12 == 6'hf; // @[Switch.scala 41:52:@24510.4]
  assign output_15_12 = io_outValid_12 & _T_63351; // @[Switch.scala 41:38:@24511.4]
  assign _T_63354 = select_13 == 6'hf; // @[Switch.scala 41:52:@24513.4]
  assign output_15_13 = io_outValid_13 & _T_63354; // @[Switch.scala 41:38:@24514.4]
  assign _T_63357 = select_14 == 6'hf; // @[Switch.scala 41:52:@24516.4]
  assign output_15_14 = io_outValid_14 & _T_63357; // @[Switch.scala 41:38:@24517.4]
  assign _T_63360 = select_15 == 6'hf; // @[Switch.scala 41:52:@24519.4]
  assign output_15_15 = io_outValid_15 & _T_63360; // @[Switch.scala 41:38:@24520.4]
  assign _T_63363 = select_16 == 6'hf; // @[Switch.scala 41:52:@24522.4]
  assign output_15_16 = io_outValid_16 & _T_63363; // @[Switch.scala 41:38:@24523.4]
  assign _T_63366 = select_17 == 6'hf; // @[Switch.scala 41:52:@24525.4]
  assign output_15_17 = io_outValid_17 & _T_63366; // @[Switch.scala 41:38:@24526.4]
  assign _T_63369 = select_18 == 6'hf; // @[Switch.scala 41:52:@24528.4]
  assign output_15_18 = io_outValid_18 & _T_63369; // @[Switch.scala 41:38:@24529.4]
  assign _T_63372 = select_19 == 6'hf; // @[Switch.scala 41:52:@24531.4]
  assign output_15_19 = io_outValid_19 & _T_63372; // @[Switch.scala 41:38:@24532.4]
  assign _T_63375 = select_20 == 6'hf; // @[Switch.scala 41:52:@24534.4]
  assign output_15_20 = io_outValid_20 & _T_63375; // @[Switch.scala 41:38:@24535.4]
  assign _T_63378 = select_21 == 6'hf; // @[Switch.scala 41:52:@24537.4]
  assign output_15_21 = io_outValid_21 & _T_63378; // @[Switch.scala 41:38:@24538.4]
  assign _T_63381 = select_22 == 6'hf; // @[Switch.scala 41:52:@24540.4]
  assign output_15_22 = io_outValid_22 & _T_63381; // @[Switch.scala 41:38:@24541.4]
  assign _T_63384 = select_23 == 6'hf; // @[Switch.scala 41:52:@24543.4]
  assign output_15_23 = io_outValid_23 & _T_63384; // @[Switch.scala 41:38:@24544.4]
  assign _T_63387 = select_24 == 6'hf; // @[Switch.scala 41:52:@24546.4]
  assign output_15_24 = io_outValid_24 & _T_63387; // @[Switch.scala 41:38:@24547.4]
  assign _T_63390 = select_25 == 6'hf; // @[Switch.scala 41:52:@24549.4]
  assign output_15_25 = io_outValid_25 & _T_63390; // @[Switch.scala 41:38:@24550.4]
  assign _T_63393 = select_26 == 6'hf; // @[Switch.scala 41:52:@24552.4]
  assign output_15_26 = io_outValid_26 & _T_63393; // @[Switch.scala 41:38:@24553.4]
  assign _T_63396 = select_27 == 6'hf; // @[Switch.scala 41:52:@24555.4]
  assign output_15_27 = io_outValid_27 & _T_63396; // @[Switch.scala 41:38:@24556.4]
  assign _T_63399 = select_28 == 6'hf; // @[Switch.scala 41:52:@24558.4]
  assign output_15_28 = io_outValid_28 & _T_63399; // @[Switch.scala 41:38:@24559.4]
  assign _T_63402 = select_29 == 6'hf; // @[Switch.scala 41:52:@24561.4]
  assign output_15_29 = io_outValid_29 & _T_63402; // @[Switch.scala 41:38:@24562.4]
  assign _T_63405 = select_30 == 6'hf; // @[Switch.scala 41:52:@24564.4]
  assign output_15_30 = io_outValid_30 & _T_63405; // @[Switch.scala 41:38:@24565.4]
  assign _T_63408 = select_31 == 6'hf; // @[Switch.scala 41:52:@24567.4]
  assign output_15_31 = io_outValid_31 & _T_63408; // @[Switch.scala 41:38:@24568.4]
  assign _T_63411 = select_32 == 6'hf; // @[Switch.scala 41:52:@24570.4]
  assign output_15_32 = io_outValid_32 & _T_63411; // @[Switch.scala 41:38:@24571.4]
  assign _T_63414 = select_33 == 6'hf; // @[Switch.scala 41:52:@24573.4]
  assign output_15_33 = io_outValid_33 & _T_63414; // @[Switch.scala 41:38:@24574.4]
  assign _T_63417 = select_34 == 6'hf; // @[Switch.scala 41:52:@24576.4]
  assign output_15_34 = io_outValid_34 & _T_63417; // @[Switch.scala 41:38:@24577.4]
  assign _T_63420 = select_35 == 6'hf; // @[Switch.scala 41:52:@24579.4]
  assign output_15_35 = io_outValid_35 & _T_63420; // @[Switch.scala 41:38:@24580.4]
  assign _T_63423 = select_36 == 6'hf; // @[Switch.scala 41:52:@24582.4]
  assign output_15_36 = io_outValid_36 & _T_63423; // @[Switch.scala 41:38:@24583.4]
  assign _T_63426 = select_37 == 6'hf; // @[Switch.scala 41:52:@24585.4]
  assign output_15_37 = io_outValid_37 & _T_63426; // @[Switch.scala 41:38:@24586.4]
  assign _T_63429 = select_38 == 6'hf; // @[Switch.scala 41:52:@24588.4]
  assign output_15_38 = io_outValid_38 & _T_63429; // @[Switch.scala 41:38:@24589.4]
  assign _T_63432 = select_39 == 6'hf; // @[Switch.scala 41:52:@24591.4]
  assign output_15_39 = io_outValid_39 & _T_63432; // @[Switch.scala 41:38:@24592.4]
  assign _T_63435 = select_40 == 6'hf; // @[Switch.scala 41:52:@24594.4]
  assign output_15_40 = io_outValid_40 & _T_63435; // @[Switch.scala 41:38:@24595.4]
  assign _T_63438 = select_41 == 6'hf; // @[Switch.scala 41:52:@24597.4]
  assign output_15_41 = io_outValid_41 & _T_63438; // @[Switch.scala 41:38:@24598.4]
  assign _T_63441 = select_42 == 6'hf; // @[Switch.scala 41:52:@24600.4]
  assign output_15_42 = io_outValid_42 & _T_63441; // @[Switch.scala 41:38:@24601.4]
  assign _T_63444 = select_43 == 6'hf; // @[Switch.scala 41:52:@24603.4]
  assign output_15_43 = io_outValid_43 & _T_63444; // @[Switch.scala 41:38:@24604.4]
  assign _T_63447 = select_44 == 6'hf; // @[Switch.scala 41:52:@24606.4]
  assign output_15_44 = io_outValid_44 & _T_63447; // @[Switch.scala 41:38:@24607.4]
  assign _T_63450 = select_45 == 6'hf; // @[Switch.scala 41:52:@24609.4]
  assign output_15_45 = io_outValid_45 & _T_63450; // @[Switch.scala 41:38:@24610.4]
  assign _T_63453 = select_46 == 6'hf; // @[Switch.scala 41:52:@24612.4]
  assign output_15_46 = io_outValid_46 & _T_63453; // @[Switch.scala 41:38:@24613.4]
  assign _T_63456 = select_47 == 6'hf; // @[Switch.scala 41:52:@24615.4]
  assign output_15_47 = io_outValid_47 & _T_63456; // @[Switch.scala 41:38:@24616.4]
  assign _T_63459 = select_48 == 6'hf; // @[Switch.scala 41:52:@24618.4]
  assign output_15_48 = io_outValid_48 & _T_63459; // @[Switch.scala 41:38:@24619.4]
  assign _T_63462 = select_49 == 6'hf; // @[Switch.scala 41:52:@24621.4]
  assign output_15_49 = io_outValid_49 & _T_63462; // @[Switch.scala 41:38:@24622.4]
  assign _T_63465 = select_50 == 6'hf; // @[Switch.scala 41:52:@24624.4]
  assign output_15_50 = io_outValid_50 & _T_63465; // @[Switch.scala 41:38:@24625.4]
  assign _T_63468 = select_51 == 6'hf; // @[Switch.scala 41:52:@24627.4]
  assign output_15_51 = io_outValid_51 & _T_63468; // @[Switch.scala 41:38:@24628.4]
  assign _T_63471 = select_52 == 6'hf; // @[Switch.scala 41:52:@24630.4]
  assign output_15_52 = io_outValid_52 & _T_63471; // @[Switch.scala 41:38:@24631.4]
  assign _T_63474 = select_53 == 6'hf; // @[Switch.scala 41:52:@24633.4]
  assign output_15_53 = io_outValid_53 & _T_63474; // @[Switch.scala 41:38:@24634.4]
  assign _T_63477 = select_54 == 6'hf; // @[Switch.scala 41:52:@24636.4]
  assign output_15_54 = io_outValid_54 & _T_63477; // @[Switch.scala 41:38:@24637.4]
  assign _T_63480 = select_55 == 6'hf; // @[Switch.scala 41:52:@24639.4]
  assign output_15_55 = io_outValid_55 & _T_63480; // @[Switch.scala 41:38:@24640.4]
  assign _T_63483 = select_56 == 6'hf; // @[Switch.scala 41:52:@24642.4]
  assign output_15_56 = io_outValid_56 & _T_63483; // @[Switch.scala 41:38:@24643.4]
  assign _T_63486 = select_57 == 6'hf; // @[Switch.scala 41:52:@24645.4]
  assign output_15_57 = io_outValid_57 & _T_63486; // @[Switch.scala 41:38:@24646.4]
  assign _T_63489 = select_58 == 6'hf; // @[Switch.scala 41:52:@24648.4]
  assign output_15_58 = io_outValid_58 & _T_63489; // @[Switch.scala 41:38:@24649.4]
  assign _T_63492 = select_59 == 6'hf; // @[Switch.scala 41:52:@24651.4]
  assign output_15_59 = io_outValid_59 & _T_63492; // @[Switch.scala 41:38:@24652.4]
  assign _T_63495 = select_60 == 6'hf; // @[Switch.scala 41:52:@24654.4]
  assign output_15_60 = io_outValid_60 & _T_63495; // @[Switch.scala 41:38:@24655.4]
  assign _T_63498 = select_61 == 6'hf; // @[Switch.scala 41:52:@24657.4]
  assign output_15_61 = io_outValid_61 & _T_63498; // @[Switch.scala 41:38:@24658.4]
  assign _T_63501 = select_62 == 6'hf; // @[Switch.scala 41:52:@24660.4]
  assign output_15_62 = io_outValid_62 & _T_63501; // @[Switch.scala 41:38:@24661.4]
  assign _T_63504 = select_63 == 6'hf; // @[Switch.scala 41:52:@24663.4]
  assign output_15_63 = io_outValid_63 & _T_63504; // @[Switch.scala 41:38:@24664.4]
  assign _T_63512 = {output_15_7,output_15_6,output_15_5,output_15_4,output_15_3,output_15_2,output_15_1,output_15_0}; // @[Switch.scala 43:31:@24672.4]
  assign _T_63520 = {output_15_15,output_15_14,output_15_13,output_15_12,output_15_11,output_15_10,output_15_9,output_15_8,_T_63512}; // @[Switch.scala 43:31:@24680.4]
  assign _T_63527 = {output_15_23,output_15_22,output_15_21,output_15_20,output_15_19,output_15_18,output_15_17,output_15_16}; // @[Switch.scala 43:31:@24687.4]
  assign _T_63536 = {output_15_31,output_15_30,output_15_29,output_15_28,output_15_27,output_15_26,output_15_25,output_15_24,_T_63527,_T_63520}; // @[Switch.scala 43:31:@24696.4]
  assign _T_63543 = {output_15_39,output_15_38,output_15_37,output_15_36,output_15_35,output_15_34,output_15_33,output_15_32}; // @[Switch.scala 43:31:@24703.4]
  assign _T_63551 = {output_15_47,output_15_46,output_15_45,output_15_44,output_15_43,output_15_42,output_15_41,output_15_40,_T_63543}; // @[Switch.scala 43:31:@24711.4]
  assign _T_63558 = {output_15_55,output_15_54,output_15_53,output_15_52,output_15_51,output_15_50,output_15_49,output_15_48}; // @[Switch.scala 43:31:@24718.4]
  assign _T_63567 = {output_15_63,output_15_62,output_15_61,output_15_60,output_15_59,output_15_58,output_15_57,output_15_56,_T_63558,_T_63551}; // @[Switch.scala 43:31:@24727.4]
  assign _T_63568 = {_T_63567,_T_63536}; // @[Switch.scala 43:31:@24728.4]
  assign _T_63572 = select_0 == 6'h10; // @[Switch.scala 41:52:@24731.4]
  assign output_16_0 = io_outValid_0 & _T_63572; // @[Switch.scala 41:38:@24732.4]
  assign _T_63575 = select_1 == 6'h10; // @[Switch.scala 41:52:@24734.4]
  assign output_16_1 = io_outValid_1 & _T_63575; // @[Switch.scala 41:38:@24735.4]
  assign _T_63578 = select_2 == 6'h10; // @[Switch.scala 41:52:@24737.4]
  assign output_16_2 = io_outValid_2 & _T_63578; // @[Switch.scala 41:38:@24738.4]
  assign _T_63581 = select_3 == 6'h10; // @[Switch.scala 41:52:@24740.4]
  assign output_16_3 = io_outValid_3 & _T_63581; // @[Switch.scala 41:38:@24741.4]
  assign _T_63584 = select_4 == 6'h10; // @[Switch.scala 41:52:@24743.4]
  assign output_16_4 = io_outValid_4 & _T_63584; // @[Switch.scala 41:38:@24744.4]
  assign _T_63587 = select_5 == 6'h10; // @[Switch.scala 41:52:@24746.4]
  assign output_16_5 = io_outValid_5 & _T_63587; // @[Switch.scala 41:38:@24747.4]
  assign _T_63590 = select_6 == 6'h10; // @[Switch.scala 41:52:@24749.4]
  assign output_16_6 = io_outValid_6 & _T_63590; // @[Switch.scala 41:38:@24750.4]
  assign _T_63593 = select_7 == 6'h10; // @[Switch.scala 41:52:@24752.4]
  assign output_16_7 = io_outValid_7 & _T_63593; // @[Switch.scala 41:38:@24753.4]
  assign _T_63596 = select_8 == 6'h10; // @[Switch.scala 41:52:@24755.4]
  assign output_16_8 = io_outValid_8 & _T_63596; // @[Switch.scala 41:38:@24756.4]
  assign _T_63599 = select_9 == 6'h10; // @[Switch.scala 41:52:@24758.4]
  assign output_16_9 = io_outValid_9 & _T_63599; // @[Switch.scala 41:38:@24759.4]
  assign _T_63602 = select_10 == 6'h10; // @[Switch.scala 41:52:@24761.4]
  assign output_16_10 = io_outValid_10 & _T_63602; // @[Switch.scala 41:38:@24762.4]
  assign _T_63605 = select_11 == 6'h10; // @[Switch.scala 41:52:@24764.4]
  assign output_16_11 = io_outValid_11 & _T_63605; // @[Switch.scala 41:38:@24765.4]
  assign _T_63608 = select_12 == 6'h10; // @[Switch.scala 41:52:@24767.4]
  assign output_16_12 = io_outValid_12 & _T_63608; // @[Switch.scala 41:38:@24768.4]
  assign _T_63611 = select_13 == 6'h10; // @[Switch.scala 41:52:@24770.4]
  assign output_16_13 = io_outValid_13 & _T_63611; // @[Switch.scala 41:38:@24771.4]
  assign _T_63614 = select_14 == 6'h10; // @[Switch.scala 41:52:@24773.4]
  assign output_16_14 = io_outValid_14 & _T_63614; // @[Switch.scala 41:38:@24774.4]
  assign _T_63617 = select_15 == 6'h10; // @[Switch.scala 41:52:@24776.4]
  assign output_16_15 = io_outValid_15 & _T_63617; // @[Switch.scala 41:38:@24777.4]
  assign _T_63620 = select_16 == 6'h10; // @[Switch.scala 41:52:@24779.4]
  assign output_16_16 = io_outValid_16 & _T_63620; // @[Switch.scala 41:38:@24780.4]
  assign _T_63623 = select_17 == 6'h10; // @[Switch.scala 41:52:@24782.4]
  assign output_16_17 = io_outValid_17 & _T_63623; // @[Switch.scala 41:38:@24783.4]
  assign _T_63626 = select_18 == 6'h10; // @[Switch.scala 41:52:@24785.4]
  assign output_16_18 = io_outValid_18 & _T_63626; // @[Switch.scala 41:38:@24786.4]
  assign _T_63629 = select_19 == 6'h10; // @[Switch.scala 41:52:@24788.4]
  assign output_16_19 = io_outValid_19 & _T_63629; // @[Switch.scala 41:38:@24789.4]
  assign _T_63632 = select_20 == 6'h10; // @[Switch.scala 41:52:@24791.4]
  assign output_16_20 = io_outValid_20 & _T_63632; // @[Switch.scala 41:38:@24792.4]
  assign _T_63635 = select_21 == 6'h10; // @[Switch.scala 41:52:@24794.4]
  assign output_16_21 = io_outValid_21 & _T_63635; // @[Switch.scala 41:38:@24795.4]
  assign _T_63638 = select_22 == 6'h10; // @[Switch.scala 41:52:@24797.4]
  assign output_16_22 = io_outValid_22 & _T_63638; // @[Switch.scala 41:38:@24798.4]
  assign _T_63641 = select_23 == 6'h10; // @[Switch.scala 41:52:@24800.4]
  assign output_16_23 = io_outValid_23 & _T_63641; // @[Switch.scala 41:38:@24801.4]
  assign _T_63644 = select_24 == 6'h10; // @[Switch.scala 41:52:@24803.4]
  assign output_16_24 = io_outValid_24 & _T_63644; // @[Switch.scala 41:38:@24804.4]
  assign _T_63647 = select_25 == 6'h10; // @[Switch.scala 41:52:@24806.4]
  assign output_16_25 = io_outValid_25 & _T_63647; // @[Switch.scala 41:38:@24807.4]
  assign _T_63650 = select_26 == 6'h10; // @[Switch.scala 41:52:@24809.4]
  assign output_16_26 = io_outValid_26 & _T_63650; // @[Switch.scala 41:38:@24810.4]
  assign _T_63653 = select_27 == 6'h10; // @[Switch.scala 41:52:@24812.4]
  assign output_16_27 = io_outValid_27 & _T_63653; // @[Switch.scala 41:38:@24813.4]
  assign _T_63656 = select_28 == 6'h10; // @[Switch.scala 41:52:@24815.4]
  assign output_16_28 = io_outValid_28 & _T_63656; // @[Switch.scala 41:38:@24816.4]
  assign _T_63659 = select_29 == 6'h10; // @[Switch.scala 41:52:@24818.4]
  assign output_16_29 = io_outValid_29 & _T_63659; // @[Switch.scala 41:38:@24819.4]
  assign _T_63662 = select_30 == 6'h10; // @[Switch.scala 41:52:@24821.4]
  assign output_16_30 = io_outValid_30 & _T_63662; // @[Switch.scala 41:38:@24822.4]
  assign _T_63665 = select_31 == 6'h10; // @[Switch.scala 41:52:@24824.4]
  assign output_16_31 = io_outValid_31 & _T_63665; // @[Switch.scala 41:38:@24825.4]
  assign _T_63668 = select_32 == 6'h10; // @[Switch.scala 41:52:@24827.4]
  assign output_16_32 = io_outValid_32 & _T_63668; // @[Switch.scala 41:38:@24828.4]
  assign _T_63671 = select_33 == 6'h10; // @[Switch.scala 41:52:@24830.4]
  assign output_16_33 = io_outValid_33 & _T_63671; // @[Switch.scala 41:38:@24831.4]
  assign _T_63674 = select_34 == 6'h10; // @[Switch.scala 41:52:@24833.4]
  assign output_16_34 = io_outValid_34 & _T_63674; // @[Switch.scala 41:38:@24834.4]
  assign _T_63677 = select_35 == 6'h10; // @[Switch.scala 41:52:@24836.4]
  assign output_16_35 = io_outValid_35 & _T_63677; // @[Switch.scala 41:38:@24837.4]
  assign _T_63680 = select_36 == 6'h10; // @[Switch.scala 41:52:@24839.4]
  assign output_16_36 = io_outValid_36 & _T_63680; // @[Switch.scala 41:38:@24840.4]
  assign _T_63683 = select_37 == 6'h10; // @[Switch.scala 41:52:@24842.4]
  assign output_16_37 = io_outValid_37 & _T_63683; // @[Switch.scala 41:38:@24843.4]
  assign _T_63686 = select_38 == 6'h10; // @[Switch.scala 41:52:@24845.4]
  assign output_16_38 = io_outValid_38 & _T_63686; // @[Switch.scala 41:38:@24846.4]
  assign _T_63689 = select_39 == 6'h10; // @[Switch.scala 41:52:@24848.4]
  assign output_16_39 = io_outValid_39 & _T_63689; // @[Switch.scala 41:38:@24849.4]
  assign _T_63692 = select_40 == 6'h10; // @[Switch.scala 41:52:@24851.4]
  assign output_16_40 = io_outValid_40 & _T_63692; // @[Switch.scala 41:38:@24852.4]
  assign _T_63695 = select_41 == 6'h10; // @[Switch.scala 41:52:@24854.4]
  assign output_16_41 = io_outValid_41 & _T_63695; // @[Switch.scala 41:38:@24855.4]
  assign _T_63698 = select_42 == 6'h10; // @[Switch.scala 41:52:@24857.4]
  assign output_16_42 = io_outValid_42 & _T_63698; // @[Switch.scala 41:38:@24858.4]
  assign _T_63701 = select_43 == 6'h10; // @[Switch.scala 41:52:@24860.4]
  assign output_16_43 = io_outValid_43 & _T_63701; // @[Switch.scala 41:38:@24861.4]
  assign _T_63704 = select_44 == 6'h10; // @[Switch.scala 41:52:@24863.4]
  assign output_16_44 = io_outValid_44 & _T_63704; // @[Switch.scala 41:38:@24864.4]
  assign _T_63707 = select_45 == 6'h10; // @[Switch.scala 41:52:@24866.4]
  assign output_16_45 = io_outValid_45 & _T_63707; // @[Switch.scala 41:38:@24867.4]
  assign _T_63710 = select_46 == 6'h10; // @[Switch.scala 41:52:@24869.4]
  assign output_16_46 = io_outValid_46 & _T_63710; // @[Switch.scala 41:38:@24870.4]
  assign _T_63713 = select_47 == 6'h10; // @[Switch.scala 41:52:@24872.4]
  assign output_16_47 = io_outValid_47 & _T_63713; // @[Switch.scala 41:38:@24873.4]
  assign _T_63716 = select_48 == 6'h10; // @[Switch.scala 41:52:@24875.4]
  assign output_16_48 = io_outValid_48 & _T_63716; // @[Switch.scala 41:38:@24876.4]
  assign _T_63719 = select_49 == 6'h10; // @[Switch.scala 41:52:@24878.4]
  assign output_16_49 = io_outValid_49 & _T_63719; // @[Switch.scala 41:38:@24879.4]
  assign _T_63722 = select_50 == 6'h10; // @[Switch.scala 41:52:@24881.4]
  assign output_16_50 = io_outValid_50 & _T_63722; // @[Switch.scala 41:38:@24882.4]
  assign _T_63725 = select_51 == 6'h10; // @[Switch.scala 41:52:@24884.4]
  assign output_16_51 = io_outValid_51 & _T_63725; // @[Switch.scala 41:38:@24885.4]
  assign _T_63728 = select_52 == 6'h10; // @[Switch.scala 41:52:@24887.4]
  assign output_16_52 = io_outValid_52 & _T_63728; // @[Switch.scala 41:38:@24888.4]
  assign _T_63731 = select_53 == 6'h10; // @[Switch.scala 41:52:@24890.4]
  assign output_16_53 = io_outValid_53 & _T_63731; // @[Switch.scala 41:38:@24891.4]
  assign _T_63734 = select_54 == 6'h10; // @[Switch.scala 41:52:@24893.4]
  assign output_16_54 = io_outValid_54 & _T_63734; // @[Switch.scala 41:38:@24894.4]
  assign _T_63737 = select_55 == 6'h10; // @[Switch.scala 41:52:@24896.4]
  assign output_16_55 = io_outValid_55 & _T_63737; // @[Switch.scala 41:38:@24897.4]
  assign _T_63740 = select_56 == 6'h10; // @[Switch.scala 41:52:@24899.4]
  assign output_16_56 = io_outValid_56 & _T_63740; // @[Switch.scala 41:38:@24900.4]
  assign _T_63743 = select_57 == 6'h10; // @[Switch.scala 41:52:@24902.4]
  assign output_16_57 = io_outValid_57 & _T_63743; // @[Switch.scala 41:38:@24903.4]
  assign _T_63746 = select_58 == 6'h10; // @[Switch.scala 41:52:@24905.4]
  assign output_16_58 = io_outValid_58 & _T_63746; // @[Switch.scala 41:38:@24906.4]
  assign _T_63749 = select_59 == 6'h10; // @[Switch.scala 41:52:@24908.4]
  assign output_16_59 = io_outValid_59 & _T_63749; // @[Switch.scala 41:38:@24909.4]
  assign _T_63752 = select_60 == 6'h10; // @[Switch.scala 41:52:@24911.4]
  assign output_16_60 = io_outValid_60 & _T_63752; // @[Switch.scala 41:38:@24912.4]
  assign _T_63755 = select_61 == 6'h10; // @[Switch.scala 41:52:@24914.4]
  assign output_16_61 = io_outValid_61 & _T_63755; // @[Switch.scala 41:38:@24915.4]
  assign _T_63758 = select_62 == 6'h10; // @[Switch.scala 41:52:@24917.4]
  assign output_16_62 = io_outValid_62 & _T_63758; // @[Switch.scala 41:38:@24918.4]
  assign _T_63761 = select_63 == 6'h10; // @[Switch.scala 41:52:@24920.4]
  assign output_16_63 = io_outValid_63 & _T_63761; // @[Switch.scala 41:38:@24921.4]
  assign _T_63769 = {output_16_7,output_16_6,output_16_5,output_16_4,output_16_3,output_16_2,output_16_1,output_16_0}; // @[Switch.scala 43:31:@24929.4]
  assign _T_63777 = {output_16_15,output_16_14,output_16_13,output_16_12,output_16_11,output_16_10,output_16_9,output_16_8,_T_63769}; // @[Switch.scala 43:31:@24937.4]
  assign _T_63784 = {output_16_23,output_16_22,output_16_21,output_16_20,output_16_19,output_16_18,output_16_17,output_16_16}; // @[Switch.scala 43:31:@24944.4]
  assign _T_63793 = {output_16_31,output_16_30,output_16_29,output_16_28,output_16_27,output_16_26,output_16_25,output_16_24,_T_63784,_T_63777}; // @[Switch.scala 43:31:@24953.4]
  assign _T_63800 = {output_16_39,output_16_38,output_16_37,output_16_36,output_16_35,output_16_34,output_16_33,output_16_32}; // @[Switch.scala 43:31:@24960.4]
  assign _T_63808 = {output_16_47,output_16_46,output_16_45,output_16_44,output_16_43,output_16_42,output_16_41,output_16_40,_T_63800}; // @[Switch.scala 43:31:@24968.4]
  assign _T_63815 = {output_16_55,output_16_54,output_16_53,output_16_52,output_16_51,output_16_50,output_16_49,output_16_48}; // @[Switch.scala 43:31:@24975.4]
  assign _T_63824 = {output_16_63,output_16_62,output_16_61,output_16_60,output_16_59,output_16_58,output_16_57,output_16_56,_T_63815,_T_63808}; // @[Switch.scala 43:31:@24984.4]
  assign _T_63825 = {_T_63824,_T_63793}; // @[Switch.scala 43:31:@24985.4]
  assign _T_63829 = select_0 == 6'h11; // @[Switch.scala 41:52:@24988.4]
  assign output_17_0 = io_outValid_0 & _T_63829; // @[Switch.scala 41:38:@24989.4]
  assign _T_63832 = select_1 == 6'h11; // @[Switch.scala 41:52:@24991.4]
  assign output_17_1 = io_outValid_1 & _T_63832; // @[Switch.scala 41:38:@24992.4]
  assign _T_63835 = select_2 == 6'h11; // @[Switch.scala 41:52:@24994.4]
  assign output_17_2 = io_outValid_2 & _T_63835; // @[Switch.scala 41:38:@24995.4]
  assign _T_63838 = select_3 == 6'h11; // @[Switch.scala 41:52:@24997.4]
  assign output_17_3 = io_outValid_3 & _T_63838; // @[Switch.scala 41:38:@24998.4]
  assign _T_63841 = select_4 == 6'h11; // @[Switch.scala 41:52:@25000.4]
  assign output_17_4 = io_outValid_4 & _T_63841; // @[Switch.scala 41:38:@25001.4]
  assign _T_63844 = select_5 == 6'h11; // @[Switch.scala 41:52:@25003.4]
  assign output_17_5 = io_outValid_5 & _T_63844; // @[Switch.scala 41:38:@25004.4]
  assign _T_63847 = select_6 == 6'h11; // @[Switch.scala 41:52:@25006.4]
  assign output_17_6 = io_outValid_6 & _T_63847; // @[Switch.scala 41:38:@25007.4]
  assign _T_63850 = select_7 == 6'h11; // @[Switch.scala 41:52:@25009.4]
  assign output_17_7 = io_outValid_7 & _T_63850; // @[Switch.scala 41:38:@25010.4]
  assign _T_63853 = select_8 == 6'h11; // @[Switch.scala 41:52:@25012.4]
  assign output_17_8 = io_outValid_8 & _T_63853; // @[Switch.scala 41:38:@25013.4]
  assign _T_63856 = select_9 == 6'h11; // @[Switch.scala 41:52:@25015.4]
  assign output_17_9 = io_outValid_9 & _T_63856; // @[Switch.scala 41:38:@25016.4]
  assign _T_63859 = select_10 == 6'h11; // @[Switch.scala 41:52:@25018.4]
  assign output_17_10 = io_outValid_10 & _T_63859; // @[Switch.scala 41:38:@25019.4]
  assign _T_63862 = select_11 == 6'h11; // @[Switch.scala 41:52:@25021.4]
  assign output_17_11 = io_outValid_11 & _T_63862; // @[Switch.scala 41:38:@25022.4]
  assign _T_63865 = select_12 == 6'h11; // @[Switch.scala 41:52:@25024.4]
  assign output_17_12 = io_outValid_12 & _T_63865; // @[Switch.scala 41:38:@25025.4]
  assign _T_63868 = select_13 == 6'h11; // @[Switch.scala 41:52:@25027.4]
  assign output_17_13 = io_outValid_13 & _T_63868; // @[Switch.scala 41:38:@25028.4]
  assign _T_63871 = select_14 == 6'h11; // @[Switch.scala 41:52:@25030.4]
  assign output_17_14 = io_outValid_14 & _T_63871; // @[Switch.scala 41:38:@25031.4]
  assign _T_63874 = select_15 == 6'h11; // @[Switch.scala 41:52:@25033.4]
  assign output_17_15 = io_outValid_15 & _T_63874; // @[Switch.scala 41:38:@25034.4]
  assign _T_63877 = select_16 == 6'h11; // @[Switch.scala 41:52:@25036.4]
  assign output_17_16 = io_outValid_16 & _T_63877; // @[Switch.scala 41:38:@25037.4]
  assign _T_63880 = select_17 == 6'h11; // @[Switch.scala 41:52:@25039.4]
  assign output_17_17 = io_outValid_17 & _T_63880; // @[Switch.scala 41:38:@25040.4]
  assign _T_63883 = select_18 == 6'h11; // @[Switch.scala 41:52:@25042.4]
  assign output_17_18 = io_outValid_18 & _T_63883; // @[Switch.scala 41:38:@25043.4]
  assign _T_63886 = select_19 == 6'h11; // @[Switch.scala 41:52:@25045.4]
  assign output_17_19 = io_outValid_19 & _T_63886; // @[Switch.scala 41:38:@25046.4]
  assign _T_63889 = select_20 == 6'h11; // @[Switch.scala 41:52:@25048.4]
  assign output_17_20 = io_outValid_20 & _T_63889; // @[Switch.scala 41:38:@25049.4]
  assign _T_63892 = select_21 == 6'h11; // @[Switch.scala 41:52:@25051.4]
  assign output_17_21 = io_outValid_21 & _T_63892; // @[Switch.scala 41:38:@25052.4]
  assign _T_63895 = select_22 == 6'h11; // @[Switch.scala 41:52:@25054.4]
  assign output_17_22 = io_outValid_22 & _T_63895; // @[Switch.scala 41:38:@25055.4]
  assign _T_63898 = select_23 == 6'h11; // @[Switch.scala 41:52:@25057.4]
  assign output_17_23 = io_outValid_23 & _T_63898; // @[Switch.scala 41:38:@25058.4]
  assign _T_63901 = select_24 == 6'h11; // @[Switch.scala 41:52:@25060.4]
  assign output_17_24 = io_outValid_24 & _T_63901; // @[Switch.scala 41:38:@25061.4]
  assign _T_63904 = select_25 == 6'h11; // @[Switch.scala 41:52:@25063.4]
  assign output_17_25 = io_outValid_25 & _T_63904; // @[Switch.scala 41:38:@25064.4]
  assign _T_63907 = select_26 == 6'h11; // @[Switch.scala 41:52:@25066.4]
  assign output_17_26 = io_outValid_26 & _T_63907; // @[Switch.scala 41:38:@25067.4]
  assign _T_63910 = select_27 == 6'h11; // @[Switch.scala 41:52:@25069.4]
  assign output_17_27 = io_outValid_27 & _T_63910; // @[Switch.scala 41:38:@25070.4]
  assign _T_63913 = select_28 == 6'h11; // @[Switch.scala 41:52:@25072.4]
  assign output_17_28 = io_outValid_28 & _T_63913; // @[Switch.scala 41:38:@25073.4]
  assign _T_63916 = select_29 == 6'h11; // @[Switch.scala 41:52:@25075.4]
  assign output_17_29 = io_outValid_29 & _T_63916; // @[Switch.scala 41:38:@25076.4]
  assign _T_63919 = select_30 == 6'h11; // @[Switch.scala 41:52:@25078.4]
  assign output_17_30 = io_outValid_30 & _T_63919; // @[Switch.scala 41:38:@25079.4]
  assign _T_63922 = select_31 == 6'h11; // @[Switch.scala 41:52:@25081.4]
  assign output_17_31 = io_outValid_31 & _T_63922; // @[Switch.scala 41:38:@25082.4]
  assign _T_63925 = select_32 == 6'h11; // @[Switch.scala 41:52:@25084.4]
  assign output_17_32 = io_outValid_32 & _T_63925; // @[Switch.scala 41:38:@25085.4]
  assign _T_63928 = select_33 == 6'h11; // @[Switch.scala 41:52:@25087.4]
  assign output_17_33 = io_outValid_33 & _T_63928; // @[Switch.scala 41:38:@25088.4]
  assign _T_63931 = select_34 == 6'h11; // @[Switch.scala 41:52:@25090.4]
  assign output_17_34 = io_outValid_34 & _T_63931; // @[Switch.scala 41:38:@25091.4]
  assign _T_63934 = select_35 == 6'h11; // @[Switch.scala 41:52:@25093.4]
  assign output_17_35 = io_outValid_35 & _T_63934; // @[Switch.scala 41:38:@25094.4]
  assign _T_63937 = select_36 == 6'h11; // @[Switch.scala 41:52:@25096.4]
  assign output_17_36 = io_outValid_36 & _T_63937; // @[Switch.scala 41:38:@25097.4]
  assign _T_63940 = select_37 == 6'h11; // @[Switch.scala 41:52:@25099.4]
  assign output_17_37 = io_outValid_37 & _T_63940; // @[Switch.scala 41:38:@25100.4]
  assign _T_63943 = select_38 == 6'h11; // @[Switch.scala 41:52:@25102.4]
  assign output_17_38 = io_outValid_38 & _T_63943; // @[Switch.scala 41:38:@25103.4]
  assign _T_63946 = select_39 == 6'h11; // @[Switch.scala 41:52:@25105.4]
  assign output_17_39 = io_outValid_39 & _T_63946; // @[Switch.scala 41:38:@25106.4]
  assign _T_63949 = select_40 == 6'h11; // @[Switch.scala 41:52:@25108.4]
  assign output_17_40 = io_outValid_40 & _T_63949; // @[Switch.scala 41:38:@25109.4]
  assign _T_63952 = select_41 == 6'h11; // @[Switch.scala 41:52:@25111.4]
  assign output_17_41 = io_outValid_41 & _T_63952; // @[Switch.scala 41:38:@25112.4]
  assign _T_63955 = select_42 == 6'h11; // @[Switch.scala 41:52:@25114.4]
  assign output_17_42 = io_outValid_42 & _T_63955; // @[Switch.scala 41:38:@25115.4]
  assign _T_63958 = select_43 == 6'h11; // @[Switch.scala 41:52:@25117.4]
  assign output_17_43 = io_outValid_43 & _T_63958; // @[Switch.scala 41:38:@25118.4]
  assign _T_63961 = select_44 == 6'h11; // @[Switch.scala 41:52:@25120.4]
  assign output_17_44 = io_outValid_44 & _T_63961; // @[Switch.scala 41:38:@25121.4]
  assign _T_63964 = select_45 == 6'h11; // @[Switch.scala 41:52:@25123.4]
  assign output_17_45 = io_outValid_45 & _T_63964; // @[Switch.scala 41:38:@25124.4]
  assign _T_63967 = select_46 == 6'h11; // @[Switch.scala 41:52:@25126.4]
  assign output_17_46 = io_outValid_46 & _T_63967; // @[Switch.scala 41:38:@25127.4]
  assign _T_63970 = select_47 == 6'h11; // @[Switch.scala 41:52:@25129.4]
  assign output_17_47 = io_outValid_47 & _T_63970; // @[Switch.scala 41:38:@25130.4]
  assign _T_63973 = select_48 == 6'h11; // @[Switch.scala 41:52:@25132.4]
  assign output_17_48 = io_outValid_48 & _T_63973; // @[Switch.scala 41:38:@25133.4]
  assign _T_63976 = select_49 == 6'h11; // @[Switch.scala 41:52:@25135.4]
  assign output_17_49 = io_outValid_49 & _T_63976; // @[Switch.scala 41:38:@25136.4]
  assign _T_63979 = select_50 == 6'h11; // @[Switch.scala 41:52:@25138.4]
  assign output_17_50 = io_outValid_50 & _T_63979; // @[Switch.scala 41:38:@25139.4]
  assign _T_63982 = select_51 == 6'h11; // @[Switch.scala 41:52:@25141.4]
  assign output_17_51 = io_outValid_51 & _T_63982; // @[Switch.scala 41:38:@25142.4]
  assign _T_63985 = select_52 == 6'h11; // @[Switch.scala 41:52:@25144.4]
  assign output_17_52 = io_outValid_52 & _T_63985; // @[Switch.scala 41:38:@25145.4]
  assign _T_63988 = select_53 == 6'h11; // @[Switch.scala 41:52:@25147.4]
  assign output_17_53 = io_outValid_53 & _T_63988; // @[Switch.scala 41:38:@25148.4]
  assign _T_63991 = select_54 == 6'h11; // @[Switch.scala 41:52:@25150.4]
  assign output_17_54 = io_outValid_54 & _T_63991; // @[Switch.scala 41:38:@25151.4]
  assign _T_63994 = select_55 == 6'h11; // @[Switch.scala 41:52:@25153.4]
  assign output_17_55 = io_outValid_55 & _T_63994; // @[Switch.scala 41:38:@25154.4]
  assign _T_63997 = select_56 == 6'h11; // @[Switch.scala 41:52:@25156.4]
  assign output_17_56 = io_outValid_56 & _T_63997; // @[Switch.scala 41:38:@25157.4]
  assign _T_64000 = select_57 == 6'h11; // @[Switch.scala 41:52:@25159.4]
  assign output_17_57 = io_outValid_57 & _T_64000; // @[Switch.scala 41:38:@25160.4]
  assign _T_64003 = select_58 == 6'h11; // @[Switch.scala 41:52:@25162.4]
  assign output_17_58 = io_outValid_58 & _T_64003; // @[Switch.scala 41:38:@25163.4]
  assign _T_64006 = select_59 == 6'h11; // @[Switch.scala 41:52:@25165.4]
  assign output_17_59 = io_outValid_59 & _T_64006; // @[Switch.scala 41:38:@25166.4]
  assign _T_64009 = select_60 == 6'h11; // @[Switch.scala 41:52:@25168.4]
  assign output_17_60 = io_outValid_60 & _T_64009; // @[Switch.scala 41:38:@25169.4]
  assign _T_64012 = select_61 == 6'h11; // @[Switch.scala 41:52:@25171.4]
  assign output_17_61 = io_outValid_61 & _T_64012; // @[Switch.scala 41:38:@25172.4]
  assign _T_64015 = select_62 == 6'h11; // @[Switch.scala 41:52:@25174.4]
  assign output_17_62 = io_outValid_62 & _T_64015; // @[Switch.scala 41:38:@25175.4]
  assign _T_64018 = select_63 == 6'h11; // @[Switch.scala 41:52:@25177.4]
  assign output_17_63 = io_outValid_63 & _T_64018; // @[Switch.scala 41:38:@25178.4]
  assign _T_64026 = {output_17_7,output_17_6,output_17_5,output_17_4,output_17_3,output_17_2,output_17_1,output_17_0}; // @[Switch.scala 43:31:@25186.4]
  assign _T_64034 = {output_17_15,output_17_14,output_17_13,output_17_12,output_17_11,output_17_10,output_17_9,output_17_8,_T_64026}; // @[Switch.scala 43:31:@25194.4]
  assign _T_64041 = {output_17_23,output_17_22,output_17_21,output_17_20,output_17_19,output_17_18,output_17_17,output_17_16}; // @[Switch.scala 43:31:@25201.4]
  assign _T_64050 = {output_17_31,output_17_30,output_17_29,output_17_28,output_17_27,output_17_26,output_17_25,output_17_24,_T_64041,_T_64034}; // @[Switch.scala 43:31:@25210.4]
  assign _T_64057 = {output_17_39,output_17_38,output_17_37,output_17_36,output_17_35,output_17_34,output_17_33,output_17_32}; // @[Switch.scala 43:31:@25217.4]
  assign _T_64065 = {output_17_47,output_17_46,output_17_45,output_17_44,output_17_43,output_17_42,output_17_41,output_17_40,_T_64057}; // @[Switch.scala 43:31:@25225.4]
  assign _T_64072 = {output_17_55,output_17_54,output_17_53,output_17_52,output_17_51,output_17_50,output_17_49,output_17_48}; // @[Switch.scala 43:31:@25232.4]
  assign _T_64081 = {output_17_63,output_17_62,output_17_61,output_17_60,output_17_59,output_17_58,output_17_57,output_17_56,_T_64072,_T_64065}; // @[Switch.scala 43:31:@25241.4]
  assign _T_64082 = {_T_64081,_T_64050}; // @[Switch.scala 43:31:@25242.4]
  assign _T_64086 = select_0 == 6'h12; // @[Switch.scala 41:52:@25245.4]
  assign output_18_0 = io_outValid_0 & _T_64086; // @[Switch.scala 41:38:@25246.4]
  assign _T_64089 = select_1 == 6'h12; // @[Switch.scala 41:52:@25248.4]
  assign output_18_1 = io_outValid_1 & _T_64089; // @[Switch.scala 41:38:@25249.4]
  assign _T_64092 = select_2 == 6'h12; // @[Switch.scala 41:52:@25251.4]
  assign output_18_2 = io_outValid_2 & _T_64092; // @[Switch.scala 41:38:@25252.4]
  assign _T_64095 = select_3 == 6'h12; // @[Switch.scala 41:52:@25254.4]
  assign output_18_3 = io_outValid_3 & _T_64095; // @[Switch.scala 41:38:@25255.4]
  assign _T_64098 = select_4 == 6'h12; // @[Switch.scala 41:52:@25257.4]
  assign output_18_4 = io_outValid_4 & _T_64098; // @[Switch.scala 41:38:@25258.4]
  assign _T_64101 = select_5 == 6'h12; // @[Switch.scala 41:52:@25260.4]
  assign output_18_5 = io_outValid_5 & _T_64101; // @[Switch.scala 41:38:@25261.4]
  assign _T_64104 = select_6 == 6'h12; // @[Switch.scala 41:52:@25263.4]
  assign output_18_6 = io_outValid_6 & _T_64104; // @[Switch.scala 41:38:@25264.4]
  assign _T_64107 = select_7 == 6'h12; // @[Switch.scala 41:52:@25266.4]
  assign output_18_7 = io_outValid_7 & _T_64107; // @[Switch.scala 41:38:@25267.4]
  assign _T_64110 = select_8 == 6'h12; // @[Switch.scala 41:52:@25269.4]
  assign output_18_8 = io_outValid_8 & _T_64110; // @[Switch.scala 41:38:@25270.4]
  assign _T_64113 = select_9 == 6'h12; // @[Switch.scala 41:52:@25272.4]
  assign output_18_9 = io_outValid_9 & _T_64113; // @[Switch.scala 41:38:@25273.4]
  assign _T_64116 = select_10 == 6'h12; // @[Switch.scala 41:52:@25275.4]
  assign output_18_10 = io_outValid_10 & _T_64116; // @[Switch.scala 41:38:@25276.4]
  assign _T_64119 = select_11 == 6'h12; // @[Switch.scala 41:52:@25278.4]
  assign output_18_11 = io_outValid_11 & _T_64119; // @[Switch.scala 41:38:@25279.4]
  assign _T_64122 = select_12 == 6'h12; // @[Switch.scala 41:52:@25281.4]
  assign output_18_12 = io_outValid_12 & _T_64122; // @[Switch.scala 41:38:@25282.4]
  assign _T_64125 = select_13 == 6'h12; // @[Switch.scala 41:52:@25284.4]
  assign output_18_13 = io_outValid_13 & _T_64125; // @[Switch.scala 41:38:@25285.4]
  assign _T_64128 = select_14 == 6'h12; // @[Switch.scala 41:52:@25287.4]
  assign output_18_14 = io_outValid_14 & _T_64128; // @[Switch.scala 41:38:@25288.4]
  assign _T_64131 = select_15 == 6'h12; // @[Switch.scala 41:52:@25290.4]
  assign output_18_15 = io_outValid_15 & _T_64131; // @[Switch.scala 41:38:@25291.4]
  assign _T_64134 = select_16 == 6'h12; // @[Switch.scala 41:52:@25293.4]
  assign output_18_16 = io_outValid_16 & _T_64134; // @[Switch.scala 41:38:@25294.4]
  assign _T_64137 = select_17 == 6'h12; // @[Switch.scala 41:52:@25296.4]
  assign output_18_17 = io_outValid_17 & _T_64137; // @[Switch.scala 41:38:@25297.4]
  assign _T_64140 = select_18 == 6'h12; // @[Switch.scala 41:52:@25299.4]
  assign output_18_18 = io_outValid_18 & _T_64140; // @[Switch.scala 41:38:@25300.4]
  assign _T_64143 = select_19 == 6'h12; // @[Switch.scala 41:52:@25302.4]
  assign output_18_19 = io_outValid_19 & _T_64143; // @[Switch.scala 41:38:@25303.4]
  assign _T_64146 = select_20 == 6'h12; // @[Switch.scala 41:52:@25305.4]
  assign output_18_20 = io_outValid_20 & _T_64146; // @[Switch.scala 41:38:@25306.4]
  assign _T_64149 = select_21 == 6'h12; // @[Switch.scala 41:52:@25308.4]
  assign output_18_21 = io_outValid_21 & _T_64149; // @[Switch.scala 41:38:@25309.4]
  assign _T_64152 = select_22 == 6'h12; // @[Switch.scala 41:52:@25311.4]
  assign output_18_22 = io_outValid_22 & _T_64152; // @[Switch.scala 41:38:@25312.4]
  assign _T_64155 = select_23 == 6'h12; // @[Switch.scala 41:52:@25314.4]
  assign output_18_23 = io_outValid_23 & _T_64155; // @[Switch.scala 41:38:@25315.4]
  assign _T_64158 = select_24 == 6'h12; // @[Switch.scala 41:52:@25317.4]
  assign output_18_24 = io_outValid_24 & _T_64158; // @[Switch.scala 41:38:@25318.4]
  assign _T_64161 = select_25 == 6'h12; // @[Switch.scala 41:52:@25320.4]
  assign output_18_25 = io_outValid_25 & _T_64161; // @[Switch.scala 41:38:@25321.4]
  assign _T_64164 = select_26 == 6'h12; // @[Switch.scala 41:52:@25323.4]
  assign output_18_26 = io_outValid_26 & _T_64164; // @[Switch.scala 41:38:@25324.4]
  assign _T_64167 = select_27 == 6'h12; // @[Switch.scala 41:52:@25326.4]
  assign output_18_27 = io_outValid_27 & _T_64167; // @[Switch.scala 41:38:@25327.4]
  assign _T_64170 = select_28 == 6'h12; // @[Switch.scala 41:52:@25329.4]
  assign output_18_28 = io_outValid_28 & _T_64170; // @[Switch.scala 41:38:@25330.4]
  assign _T_64173 = select_29 == 6'h12; // @[Switch.scala 41:52:@25332.4]
  assign output_18_29 = io_outValid_29 & _T_64173; // @[Switch.scala 41:38:@25333.4]
  assign _T_64176 = select_30 == 6'h12; // @[Switch.scala 41:52:@25335.4]
  assign output_18_30 = io_outValid_30 & _T_64176; // @[Switch.scala 41:38:@25336.4]
  assign _T_64179 = select_31 == 6'h12; // @[Switch.scala 41:52:@25338.4]
  assign output_18_31 = io_outValid_31 & _T_64179; // @[Switch.scala 41:38:@25339.4]
  assign _T_64182 = select_32 == 6'h12; // @[Switch.scala 41:52:@25341.4]
  assign output_18_32 = io_outValid_32 & _T_64182; // @[Switch.scala 41:38:@25342.4]
  assign _T_64185 = select_33 == 6'h12; // @[Switch.scala 41:52:@25344.4]
  assign output_18_33 = io_outValid_33 & _T_64185; // @[Switch.scala 41:38:@25345.4]
  assign _T_64188 = select_34 == 6'h12; // @[Switch.scala 41:52:@25347.4]
  assign output_18_34 = io_outValid_34 & _T_64188; // @[Switch.scala 41:38:@25348.4]
  assign _T_64191 = select_35 == 6'h12; // @[Switch.scala 41:52:@25350.4]
  assign output_18_35 = io_outValid_35 & _T_64191; // @[Switch.scala 41:38:@25351.4]
  assign _T_64194 = select_36 == 6'h12; // @[Switch.scala 41:52:@25353.4]
  assign output_18_36 = io_outValid_36 & _T_64194; // @[Switch.scala 41:38:@25354.4]
  assign _T_64197 = select_37 == 6'h12; // @[Switch.scala 41:52:@25356.4]
  assign output_18_37 = io_outValid_37 & _T_64197; // @[Switch.scala 41:38:@25357.4]
  assign _T_64200 = select_38 == 6'h12; // @[Switch.scala 41:52:@25359.4]
  assign output_18_38 = io_outValid_38 & _T_64200; // @[Switch.scala 41:38:@25360.4]
  assign _T_64203 = select_39 == 6'h12; // @[Switch.scala 41:52:@25362.4]
  assign output_18_39 = io_outValid_39 & _T_64203; // @[Switch.scala 41:38:@25363.4]
  assign _T_64206 = select_40 == 6'h12; // @[Switch.scala 41:52:@25365.4]
  assign output_18_40 = io_outValid_40 & _T_64206; // @[Switch.scala 41:38:@25366.4]
  assign _T_64209 = select_41 == 6'h12; // @[Switch.scala 41:52:@25368.4]
  assign output_18_41 = io_outValid_41 & _T_64209; // @[Switch.scala 41:38:@25369.4]
  assign _T_64212 = select_42 == 6'h12; // @[Switch.scala 41:52:@25371.4]
  assign output_18_42 = io_outValid_42 & _T_64212; // @[Switch.scala 41:38:@25372.4]
  assign _T_64215 = select_43 == 6'h12; // @[Switch.scala 41:52:@25374.4]
  assign output_18_43 = io_outValid_43 & _T_64215; // @[Switch.scala 41:38:@25375.4]
  assign _T_64218 = select_44 == 6'h12; // @[Switch.scala 41:52:@25377.4]
  assign output_18_44 = io_outValid_44 & _T_64218; // @[Switch.scala 41:38:@25378.4]
  assign _T_64221 = select_45 == 6'h12; // @[Switch.scala 41:52:@25380.4]
  assign output_18_45 = io_outValid_45 & _T_64221; // @[Switch.scala 41:38:@25381.4]
  assign _T_64224 = select_46 == 6'h12; // @[Switch.scala 41:52:@25383.4]
  assign output_18_46 = io_outValid_46 & _T_64224; // @[Switch.scala 41:38:@25384.4]
  assign _T_64227 = select_47 == 6'h12; // @[Switch.scala 41:52:@25386.4]
  assign output_18_47 = io_outValid_47 & _T_64227; // @[Switch.scala 41:38:@25387.4]
  assign _T_64230 = select_48 == 6'h12; // @[Switch.scala 41:52:@25389.4]
  assign output_18_48 = io_outValid_48 & _T_64230; // @[Switch.scala 41:38:@25390.4]
  assign _T_64233 = select_49 == 6'h12; // @[Switch.scala 41:52:@25392.4]
  assign output_18_49 = io_outValid_49 & _T_64233; // @[Switch.scala 41:38:@25393.4]
  assign _T_64236 = select_50 == 6'h12; // @[Switch.scala 41:52:@25395.4]
  assign output_18_50 = io_outValid_50 & _T_64236; // @[Switch.scala 41:38:@25396.4]
  assign _T_64239 = select_51 == 6'h12; // @[Switch.scala 41:52:@25398.4]
  assign output_18_51 = io_outValid_51 & _T_64239; // @[Switch.scala 41:38:@25399.4]
  assign _T_64242 = select_52 == 6'h12; // @[Switch.scala 41:52:@25401.4]
  assign output_18_52 = io_outValid_52 & _T_64242; // @[Switch.scala 41:38:@25402.4]
  assign _T_64245 = select_53 == 6'h12; // @[Switch.scala 41:52:@25404.4]
  assign output_18_53 = io_outValid_53 & _T_64245; // @[Switch.scala 41:38:@25405.4]
  assign _T_64248 = select_54 == 6'h12; // @[Switch.scala 41:52:@25407.4]
  assign output_18_54 = io_outValid_54 & _T_64248; // @[Switch.scala 41:38:@25408.4]
  assign _T_64251 = select_55 == 6'h12; // @[Switch.scala 41:52:@25410.4]
  assign output_18_55 = io_outValid_55 & _T_64251; // @[Switch.scala 41:38:@25411.4]
  assign _T_64254 = select_56 == 6'h12; // @[Switch.scala 41:52:@25413.4]
  assign output_18_56 = io_outValid_56 & _T_64254; // @[Switch.scala 41:38:@25414.4]
  assign _T_64257 = select_57 == 6'h12; // @[Switch.scala 41:52:@25416.4]
  assign output_18_57 = io_outValid_57 & _T_64257; // @[Switch.scala 41:38:@25417.4]
  assign _T_64260 = select_58 == 6'h12; // @[Switch.scala 41:52:@25419.4]
  assign output_18_58 = io_outValid_58 & _T_64260; // @[Switch.scala 41:38:@25420.4]
  assign _T_64263 = select_59 == 6'h12; // @[Switch.scala 41:52:@25422.4]
  assign output_18_59 = io_outValid_59 & _T_64263; // @[Switch.scala 41:38:@25423.4]
  assign _T_64266 = select_60 == 6'h12; // @[Switch.scala 41:52:@25425.4]
  assign output_18_60 = io_outValid_60 & _T_64266; // @[Switch.scala 41:38:@25426.4]
  assign _T_64269 = select_61 == 6'h12; // @[Switch.scala 41:52:@25428.4]
  assign output_18_61 = io_outValid_61 & _T_64269; // @[Switch.scala 41:38:@25429.4]
  assign _T_64272 = select_62 == 6'h12; // @[Switch.scala 41:52:@25431.4]
  assign output_18_62 = io_outValid_62 & _T_64272; // @[Switch.scala 41:38:@25432.4]
  assign _T_64275 = select_63 == 6'h12; // @[Switch.scala 41:52:@25434.4]
  assign output_18_63 = io_outValid_63 & _T_64275; // @[Switch.scala 41:38:@25435.4]
  assign _T_64283 = {output_18_7,output_18_6,output_18_5,output_18_4,output_18_3,output_18_2,output_18_1,output_18_0}; // @[Switch.scala 43:31:@25443.4]
  assign _T_64291 = {output_18_15,output_18_14,output_18_13,output_18_12,output_18_11,output_18_10,output_18_9,output_18_8,_T_64283}; // @[Switch.scala 43:31:@25451.4]
  assign _T_64298 = {output_18_23,output_18_22,output_18_21,output_18_20,output_18_19,output_18_18,output_18_17,output_18_16}; // @[Switch.scala 43:31:@25458.4]
  assign _T_64307 = {output_18_31,output_18_30,output_18_29,output_18_28,output_18_27,output_18_26,output_18_25,output_18_24,_T_64298,_T_64291}; // @[Switch.scala 43:31:@25467.4]
  assign _T_64314 = {output_18_39,output_18_38,output_18_37,output_18_36,output_18_35,output_18_34,output_18_33,output_18_32}; // @[Switch.scala 43:31:@25474.4]
  assign _T_64322 = {output_18_47,output_18_46,output_18_45,output_18_44,output_18_43,output_18_42,output_18_41,output_18_40,_T_64314}; // @[Switch.scala 43:31:@25482.4]
  assign _T_64329 = {output_18_55,output_18_54,output_18_53,output_18_52,output_18_51,output_18_50,output_18_49,output_18_48}; // @[Switch.scala 43:31:@25489.4]
  assign _T_64338 = {output_18_63,output_18_62,output_18_61,output_18_60,output_18_59,output_18_58,output_18_57,output_18_56,_T_64329,_T_64322}; // @[Switch.scala 43:31:@25498.4]
  assign _T_64339 = {_T_64338,_T_64307}; // @[Switch.scala 43:31:@25499.4]
  assign _T_64343 = select_0 == 6'h13; // @[Switch.scala 41:52:@25502.4]
  assign output_19_0 = io_outValid_0 & _T_64343; // @[Switch.scala 41:38:@25503.4]
  assign _T_64346 = select_1 == 6'h13; // @[Switch.scala 41:52:@25505.4]
  assign output_19_1 = io_outValid_1 & _T_64346; // @[Switch.scala 41:38:@25506.4]
  assign _T_64349 = select_2 == 6'h13; // @[Switch.scala 41:52:@25508.4]
  assign output_19_2 = io_outValid_2 & _T_64349; // @[Switch.scala 41:38:@25509.4]
  assign _T_64352 = select_3 == 6'h13; // @[Switch.scala 41:52:@25511.4]
  assign output_19_3 = io_outValid_3 & _T_64352; // @[Switch.scala 41:38:@25512.4]
  assign _T_64355 = select_4 == 6'h13; // @[Switch.scala 41:52:@25514.4]
  assign output_19_4 = io_outValid_4 & _T_64355; // @[Switch.scala 41:38:@25515.4]
  assign _T_64358 = select_5 == 6'h13; // @[Switch.scala 41:52:@25517.4]
  assign output_19_5 = io_outValid_5 & _T_64358; // @[Switch.scala 41:38:@25518.4]
  assign _T_64361 = select_6 == 6'h13; // @[Switch.scala 41:52:@25520.4]
  assign output_19_6 = io_outValid_6 & _T_64361; // @[Switch.scala 41:38:@25521.4]
  assign _T_64364 = select_7 == 6'h13; // @[Switch.scala 41:52:@25523.4]
  assign output_19_7 = io_outValid_7 & _T_64364; // @[Switch.scala 41:38:@25524.4]
  assign _T_64367 = select_8 == 6'h13; // @[Switch.scala 41:52:@25526.4]
  assign output_19_8 = io_outValid_8 & _T_64367; // @[Switch.scala 41:38:@25527.4]
  assign _T_64370 = select_9 == 6'h13; // @[Switch.scala 41:52:@25529.4]
  assign output_19_9 = io_outValid_9 & _T_64370; // @[Switch.scala 41:38:@25530.4]
  assign _T_64373 = select_10 == 6'h13; // @[Switch.scala 41:52:@25532.4]
  assign output_19_10 = io_outValid_10 & _T_64373; // @[Switch.scala 41:38:@25533.4]
  assign _T_64376 = select_11 == 6'h13; // @[Switch.scala 41:52:@25535.4]
  assign output_19_11 = io_outValid_11 & _T_64376; // @[Switch.scala 41:38:@25536.4]
  assign _T_64379 = select_12 == 6'h13; // @[Switch.scala 41:52:@25538.4]
  assign output_19_12 = io_outValid_12 & _T_64379; // @[Switch.scala 41:38:@25539.4]
  assign _T_64382 = select_13 == 6'h13; // @[Switch.scala 41:52:@25541.4]
  assign output_19_13 = io_outValid_13 & _T_64382; // @[Switch.scala 41:38:@25542.4]
  assign _T_64385 = select_14 == 6'h13; // @[Switch.scala 41:52:@25544.4]
  assign output_19_14 = io_outValid_14 & _T_64385; // @[Switch.scala 41:38:@25545.4]
  assign _T_64388 = select_15 == 6'h13; // @[Switch.scala 41:52:@25547.4]
  assign output_19_15 = io_outValid_15 & _T_64388; // @[Switch.scala 41:38:@25548.4]
  assign _T_64391 = select_16 == 6'h13; // @[Switch.scala 41:52:@25550.4]
  assign output_19_16 = io_outValid_16 & _T_64391; // @[Switch.scala 41:38:@25551.4]
  assign _T_64394 = select_17 == 6'h13; // @[Switch.scala 41:52:@25553.4]
  assign output_19_17 = io_outValid_17 & _T_64394; // @[Switch.scala 41:38:@25554.4]
  assign _T_64397 = select_18 == 6'h13; // @[Switch.scala 41:52:@25556.4]
  assign output_19_18 = io_outValid_18 & _T_64397; // @[Switch.scala 41:38:@25557.4]
  assign _T_64400 = select_19 == 6'h13; // @[Switch.scala 41:52:@25559.4]
  assign output_19_19 = io_outValid_19 & _T_64400; // @[Switch.scala 41:38:@25560.4]
  assign _T_64403 = select_20 == 6'h13; // @[Switch.scala 41:52:@25562.4]
  assign output_19_20 = io_outValid_20 & _T_64403; // @[Switch.scala 41:38:@25563.4]
  assign _T_64406 = select_21 == 6'h13; // @[Switch.scala 41:52:@25565.4]
  assign output_19_21 = io_outValid_21 & _T_64406; // @[Switch.scala 41:38:@25566.4]
  assign _T_64409 = select_22 == 6'h13; // @[Switch.scala 41:52:@25568.4]
  assign output_19_22 = io_outValid_22 & _T_64409; // @[Switch.scala 41:38:@25569.4]
  assign _T_64412 = select_23 == 6'h13; // @[Switch.scala 41:52:@25571.4]
  assign output_19_23 = io_outValid_23 & _T_64412; // @[Switch.scala 41:38:@25572.4]
  assign _T_64415 = select_24 == 6'h13; // @[Switch.scala 41:52:@25574.4]
  assign output_19_24 = io_outValid_24 & _T_64415; // @[Switch.scala 41:38:@25575.4]
  assign _T_64418 = select_25 == 6'h13; // @[Switch.scala 41:52:@25577.4]
  assign output_19_25 = io_outValid_25 & _T_64418; // @[Switch.scala 41:38:@25578.4]
  assign _T_64421 = select_26 == 6'h13; // @[Switch.scala 41:52:@25580.4]
  assign output_19_26 = io_outValid_26 & _T_64421; // @[Switch.scala 41:38:@25581.4]
  assign _T_64424 = select_27 == 6'h13; // @[Switch.scala 41:52:@25583.4]
  assign output_19_27 = io_outValid_27 & _T_64424; // @[Switch.scala 41:38:@25584.4]
  assign _T_64427 = select_28 == 6'h13; // @[Switch.scala 41:52:@25586.4]
  assign output_19_28 = io_outValid_28 & _T_64427; // @[Switch.scala 41:38:@25587.4]
  assign _T_64430 = select_29 == 6'h13; // @[Switch.scala 41:52:@25589.4]
  assign output_19_29 = io_outValid_29 & _T_64430; // @[Switch.scala 41:38:@25590.4]
  assign _T_64433 = select_30 == 6'h13; // @[Switch.scala 41:52:@25592.4]
  assign output_19_30 = io_outValid_30 & _T_64433; // @[Switch.scala 41:38:@25593.4]
  assign _T_64436 = select_31 == 6'h13; // @[Switch.scala 41:52:@25595.4]
  assign output_19_31 = io_outValid_31 & _T_64436; // @[Switch.scala 41:38:@25596.4]
  assign _T_64439 = select_32 == 6'h13; // @[Switch.scala 41:52:@25598.4]
  assign output_19_32 = io_outValid_32 & _T_64439; // @[Switch.scala 41:38:@25599.4]
  assign _T_64442 = select_33 == 6'h13; // @[Switch.scala 41:52:@25601.4]
  assign output_19_33 = io_outValid_33 & _T_64442; // @[Switch.scala 41:38:@25602.4]
  assign _T_64445 = select_34 == 6'h13; // @[Switch.scala 41:52:@25604.4]
  assign output_19_34 = io_outValid_34 & _T_64445; // @[Switch.scala 41:38:@25605.4]
  assign _T_64448 = select_35 == 6'h13; // @[Switch.scala 41:52:@25607.4]
  assign output_19_35 = io_outValid_35 & _T_64448; // @[Switch.scala 41:38:@25608.4]
  assign _T_64451 = select_36 == 6'h13; // @[Switch.scala 41:52:@25610.4]
  assign output_19_36 = io_outValid_36 & _T_64451; // @[Switch.scala 41:38:@25611.4]
  assign _T_64454 = select_37 == 6'h13; // @[Switch.scala 41:52:@25613.4]
  assign output_19_37 = io_outValid_37 & _T_64454; // @[Switch.scala 41:38:@25614.4]
  assign _T_64457 = select_38 == 6'h13; // @[Switch.scala 41:52:@25616.4]
  assign output_19_38 = io_outValid_38 & _T_64457; // @[Switch.scala 41:38:@25617.4]
  assign _T_64460 = select_39 == 6'h13; // @[Switch.scala 41:52:@25619.4]
  assign output_19_39 = io_outValid_39 & _T_64460; // @[Switch.scala 41:38:@25620.4]
  assign _T_64463 = select_40 == 6'h13; // @[Switch.scala 41:52:@25622.4]
  assign output_19_40 = io_outValid_40 & _T_64463; // @[Switch.scala 41:38:@25623.4]
  assign _T_64466 = select_41 == 6'h13; // @[Switch.scala 41:52:@25625.4]
  assign output_19_41 = io_outValid_41 & _T_64466; // @[Switch.scala 41:38:@25626.4]
  assign _T_64469 = select_42 == 6'h13; // @[Switch.scala 41:52:@25628.4]
  assign output_19_42 = io_outValid_42 & _T_64469; // @[Switch.scala 41:38:@25629.4]
  assign _T_64472 = select_43 == 6'h13; // @[Switch.scala 41:52:@25631.4]
  assign output_19_43 = io_outValid_43 & _T_64472; // @[Switch.scala 41:38:@25632.4]
  assign _T_64475 = select_44 == 6'h13; // @[Switch.scala 41:52:@25634.4]
  assign output_19_44 = io_outValid_44 & _T_64475; // @[Switch.scala 41:38:@25635.4]
  assign _T_64478 = select_45 == 6'h13; // @[Switch.scala 41:52:@25637.4]
  assign output_19_45 = io_outValid_45 & _T_64478; // @[Switch.scala 41:38:@25638.4]
  assign _T_64481 = select_46 == 6'h13; // @[Switch.scala 41:52:@25640.4]
  assign output_19_46 = io_outValid_46 & _T_64481; // @[Switch.scala 41:38:@25641.4]
  assign _T_64484 = select_47 == 6'h13; // @[Switch.scala 41:52:@25643.4]
  assign output_19_47 = io_outValid_47 & _T_64484; // @[Switch.scala 41:38:@25644.4]
  assign _T_64487 = select_48 == 6'h13; // @[Switch.scala 41:52:@25646.4]
  assign output_19_48 = io_outValid_48 & _T_64487; // @[Switch.scala 41:38:@25647.4]
  assign _T_64490 = select_49 == 6'h13; // @[Switch.scala 41:52:@25649.4]
  assign output_19_49 = io_outValid_49 & _T_64490; // @[Switch.scala 41:38:@25650.4]
  assign _T_64493 = select_50 == 6'h13; // @[Switch.scala 41:52:@25652.4]
  assign output_19_50 = io_outValid_50 & _T_64493; // @[Switch.scala 41:38:@25653.4]
  assign _T_64496 = select_51 == 6'h13; // @[Switch.scala 41:52:@25655.4]
  assign output_19_51 = io_outValid_51 & _T_64496; // @[Switch.scala 41:38:@25656.4]
  assign _T_64499 = select_52 == 6'h13; // @[Switch.scala 41:52:@25658.4]
  assign output_19_52 = io_outValid_52 & _T_64499; // @[Switch.scala 41:38:@25659.4]
  assign _T_64502 = select_53 == 6'h13; // @[Switch.scala 41:52:@25661.4]
  assign output_19_53 = io_outValid_53 & _T_64502; // @[Switch.scala 41:38:@25662.4]
  assign _T_64505 = select_54 == 6'h13; // @[Switch.scala 41:52:@25664.4]
  assign output_19_54 = io_outValid_54 & _T_64505; // @[Switch.scala 41:38:@25665.4]
  assign _T_64508 = select_55 == 6'h13; // @[Switch.scala 41:52:@25667.4]
  assign output_19_55 = io_outValid_55 & _T_64508; // @[Switch.scala 41:38:@25668.4]
  assign _T_64511 = select_56 == 6'h13; // @[Switch.scala 41:52:@25670.4]
  assign output_19_56 = io_outValid_56 & _T_64511; // @[Switch.scala 41:38:@25671.4]
  assign _T_64514 = select_57 == 6'h13; // @[Switch.scala 41:52:@25673.4]
  assign output_19_57 = io_outValid_57 & _T_64514; // @[Switch.scala 41:38:@25674.4]
  assign _T_64517 = select_58 == 6'h13; // @[Switch.scala 41:52:@25676.4]
  assign output_19_58 = io_outValid_58 & _T_64517; // @[Switch.scala 41:38:@25677.4]
  assign _T_64520 = select_59 == 6'h13; // @[Switch.scala 41:52:@25679.4]
  assign output_19_59 = io_outValid_59 & _T_64520; // @[Switch.scala 41:38:@25680.4]
  assign _T_64523 = select_60 == 6'h13; // @[Switch.scala 41:52:@25682.4]
  assign output_19_60 = io_outValid_60 & _T_64523; // @[Switch.scala 41:38:@25683.4]
  assign _T_64526 = select_61 == 6'h13; // @[Switch.scala 41:52:@25685.4]
  assign output_19_61 = io_outValid_61 & _T_64526; // @[Switch.scala 41:38:@25686.4]
  assign _T_64529 = select_62 == 6'h13; // @[Switch.scala 41:52:@25688.4]
  assign output_19_62 = io_outValid_62 & _T_64529; // @[Switch.scala 41:38:@25689.4]
  assign _T_64532 = select_63 == 6'h13; // @[Switch.scala 41:52:@25691.4]
  assign output_19_63 = io_outValid_63 & _T_64532; // @[Switch.scala 41:38:@25692.4]
  assign _T_64540 = {output_19_7,output_19_6,output_19_5,output_19_4,output_19_3,output_19_2,output_19_1,output_19_0}; // @[Switch.scala 43:31:@25700.4]
  assign _T_64548 = {output_19_15,output_19_14,output_19_13,output_19_12,output_19_11,output_19_10,output_19_9,output_19_8,_T_64540}; // @[Switch.scala 43:31:@25708.4]
  assign _T_64555 = {output_19_23,output_19_22,output_19_21,output_19_20,output_19_19,output_19_18,output_19_17,output_19_16}; // @[Switch.scala 43:31:@25715.4]
  assign _T_64564 = {output_19_31,output_19_30,output_19_29,output_19_28,output_19_27,output_19_26,output_19_25,output_19_24,_T_64555,_T_64548}; // @[Switch.scala 43:31:@25724.4]
  assign _T_64571 = {output_19_39,output_19_38,output_19_37,output_19_36,output_19_35,output_19_34,output_19_33,output_19_32}; // @[Switch.scala 43:31:@25731.4]
  assign _T_64579 = {output_19_47,output_19_46,output_19_45,output_19_44,output_19_43,output_19_42,output_19_41,output_19_40,_T_64571}; // @[Switch.scala 43:31:@25739.4]
  assign _T_64586 = {output_19_55,output_19_54,output_19_53,output_19_52,output_19_51,output_19_50,output_19_49,output_19_48}; // @[Switch.scala 43:31:@25746.4]
  assign _T_64595 = {output_19_63,output_19_62,output_19_61,output_19_60,output_19_59,output_19_58,output_19_57,output_19_56,_T_64586,_T_64579}; // @[Switch.scala 43:31:@25755.4]
  assign _T_64596 = {_T_64595,_T_64564}; // @[Switch.scala 43:31:@25756.4]
  assign _T_64600 = select_0 == 6'h14; // @[Switch.scala 41:52:@25759.4]
  assign output_20_0 = io_outValid_0 & _T_64600; // @[Switch.scala 41:38:@25760.4]
  assign _T_64603 = select_1 == 6'h14; // @[Switch.scala 41:52:@25762.4]
  assign output_20_1 = io_outValid_1 & _T_64603; // @[Switch.scala 41:38:@25763.4]
  assign _T_64606 = select_2 == 6'h14; // @[Switch.scala 41:52:@25765.4]
  assign output_20_2 = io_outValid_2 & _T_64606; // @[Switch.scala 41:38:@25766.4]
  assign _T_64609 = select_3 == 6'h14; // @[Switch.scala 41:52:@25768.4]
  assign output_20_3 = io_outValid_3 & _T_64609; // @[Switch.scala 41:38:@25769.4]
  assign _T_64612 = select_4 == 6'h14; // @[Switch.scala 41:52:@25771.4]
  assign output_20_4 = io_outValid_4 & _T_64612; // @[Switch.scala 41:38:@25772.4]
  assign _T_64615 = select_5 == 6'h14; // @[Switch.scala 41:52:@25774.4]
  assign output_20_5 = io_outValid_5 & _T_64615; // @[Switch.scala 41:38:@25775.4]
  assign _T_64618 = select_6 == 6'h14; // @[Switch.scala 41:52:@25777.4]
  assign output_20_6 = io_outValid_6 & _T_64618; // @[Switch.scala 41:38:@25778.4]
  assign _T_64621 = select_7 == 6'h14; // @[Switch.scala 41:52:@25780.4]
  assign output_20_7 = io_outValid_7 & _T_64621; // @[Switch.scala 41:38:@25781.4]
  assign _T_64624 = select_8 == 6'h14; // @[Switch.scala 41:52:@25783.4]
  assign output_20_8 = io_outValid_8 & _T_64624; // @[Switch.scala 41:38:@25784.4]
  assign _T_64627 = select_9 == 6'h14; // @[Switch.scala 41:52:@25786.4]
  assign output_20_9 = io_outValid_9 & _T_64627; // @[Switch.scala 41:38:@25787.4]
  assign _T_64630 = select_10 == 6'h14; // @[Switch.scala 41:52:@25789.4]
  assign output_20_10 = io_outValid_10 & _T_64630; // @[Switch.scala 41:38:@25790.4]
  assign _T_64633 = select_11 == 6'h14; // @[Switch.scala 41:52:@25792.4]
  assign output_20_11 = io_outValid_11 & _T_64633; // @[Switch.scala 41:38:@25793.4]
  assign _T_64636 = select_12 == 6'h14; // @[Switch.scala 41:52:@25795.4]
  assign output_20_12 = io_outValid_12 & _T_64636; // @[Switch.scala 41:38:@25796.4]
  assign _T_64639 = select_13 == 6'h14; // @[Switch.scala 41:52:@25798.4]
  assign output_20_13 = io_outValid_13 & _T_64639; // @[Switch.scala 41:38:@25799.4]
  assign _T_64642 = select_14 == 6'h14; // @[Switch.scala 41:52:@25801.4]
  assign output_20_14 = io_outValid_14 & _T_64642; // @[Switch.scala 41:38:@25802.4]
  assign _T_64645 = select_15 == 6'h14; // @[Switch.scala 41:52:@25804.4]
  assign output_20_15 = io_outValid_15 & _T_64645; // @[Switch.scala 41:38:@25805.4]
  assign _T_64648 = select_16 == 6'h14; // @[Switch.scala 41:52:@25807.4]
  assign output_20_16 = io_outValid_16 & _T_64648; // @[Switch.scala 41:38:@25808.4]
  assign _T_64651 = select_17 == 6'h14; // @[Switch.scala 41:52:@25810.4]
  assign output_20_17 = io_outValid_17 & _T_64651; // @[Switch.scala 41:38:@25811.4]
  assign _T_64654 = select_18 == 6'h14; // @[Switch.scala 41:52:@25813.4]
  assign output_20_18 = io_outValid_18 & _T_64654; // @[Switch.scala 41:38:@25814.4]
  assign _T_64657 = select_19 == 6'h14; // @[Switch.scala 41:52:@25816.4]
  assign output_20_19 = io_outValid_19 & _T_64657; // @[Switch.scala 41:38:@25817.4]
  assign _T_64660 = select_20 == 6'h14; // @[Switch.scala 41:52:@25819.4]
  assign output_20_20 = io_outValid_20 & _T_64660; // @[Switch.scala 41:38:@25820.4]
  assign _T_64663 = select_21 == 6'h14; // @[Switch.scala 41:52:@25822.4]
  assign output_20_21 = io_outValid_21 & _T_64663; // @[Switch.scala 41:38:@25823.4]
  assign _T_64666 = select_22 == 6'h14; // @[Switch.scala 41:52:@25825.4]
  assign output_20_22 = io_outValid_22 & _T_64666; // @[Switch.scala 41:38:@25826.4]
  assign _T_64669 = select_23 == 6'h14; // @[Switch.scala 41:52:@25828.4]
  assign output_20_23 = io_outValid_23 & _T_64669; // @[Switch.scala 41:38:@25829.4]
  assign _T_64672 = select_24 == 6'h14; // @[Switch.scala 41:52:@25831.4]
  assign output_20_24 = io_outValid_24 & _T_64672; // @[Switch.scala 41:38:@25832.4]
  assign _T_64675 = select_25 == 6'h14; // @[Switch.scala 41:52:@25834.4]
  assign output_20_25 = io_outValid_25 & _T_64675; // @[Switch.scala 41:38:@25835.4]
  assign _T_64678 = select_26 == 6'h14; // @[Switch.scala 41:52:@25837.4]
  assign output_20_26 = io_outValid_26 & _T_64678; // @[Switch.scala 41:38:@25838.4]
  assign _T_64681 = select_27 == 6'h14; // @[Switch.scala 41:52:@25840.4]
  assign output_20_27 = io_outValid_27 & _T_64681; // @[Switch.scala 41:38:@25841.4]
  assign _T_64684 = select_28 == 6'h14; // @[Switch.scala 41:52:@25843.4]
  assign output_20_28 = io_outValid_28 & _T_64684; // @[Switch.scala 41:38:@25844.4]
  assign _T_64687 = select_29 == 6'h14; // @[Switch.scala 41:52:@25846.4]
  assign output_20_29 = io_outValid_29 & _T_64687; // @[Switch.scala 41:38:@25847.4]
  assign _T_64690 = select_30 == 6'h14; // @[Switch.scala 41:52:@25849.4]
  assign output_20_30 = io_outValid_30 & _T_64690; // @[Switch.scala 41:38:@25850.4]
  assign _T_64693 = select_31 == 6'h14; // @[Switch.scala 41:52:@25852.4]
  assign output_20_31 = io_outValid_31 & _T_64693; // @[Switch.scala 41:38:@25853.4]
  assign _T_64696 = select_32 == 6'h14; // @[Switch.scala 41:52:@25855.4]
  assign output_20_32 = io_outValid_32 & _T_64696; // @[Switch.scala 41:38:@25856.4]
  assign _T_64699 = select_33 == 6'h14; // @[Switch.scala 41:52:@25858.4]
  assign output_20_33 = io_outValid_33 & _T_64699; // @[Switch.scala 41:38:@25859.4]
  assign _T_64702 = select_34 == 6'h14; // @[Switch.scala 41:52:@25861.4]
  assign output_20_34 = io_outValid_34 & _T_64702; // @[Switch.scala 41:38:@25862.4]
  assign _T_64705 = select_35 == 6'h14; // @[Switch.scala 41:52:@25864.4]
  assign output_20_35 = io_outValid_35 & _T_64705; // @[Switch.scala 41:38:@25865.4]
  assign _T_64708 = select_36 == 6'h14; // @[Switch.scala 41:52:@25867.4]
  assign output_20_36 = io_outValid_36 & _T_64708; // @[Switch.scala 41:38:@25868.4]
  assign _T_64711 = select_37 == 6'h14; // @[Switch.scala 41:52:@25870.4]
  assign output_20_37 = io_outValid_37 & _T_64711; // @[Switch.scala 41:38:@25871.4]
  assign _T_64714 = select_38 == 6'h14; // @[Switch.scala 41:52:@25873.4]
  assign output_20_38 = io_outValid_38 & _T_64714; // @[Switch.scala 41:38:@25874.4]
  assign _T_64717 = select_39 == 6'h14; // @[Switch.scala 41:52:@25876.4]
  assign output_20_39 = io_outValid_39 & _T_64717; // @[Switch.scala 41:38:@25877.4]
  assign _T_64720 = select_40 == 6'h14; // @[Switch.scala 41:52:@25879.4]
  assign output_20_40 = io_outValid_40 & _T_64720; // @[Switch.scala 41:38:@25880.4]
  assign _T_64723 = select_41 == 6'h14; // @[Switch.scala 41:52:@25882.4]
  assign output_20_41 = io_outValid_41 & _T_64723; // @[Switch.scala 41:38:@25883.4]
  assign _T_64726 = select_42 == 6'h14; // @[Switch.scala 41:52:@25885.4]
  assign output_20_42 = io_outValid_42 & _T_64726; // @[Switch.scala 41:38:@25886.4]
  assign _T_64729 = select_43 == 6'h14; // @[Switch.scala 41:52:@25888.4]
  assign output_20_43 = io_outValid_43 & _T_64729; // @[Switch.scala 41:38:@25889.4]
  assign _T_64732 = select_44 == 6'h14; // @[Switch.scala 41:52:@25891.4]
  assign output_20_44 = io_outValid_44 & _T_64732; // @[Switch.scala 41:38:@25892.4]
  assign _T_64735 = select_45 == 6'h14; // @[Switch.scala 41:52:@25894.4]
  assign output_20_45 = io_outValid_45 & _T_64735; // @[Switch.scala 41:38:@25895.4]
  assign _T_64738 = select_46 == 6'h14; // @[Switch.scala 41:52:@25897.4]
  assign output_20_46 = io_outValid_46 & _T_64738; // @[Switch.scala 41:38:@25898.4]
  assign _T_64741 = select_47 == 6'h14; // @[Switch.scala 41:52:@25900.4]
  assign output_20_47 = io_outValid_47 & _T_64741; // @[Switch.scala 41:38:@25901.4]
  assign _T_64744 = select_48 == 6'h14; // @[Switch.scala 41:52:@25903.4]
  assign output_20_48 = io_outValid_48 & _T_64744; // @[Switch.scala 41:38:@25904.4]
  assign _T_64747 = select_49 == 6'h14; // @[Switch.scala 41:52:@25906.4]
  assign output_20_49 = io_outValid_49 & _T_64747; // @[Switch.scala 41:38:@25907.4]
  assign _T_64750 = select_50 == 6'h14; // @[Switch.scala 41:52:@25909.4]
  assign output_20_50 = io_outValid_50 & _T_64750; // @[Switch.scala 41:38:@25910.4]
  assign _T_64753 = select_51 == 6'h14; // @[Switch.scala 41:52:@25912.4]
  assign output_20_51 = io_outValid_51 & _T_64753; // @[Switch.scala 41:38:@25913.4]
  assign _T_64756 = select_52 == 6'h14; // @[Switch.scala 41:52:@25915.4]
  assign output_20_52 = io_outValid_52 & _T_64756; // @[Switch.scala 41:38:@25916.4]
  assign _T_64759 = select_53 == 6'h14; // @[Switch.scala 41:52:@25918.4]
  assign output_20_53 = io_outValid_53 & _T_64759; // @[Switch.scala 41:38:@25919.4]
  assign _T_64762 = select_54 == 6'h14; // @[Switch.scala 41:52:@25921.4]
  assign output_20_54 = io_outValid_54 & _T_64762; // @[Switch.scala 41:38:@25922.4]
  assign _T_64765 = select_55 == 6'h14; // @[Switch.scala 41:52:@25924.4]
  assign output_20_55 = io_outValid_55 & _T_64765; // @[Switch.scala 41:38:@25925.4]
  assign _T_64768 = select_56 == 6'h14; // @[Switch.scala 41:52:@25927.4]
  assign output_20_56 = io_outValid_56 & _T_64768; // @[Switch.scala 41:38:@25928.4]
  assign _T_64771 = select_57 == 6'h14; // @[Switch.scala 41:52:@25930.4]
  assign output_20_57 = io_outValid_57 & _T_64771; // @[Switch.scala 41:38:@25931.4]
  assign _T_64774 = select_58 == 6'h14; // @[Switch.scala 41:52:@25933.4]
  assign output_20_58 = io_outValid_58 & _T_64774; // @[Switch.scala 41:38:@25934.4]
  assign _T_64777 = select_59 == 6'h14; // @[Switch.scala 41:52:@25936.4]
  assign output_20_59 = io_outValid_59 & _T_64777; // @[Switch.scala 41:38:@25937.4]
  assign _T_64780 = select_60 == 6'h14; // @[Switch.scala 41:52:@25939.4]
  assign output_20_60 = io_outValid_60 & _T_64780; // @[Switch.scala 41:38:@25940.4]
  assign _T_64783 = select_61 == 6'h14; // @[Switch.scala 41:52:@25942.4]
  assign output_20_61 = io_outValid_61 & _T_64783; // @[Switch.scala 41:38:@25943.4]
  assign _T_64786 = select_62 == 6'h14; // @[Switch.scala 41:52:@25945.4]
  assign output_20_62 = io_outValid_62 & _T_64786; // @[Switch.scala 41:38:@25946.4]
  assign _T_64789 = select_63 == 6'h14; // @[Switch.scala 41:52:@25948.4]
  assign output_20_63 = io_outValid_63 & _T_64789; // @[Switch.scala 41:38:@25949.4]
  assign _T_64797 = {output_20_7,output_20_6,output_20_5,output_20_4,output_20_3,output_20_2,output_20_1,output_20_0}; // @[Switch.scala 43:31:@25957.4]
  assign _T_64805 = {output_20_15,output_20_14,output_20_13,output_20_12,output_20_11,output_20_10,output_20_9,output_20_8,_T_64797}; // @[Switch.scala 43:31:@25965.4]
  assign _T_64812 = {output_20_23,output_20_22,output_20_21,output_20_20,output_20_19,output_20_18,output_20_17,output_20_16}; // @[Switch.scala 43:31:@25972.4]
  assign _T_64821 = {output_20_31,output_20_30,output_20_29,output_20_28,output_20_27,output_20_26,output_20_25,output_20_24,_T_64812,_T_64805}; // @[Switch.scala 43:31:@25981.4]
  assign _T_64828 = {output_20_39,output_20_38,output_20_37,output_20_36,output_20_35,output_20_34,output_20_33,output_20_32}; // @[Switch.scala 43:31:@25988.4]
  assign _T_64836 = {output_20_47,output_20_46,output_20_45,output_20_44,output_20_43,output_20_42,output_20_41,output_20_40,_T_64828}; // @[Switch.scala 43:31:@25996.4]
  assign _T_64843 = {output_20_55,output_20_54,output_20_53,output_20_52,output_20_51,output_20_50,output_20_49,output_20_48}; // @[Switch.scala 43:31:@26003.4]
  assign _T_64852 = {output_20_63,output_20_62,output_20_61,output_20_60,output_20_59,output_20_58,output_20_57,output_20_56,_T_64843,_T_64836}; // @[Switch.scala 43:31:@26012.4]
  assign _T_64853 = {_T_64852,_T_64821}; // @[Switch.scala 43:31:@26013.4]
  assign _T_64857 = select_0 == 6'h15; // @[Switch.scala 41:52:@26016.4]
  assign output_21_0 = io_outValid_0 & _T_64857; // @[Switch.scala 41:38:@26017.4]
  assign _T_64860 = select_1 == 6'h15; // @[Switch.scala 41:52:@26019.4]
  assign output_21_1 = io_outValid_1 & _T_64860; // @[Switch.scala 41:38:@26020.4]
  assign _T_64863 = select_2 == 6'h15; // @[Switch.scala 41:52:@26022.4]
  assign output_21_2 = io_outValid_2 & _T_64863; // @[Switch.scala 41:38:@26023.4]
  assign _T_64866 = select_3 == 6'h15; // @[Switch.scala 41:52:@26025.4]
  assign output_21_3 = io_outValid_3 & _T_64866; // @[Switch.scala 41:38:@26026.4]
  assign _T_64869 = select_4 == 6'h15; // @[Switch.scala 41:52:@26028.4]
  assign output_21_4 = io_outValid_4 & _T_64869; // @[Switch.scala 41:38:@26029.4]
  assign _T_64872 = select_5 == 6'h15; // @[Switch.scala 41:52:@26031.4]
  assign output_21_5 = io_outValid_5 & _T_64872; // @[Switch.scala 41:38:@26032.4]
  assign _T_64875 = select_6 == 6'h15; // @[Switch.scala 41:52:@26034.4]
  assign output_21_6 = io_outValid_6 & _T_64875; // @[Switch.scala 41:38:@26035.4]
  assign _T_64878 = select_7 == 6'h15; // @[Switch.scala 41:52:@26037.4]
  assign output_21_7 = io_outValid_7 & _T_64878; // @[Switch.scala 41:38:@26038.4]
  assign _T_64881 = select_8 == 6'h15; // @[Switch.scala 41:52:@26040.4]
  assign output_21_8 = io_outValid_8 & _T_64881; // @[Switch.scala 41:38:@26041.4]
  assign _T_64884 = select_9 == 6'h15; // @[Switch.scala 41:52:@26043.4]
  assign output_21_9 = io_outValid_9 & _T_64884; // @[Switch.scala 41:38:@26044.4]
  assign _T_64887 = select_10 == 6'h15; // @[Switch.scala 41:52:@26046.4]
  assign output_21_10 = io_outValid_10 & _T_64887; // @[Switch.scala 41:38:@26047.4]
  assign _T_64890 = select_11 == 6'h15; // @[Switch.scala 41:52:@26049.4]
  assign output_21_11 = io_outValid_11 & _T_64890; // @[Switch.scala 41:38:@26050.4]
  assign _T_64893 = select_12 == 6'h15; // @[Switch.scala 41:52:@26052.4]
  assign output_21_12 = io_outValid_12 & _T_64893; // @[Switch.scala 41:38:@26053.4]
  assign _T_64896 = select_13 == 6'h15; // @[Switch.scala 41:52:@26055.4]
  assign output_21_13 = io_outValid_13 & _T_64896; // @[Switch.scala 41:38:@26056.4]
  assign _T_64899 = select_14 == 6'h15; // @[Switch.scala 41:52:@26058.4]
  assign output_21_14 = io_outValid_14 & _T_64899; // @[Switch.scala 41:38:@26059.4]
  assign _T_64902 = select_15 == 6'h15; // @[Switch.scala 41:52:@26061.4]
  assign output_21_15 = io_outValid_15 & _T_64902; // @[Switch.scala 41:38:@26062.4]
  assign _T_64905 = select_16 == 6'h15; // @[Switch.scala 41:52:@26064.4]
  assign output_21_16 = io_outValid_16 & _T_64905; // @[Switch.scala 41:38:@26065.4]
  assign _T_64908 = select_17 == 6'h15; // @[Switch.scala 41:52:@26067.4]
  assign output_21_17 = io_outValid_17 & _T_64908; // @[Switch.scala 41:38:@26068.4]
  assign _T_64911 = select_18 == 6'h15; // @[Switch.scala 41:52:@26070.4]
  assign output_21_18 = io_outValid_18 & _T_64911; // @[Switch.scala 41:38:@26071.4]
  assign _T_64914 = select_19 == 6'h15; // @[Switch.scala 41:52:@26073.4]
  assign output_21_19 = io_outValid_19 & _T_64914; // @[Switch.scala 41:38:@26074.4]
  assign _T_64917 = select_20 == 6'h15; // @[Switch.scala 41:52:@26076.4]
  assign output_21_20 = io_outValid_20 & _T_64917; // @[Switch.scala 41:38:@26077.4]
  assign _T_64920 = select_21 == 6'h15; // @[Switch.scala 41:52:@26079.4]
  assign output_21_21 = io_outValid_21 & _T_64920; // @[Switch.scala 41:38:@26080.4]
  assign _T_64923 = select_22 == 6'h15; // @[Switch.scala 41:52:@26082.4]
  assign output_21_22 = io_outValid_22 & _T_64923; // @[Switch.scala 41:38:@26083.4]
  assign _T_64926 = select_23 == 6'h15; // @[Switch.scala 41:52:@26085.4]
  assign output_21_23 = io_outValid_23 & _T_64926; // @[Switch.scala 41:38:@26086.4]
  assign _T_64929 = select_24 == 6'h15; // @[Switch.scala 41:52:@26088.4]
  assign output_21_24 = io_outValid_24 & _T_64929; // @[Switch.scala 41:38:@26089.4]
  assign _T_64932 = select_25 == 6'h15; // @[Switch.scala 41:52:@26091.4]
  assign output_21_25 = io_outValid_25 & _T_64932; // @[Switch.scala 41:38:@26092.4]
  assign _T_64935 = select_26 == 6'h15; // @[Switch.scala 41:52:@26094.4]
  assign output_21_26 = io_outValid_26 & _T_64935; // @[Switch.scala 41:38:@26095.4]
  assign _T_64938 = select_27 == 6'h15; // @[Switch.scala 41:52:@26097.4]
  assign output_21_27 = io_outValid_27 & _T_64938; // @[Switch.scala 41:38:@26098.4]
  assign _T_64941 = select_28 == 6'h15; // @[Switch.scala 41:52:@26100.4]
  assign output_21_28 = io_outValid_28 & _T_64941; // @[Switch.scala 41:38:@26101.4]
  assign _T_64944 = select_29 == 6'h15; // @[Switch.scala 41:52:@26103.4]
  assign output_21_29 = io_outValid_29 & _T_64944; // @[Switch.scala 41:38:@26104.4]
  assign _T_64947 = select_30 == 6'h15; // @[Switch.scala 41:52:@26106.4]
  assign output_21_30 = io_outValid_30 & _T_64947; // @[Switch.scala 41:38:@26107.4]
  assign _T_64950 = select_31 == 6'h15; // @[Switch.scala 41:52:@26109.4]
  assign output_21_31 = io_outValid_31 & _T_64950; // @[Switch.scala 41:38:@26110.4]
  assign _T_64953 = select_32 == 6'h15; // @[Switch.scala 41:52:@26112.4]
  assign output_21_32 = io_outValid_32 & _T_64953; // @[Switch.scala 41:38:@26113.4]
  assign _T_64956 = select_33 == 6'h15; // @[Switch.scala 41:52:@26115.4]
  assign output_21_33 = io_outValid_33 & _T_64956; // @[Switch.scala 41:38:@26116.4]
  assign _T_64959 = select_34 == 6'h15; // @[Switch.scala 41:52:@26118.4]
  assign output_21_34 = io_outValid_34 & _T_64959; // @[Switch.scala 41:38:@26119.4]
  assign _T_64962 = select_35 == 6'h15; // @[Switch.scala 41:52:@26121.4]
  assign output_21_35 = io_outValid_35 & _T_64962; // @[Switch.scala 41:38:@26122.4]
  assign _T_64965 = select_36 == 6'h15; // @[Switch.scala 41:52:@26124.4]
  assign output_21_36 = io_outValid_36 & _T_64965; // @[Switch.scala 41:38:@26125.4]
  assign _T_64968 = select_37 == 6'h15; // @[Switch.scala 41:52:@26127.4]
  assign output_21_37 = io_outValid_37 & _T_64968; // @[Switch.scala 41:38:@26128.4]
  assign _T_64971 = select_38 == 6'h15; // @[Switch.scala 41:52:@26130.4]
  assign output_21_38 = io_outValid_38 & _T_64971; // @[Switch.scala 41:38:@26131.4]
  assign _T_64974 = select_39 == 6'h15; // @[Switch.scala 41:52:@26133.4]
  assign output_21_39 = io_outValid_39 & _T_64974; // @[Switch.scala 41:38:@26134.4]
  assign _T_64977 = select_40 == 6'h15; // @[Switch.scala 41:52:@26136.4]
  assign output_21_40 = io_outValid_40 & _T_64977; // @[Switch.scala 41:38:@26137.4]
  assign _T_64980 = select_41 == 6'h15; // @[Switch.scala 41:52:@26139.4]
  assign output_21_41 = io_outValid_41 & _T_64980; // @[Switch.scala 41:38:@26140.4]
  assign _T_64983 = select_42 == 6'h15; // @[Switch.scala 41:52:@26142.4]
  assign output_21_42 = io_outValid_42 & _T_64983; // @[Switch.scala 41:38:@26143.4]
  assign _T_64986 = select_43 == 6'h15; // @[Switch.scala 41:52:@26145.4]
  assign output_21_43 = io_outValid_43 & _T_64986; // @[Switch.scala 41:38:@26146.4]
  assign _T_64989 = select_44 == 6'h15; // @[Switch.scala 41:52:@26148.4]
  assign output_21_44 = io_outValid_44 & _T_64989; // @[Switch.scala 41:38:@26149.4]
  assign _T_64992 = select_45 == 6'h15; // @[Switch.scala 41:52:@26151.4]
  assign output_21_45 = io_outValid_45 & _T_64992; // @[Switch.scala 41:38:@26152.4]
  assign _T_64995 = select_46 == 6'h15; // @[Switch.scala 41:52:@26154.4]
  assign output_21_46 = io_outValid_46 & _T_64995; // @[Switch.scala 41:38:@26155.4]
  assign _T_64998 = select_47 == 6'h15; // @[Switch.scala 41:52:@26157.4]
  assign output_21_47 = io_outValid_47 & _T_64998; // @[Switch.scala 41:38:@26158.4]
  assign _T_65001 = select_48 == 6'h15; // @[Switch.scala 41:52:@26160.4]
  assign output_21_48 = io_outValid_48 & _T_65001; // @[Switch.scala 41:38:@26161.4]
  assign _T_65004 = select_49 == 6'h15; // @[Switch.scala 41:52:@26163.4]
  assign output_21_49 = io_outValid_49 & _T_65004; // @[Switch.scala 41:38:@26164.4]
  assign _T_65007 = select_50 == 6'h15; // @[Switch.scala 41:52:@26166.4]
  assign output_21_50 = io_outValid_50 & _T_65007; // @[Switch.scala 41:38:@26167.4]
  assign _T_65010 = select_51 == 6'h15; // @[Switch.scala 41:52:@26169.4]
  assign output_21_51 = io_outValid_51 & _T_65010; // @[Switch.scala 41:38:@26170.4]
  assign _T_65013 = select_52 == 6'h15; // @[Switch.scala 41:52:@26172.4]
  assign output_21_52 = io_outValid_52 & _T_65013; // @[Switch.scala 41:38:@26173.4]
  assign _T_65016 = select_53 == 6'h15; // @[Switch.scala 41:52:@26175.4]
  assign output_21_53 = io_outValid_53 & _T_65016; // @[Switch.scala 41:38:@26176.4]
  assign _T_65019 = select_54 == 6'h15; // @[Switch.scala 41:52:@26178.4]
  assign output_21_54 = io_outValid_54 & _T_65019; // @[Switch.scala 41:38:@26179.4]
  assign _T_65022 = select_55 == 6'h15; // @[Switch.scala 41:52:@26181.4]
  assign output_21_55 = io_outValid_55 & _T_65022; // @[Switch.scala 41:38:@26182.4]
  assign _T_65025 = select_56 == 6'h15; // @[Switch.scala 41:52:@26184.4]
  assign output_21_56 = io_outValid_56 & _T_65025; // @[Switch.scala 41:38:@26185.4]
  assign _T_65028 = select_57 == 6'h15; // @[Switch.scala 41:52:@26187.4]
  assign output_21_57 = io_outValid_57 & _T_65028; // @[Switch.scala 41:38:@26188.4]
  assign _T_65031 = select_58 == 6'h15; // @[Switch.scala 41:52:@26190.4]
  assign output_21_58 = io_outValid_58 & _T_65031; // @[Switch.scala 41:38:@26191.4]
  assign _T_65034 = select_59 == 6'h15; // @[Switch.scala 41:52:@26193.4]
  assign output_21_59 = io_outValid_59 & _T_65034; // @[Switch.scala 41:38:@26194.4]
  assign _T_65037 = select_60 == 6'h15; // @[Switch.scala 41:52:@26196.4]
  assign output_21_60 = io_outValid_60 & _T_65037; // @[Switch.scala 41:38:@26197.4]
  assign _T_65040 = select_61 == 6'h15; // @[Switch.scala 41:52:@26199.4]
  assign output_21_61 = io_outValid_61 & _T_65040; // @[Switch.scala 41:38:@26200.4]
  assign _T_65043 = select_62 == 6'h15; // @[Switch.scala 41:52:@26202.4]
  assign output_21_62 = io_outValid_62 & _T_65043; // @[Switch.scala 41:38:@26203.4]
  assign _T_65046 = select_63 == 6'h15; // @[Switch.scala 41:52:@26205.4]
  assign output_21_63 = io_outValid_63 & _T_65046; // @[Switch.scala 41:38:@26206.4]
  assign _T_65054 = {output_21_7,output_21_6,output_21_5,output_21_4,output_21_3,output_21_2,output_21_1,output_21_0}; // @[Switch.scala 43:31:@26214.4]
  assign _T_65062 = {output_21_15,output_21_14,output_21_13,output_21_12,output_21_11,output_21_10,output_21_9,output_21_8,_T_65054}; // @[Switch.scala 43:31:@26222.4]
  assign _T_65069 = {output_21_23,output_21_22,output_21_21,output_21_20,output_21_19,output_21_18,output_21_17,output_21_16}; // @[Switch.scala 43:31:@26229.4]
  assign _T_65078 = {output_21_31,output_21_30,output_21_29,output_21_28,output_21_27,output_21_26,output_21_25,output_21_24,_T_65069,_T_65062}; // @[Switch.scala 43:31:@26238.4]
  assign _T_65085 = {output_21_39,output_21_38,output_21_37,output_21_36,output_21_35,output_21_34,output_21_33,output_21_32}; // @[Switch.scala 43:31:@26245.4]
  assign _T_65093 = {output_21_47,output_21_46,output_21_45,output_21_44,output_21_43,output_21_42,output_21_41,output_21_40,_T_65085}; // @[Switch.scala 43:31:@26253.4]
  assign _T_65100 = {output_21_55,output_21_54,output_21_53,output_21_52,output_21_51,output_21_50,output_21_49,output_21_48}; // @[Switch.scala 43:31:@26260.4]
  assign _T_65109 = {output_21_63,output_21_62,output_21_61,output_21_60,output_21_59,output_21_58,output_21_57,output_21_56,_T_65100,_T_65093}; // @[Switch.scala 43:31:@26269.4]
  assign _T_65110 = {_T_65109,_T_65078}; // @[Switch.scala 43:31:@26270.4]
  assign _T_65114 = select_0 == 6'h16; // @[Switch.scala 41:52:@26273.4]
  assign output_22_0 = io_outValid_0 & _T_65114; // @[Switch.scala 41:38:@26274.4]
  assign _T_65117 = select_1 == 6'h16; // @[Switch.scala 41:52:@26276.4]
  assign output_22_1 = io_outValid_1 & _T_65117; // @[Switch.scala 41:38:@26277.4]
  assign _T_65120 = select_2 == 6'h16; // @[Switch.scala 41:52:@26279.4]
  assign output_22_2 = io_outValid_2 & _T_65120; // @[Switch.scala 41:38:@26280.4]
  assign _T_65123 = select_3 == 6'h16; // @[Switch.scala 41:52:@26282.4]
  assign output_22_3 = io_outValid_3 & _T_65123; // @[Switch.scala 41:38:@26283.4]
  assign _T_65126 = select_4 == 6'h16; // @[Switch.scala 41:52:@26285.4]
  assign output_22_4 = io_outValid_4 & _T_65126; // @[Switch.scala 41:38:@26286.4]
  assign _T_65129 = select_5 == 6'h16; // @[Switch.scala 41:52:@26288.4]
  assign output_22_5 = io_outValid_5 & _T_65129; // @[Switch.scala 41:38:@26289.4]
  assign _T_65132 = select_6 == 6'h16; // @[Switch.scala 41:52:@26291.4]
  assign output_22_6 = io_outValid_6 & _T_65132; // @[Switch.scala 41:38:@26292.4]
  assign _T_65135 = select_7 == 6'h16; // @[Switch.scala 41:52:@26294.4]
  assign output_22_7 = io_outValid_7 & _T_65135; // @[Switch.scala 41:38:@26295.4]
  assign _T_65138 = select_8 == 6'h16; // @[Switch.scala 41:52:@26297.4]
  assign output_22_8 = io_outValid_8 & _T_65138; // @[Switch.scala 41:38:@26298.4]
  assign _T_65141 = select_9 == 6'h16; // @[Switch.scala 41:52:@26300.4]
  assign output_22_9 = io_outValid_9 & _T_65141; // @[Switch.scala 41:38:@26301.4]
  assign _T_65144 = select_10 == 6'h16; // @[Switch.scala 41:52:@26303.4]
  assign output_22_10 = io_outValid_10 & _T_65144; // @[Switch.scala 41:38:@26304.4]
  assign _T_65147 = select_11 == 6'h16; // @[Switch.scala 41:52:@26306.4]
  assign output_22_11 = io_outValid_11 & _T_65147; // @[Switch.scala 41:38:@26307.4]
  assign _T_65150 = select_12 == 6'h16; // @[Switch.scala 41:52:@26309.4]
  assign output_22_12 = io_outValid_12 & _T_65150; // @[Switch.scala 41:38:@26310.4]
  assign _T_65153 = select_13 == 6'h16; // @[Switch.scala 41:52:@26312.4]
  assign output_22_13 = io_outValid_13 & _T_65153; // @[Switch.scala 41:38:@26313.4]
  assign _T_65156 = select_14 == 6'h16; // @[Switch.scala 41:52:@26315.4]
  assign output_22_14 = io_outValid_14 & _T_65156; // @[Switch.scala 41:38:@26316.4]
  assign _T_65159 = select_15 == 6'h16; // @[Switch.scala 41:52:@26318.4]
  assign output_22_15 = io_outValid_15 & _T_65159; // @[Switch.scala 41:38:@26319.4]
  assign _T_65162 = select_16 == 6'h16; // @[Switch.scala 41:52:@26321.4]
  assign output_22_16 = io_outValid_16 & _T_65162; // @[Switch.scala 41:38:@26322.4]
  assign _T_65165 = select_17 == 6'h16; // @[Switch.scala 41:52:@26324.4]
  assign output_22_17 = io_outValid_17 & _T_65165; // @[Switch.scala 41:38:@26325.4]
  assign _T_65168 = select_18 == 6'h16; // @[Switch.scala 41:52:@26327.4]
  assign output_22_18 = io_outValid_18 & _T_65168; // @[Switch.scala 41:38:@26328.4]
  assign _T_65171 = select_19 == 6'h16; // @[Switch.scala 41:52:@26330.4]
  assign output_22_19 = io_outValid_19 & _T_65171; // @[Switch.scala 41:38:@26331.4]
  assign _T_65174 = select_20 == 6'h16; // @[Switch.scala 41:52:@26333.4]
  assign output_22_20 = io_outValid_20 & _T_65174; // @[Switch.scala 41:38:@26334.4]
  assign _T_65177 = select_21 == 6'h16; // @[Switch.scala 41:52:@26336.4]
  assign output_22_21 = io_outValid_21 & _T_65177; // @[Switch.scala 41:38:@26337.4]
  assign _T_65180 = select_22 == 6'h16; // @[Switch.scala 41:52:@26339.4]
  assign output_22_22 = io_outValid_22 & _T_65180; // @[Switch.scala 41:38:@26340.4]
  assign _T_65183 = select_23 == 6'h16; // @[Switch.scala 41:52:@26342.4]
  assign output_22_23 = io_outValid_23 & _T_65183; // @[Switch.scala 41:38:@26343.4]
  assign _T_65186 = select_24 == 6'h16; // @[Switch.scala 41:52:@26345.4]
  assign output_22_24 = io_outValid_24 & _T_65186; // @[Switch.scala 41:38:@26346.4]
  assign _T_65189 = select_25 == 6'h16; // @[Switch.scala 41:52:@26348.4]
  assign output_22_25 = io_outValid_25 & _T_65189; // @[Switch.scala 41:38:@26349.4]
  assign _T_65192 = select_26 == 6'h16; // @[Switch.scala 41:52:@26351.4]
  assign output_22_26 = io_outValid_26 & _T_65192; // @[Switch.scala 41:38:@26352.4]
  assign _T_65195 = select_27 == 6'h16; // @[Switch.scala 41:52:@26354.4]
  assign output_22_27 = io_outValid_27 & _T_65195; // @[Switch.scala 41:38:@26355.4]
  assign _T_65198 = select_28 == 6'h16; // @[Switch.scala 41:52:@26357.4]
  assign output_22_28 = io_outValid_28 & _T_65198; // @[Switch.scala 41:38:@26358.4]
  assign _T_65201 = select_29 == 6'h16; // @[Switch.scala 41:52:@26360.4]
  assign output_22_29 = io_outValid_29 & _T_65201; // @[Switch.scala 41:38:@26361.4]
  assign _T_65204 = select_30 == 6'h16; // @[Switch.scala 41:52:@26363.4]
  assign output_22_30 = io_outValid_30 & _T_65204; // @[Switch.scala 41:38:@26364.4]
  assign _T_65207 = select_31 == 6'h16; // @[Switch.scala 41:52:@26366.4]
  assign output_22_31 = io_outValid_31 & _T_65207; // @[Switch.scala 41:38:@26367.4]
  assign _T_65210 = select_32 == 6'h16; // @[Switch.scala 41:52:@26369.4]
  assign output_22_32 = io_outValid_32 & _T_65210; // @[Switch.scala 41:38:@26370.4]
  assign _T_65213 = select_33 == 6'h16; // @[Switch.scala 41:52:@26372.4]
  assign output_22_33 = io_outValid_33 & _T_65213; // @[Switch.scala 41:38:@26373.4]
  assign _T_65216 = select_34 == 6'h16; // @[Switch.scala 41:52:@26375.4]
  assign output_22_34 = io_outValid_34 & _T_65216; // @[Switch.scala 41:38:@26376.4]
  assign _T_65219 = select_35 == 6'h16; // @[Switch.scala 41:52:@26378.4]
  assign output_22_35 = io_outValid_35 & _T_65219; // @[Switch.scala 41:38:@26379.4]
  assign _T_65222 = select_36 == 6'h16; // @[Switch.scala 41:52:@26381.4]
  assign output_22_36 = io_outValid_36 & _T_65222; // @[Switch.scala 41:38:@26382.4]
  assign _T_65225 = select_37 == 6'h16; // @[Switch.scala 41:52:@26384.4]
  assign output_22_37 = io_outValid_37 & _T_65225; // @[Switch.scala 41:38:@26385.4]
  assign _T_65228 = select_38 == 6'h16; // @[Switch.scala 41:52:@26387.4]
  assign output_22_38 = io_outValid_38 & _T_65228; // @[Switch.scala 41:38:@26388.4]
  assign _T_65231 = select_39 == 6'h16; // @[Switch.scala 41:52:@26390.4]
  assign output_22_39 = io_outValid_39 & _T_65231; // @[Switch.scala 41:38:@26391.4]
  assign _T_65234 = select_40 == 6'h16; // @[Switch.scala 41:52:@26393.4]
  assign output_22_40 = io_outValid_40 & _T_65234; // @[Switch.scala 41:38:@26394.4]
  assign _T_65237 = select_41 == 6'h16; // @[Switch.scala 41:52:@26396.4]
  assign output_22_41 = io_outValid_41 & _T_65237; // @[Switch.scala 41:38:@26397.4]
  assign _T_65240 = select_42 == 6'h16; // @[Switch.scala 41:52:@26399.4]
  assign output_22_42 = io_outValid_42 & _T_65240; // @[Switch.scala 41:38:@26400.4]
  assign _T_65243 = select_43 == 6'h16; // @[Switch.scala 41:52:@26402.4]
  assign output_22_43 = io_outValid_43 & _T_65243; // @[Switch.scala 41:38:@26403.4]
  assign _T_65246 = select_44 == 6'h16; // @[Switch.scala 41:52:@26405.4]
  assign output_22_44 = io_outValid_44 & _T_65246; // @[Switch.scala 41:38:@26406.4]
  assign _T_65249 = select_45 == 6'h16; // @[Switch.scala 41:52:@26408.4]
  assign output_22_45 = io_outValid_45 & _T_65249; // @[Switch.scala 41:38:@26409.4]
  assign _T_65252 = select_46 == 6'h16; // @[Switch.scala 41:52:@26411.4]
  assign output_22_46 = io_outValid_46 & _T_65252; // @[Switch.scala 41:38:@26412.4]
  assign _T_65255 = select_47 == 6'h16; // @[Switch.scala 41:52:@26414.4]
  assign output_22_47 = io_outValid_47 & _T_65255; // @[Switch.scala 41:38:@26415.4]
  assign _T_65258 = select_48 == 6'h16; // @[Switch.scala 41:52:@26417.4]
  assign output_22_48 = io_outValid_48 & _T_65258; // @[Switch.scala 41:38:@26418.4]
  assign _T_65261 = select_49 == 6'h16; // @[Switch.scala 41:52:@26420.4]
  assign output_22_49 = io_outValid_49 & _T_65261; // @[Switch.scala 41:38:@26421.4]
  assign _T_65264 = select_50 == 6'h16; // @[Switch.scala 41:52:@26423.4]
  assign output_22_50 = io_outValid_50 & _T_65264; // @[Switch.scala 41:38:@26424.4]
  assign _T_65267 = select_51 == 6'h16; // @[Switch.scala 41:52:@26426.4]
  assign output_22_51 = io_outValid_51 & _T_65267; // @[Switch.scala 41:38:@26427.4]
  assign _T_65270 = select_52 == 6'h16; // @[Switch.scala 41:52:@26429.4]
  assign output_22_52 = io_outValid_52 & _T_65270; // @[Switch.scala 41:38:@26430.4]
  assign _T_65273 = select_53 == 6'h16; // @[Switch.scala 41:52:@26432.4]
  assign output_22_53 = io_outValid_53 & _T_65273; // @[Switch.scala 41:38:@26433.4]
  assign _T_65276 = select_54 == 6'h16; // @[Switch.scala 41:52:@26435.4]
  assign output_22_54 = io_outValid_54 & _T_65276; // @[Switch.scala 41:38:@26436.4]
  assign _T_65279 = select_55 == 6'h16; // @[Switch.scala 41:52:@26438.4]
  assign output_22_55 = io_outValid_55 & _T_65279; // @[Switch.scala 41:38:@26439.4]
  assign _T_65282 = select_56 == 6'h16; // @[Switch.scala 41:52:@26441.4]
  assign output_22_56 = io_outValid_56 & _T_65282; // @[Switch.scala 41:38:@26442.4]
  assign _T_65285 = select_57 == 6'h16; // @[Switch.scala 41:52:@26444.4]
  assign output_22_57 = io_outValid_57 & _T_65285; // @[Switch.scala 41:38:@26445.4]
  assign _T_65288 = select_58 == 6'h16; // @[Switch.scala 41:52:@26447.4]
  assign output_22_58 = io_outValid_58 & _T_65288; // @[Switch.scala 41:38:@26448.4]
  assign _T_65291 = select_59 == 6'h16; // @[Switch.scala 41:52:@26450.4]
  assign output_22_59 = io_outValid_59 & _T_65291; // @[Switch.scala 41:38:@26451.4]
  assign _T_65294 = select_60 == 6'h16; // @[Switch.scala 41:52:@26453.4]
  assign output_22_60 = io_outValid_60 & _T_65294; // @[Switch.scala 41:38:@26454.4]
  assign _T_65297 = select_61 == 6'h16; // @[Switch.scala 41:52:@26456.4]
  assign output_22_61 = io_outValid_61 & _T_65297; // @[Switch.scala 41:38:@26457.4]
  assign _T_65300 = select_62 == 6'h16; // @[Switch.scala 41:52:@26459.4]
  assign output_22_62 = io_outValid_62 & _T_65300; // @[Switch.scala 41:38:@26460.4]
  assign _T_65303 = select_63 == 6'h16; // @[Switch.scala 41:52:@26462.4]
  assign output_22_63 = io_outValid_63 & _T_65303; // @[Switch.scala 41:38:@26463.4]
  assign _T_65311 = {output_22_7,output_22_6,output_22_5,output_22_4,output_22_3,output_22_2,output_22_1,output_22_0}; // @[Switch.scala 43:31:@26471.4]
  assign _T_65319 = {output_22_15,output_22_14,output_22_13,output_22_12,output_22_11,output_22_10,output_22_9,output_22_8,_T_65311}; // @[Switch.scala 43:31:@26479.4]
  assign _T_65326 = {output_22_23,output_22_22,output_22_21,output_22_20,output_22_19,output_22_18,output_22_17,output_22_16}; // @[Switch.scala 43:31:@26486.4]
  assign _T_65335 = {output_22_31,output_22_30,output_22_29,output_22_28,output_22_27,output_22_26,output_22_25,output_22_24,_T_65326,_T_65319}; // @[Switch.scala 43:31:@26495.4]
  assign _T_65342 = {output_22_39,output_22_38,output_22_37,output_22_36,output_22_35,output_22_34,output_22_33,output_22_32}; // @[Switch.scala 43:31:@26502.4]
  assign _T_65350 = {output_22_47,output_22_46,output_22_45,output_22_44,output_22_43,output_22_42,output_22_41,output_22_40,_T_65342}; // @[Switch.scala 43:31:@26510.4]
  assign _T_65357 = {output_22_55,output_22_54,output_22_53,output_22_52,output_22_51,output_22_50,output_22_49,output_22_48}; // @[Switch.scala 43:31:@26517.4]
  assign _T_65366 = {output_22_63,output_22_62,output_22_61,output_22_60,output_22_59,output_22_58,output_22_57,output_22_56,_T_65357,_T_65350}; // @[Switch.scala 43:31:@26526.4]
  assign _T_65367 = {_T_65366,_T_65335}; // @[Switch.scala 43:31:@26527.4]
  assign _T_65371 = select_0 == 6'h17; // @[Switch.scala 41:52:@26530.4]
  assign output_23_0 = io_outValid_0 & _T_65371; // @[Switch.scala 41:38:@26531.4]
  assign _T_65374 = select_1 == 6'h17; // @[Switch.scala 41:52:@26533.4]
  assign output_23_1 = io_outValid_1 & _T_65374; // @[Switch.scala 41:38:@26534.4]
  assign _T_65377 = select_2 == 6'h17; // @[Switch.scala 41:52:@26536.4]
  assign output_23_2 = io_outValid_2 & _T_65377; // @[Switch.scala 41:38:@26537.4]
  assign _T_65380 = select_3 == 6'h17; // @[Switch.scala 41:52:@26539.4]
  assign output_23_3 = io_outValid_3 & _T_65380; // @[Switch.scala 41:38:@26540.4]
  assign _T_65383 = select_4 == 6'h17; // @[Switch.scala 41:52:@26542.4]
  assign output_23_4 = io_outValid_4 & _T_65383; // @[Switch.scala 41:38:@26543.4]
  assign _T_65386 = select_5 == 6'h17; // @[Switch.scala 41:52:@26545.4]
  assign output_23_5 = io_outValid_5 & _T_65386; // @[Switch.scala 41:38:@26546.4]
  assign _T_65389 = select_6 == 6'h17; // @[Switch.scala 41:52:@26548.4]
  assign output_23_6 = io_outValid_6 & _T_65389; // @[Switch.scala 41:38:@26549.4]
  assign _T_65392 = select_7 == 6'h17; // @[Switch.scala 41:52:@26551.4]
  assign output_23_7 = io_outValid_7 & _T_65392; // @[Switch.scala 41:38:@26552.4]
  assign _T_65395 = select_8 == 6'h17; // @[Switch.scala 41:52:@26554.4]
  assign output_23_8 = io_outValid_8 & _T_65395; // @[Switch.scala 41:38:@26555.4]
  assign _T_65398 = select_9 == 6'h17; // @[Switch.scala 41:52:@26557.4]
  assign output_23_9 = io_outValid_9 & _T_65398; // @[Switch.scala 41:38:@26558.4]
  assign _T_65401 = select_10 == 6'h17; // @[Switch.scala 41:52:@26560.4]
  assign output_23_10 = io_outValid_10 & _T_65401; // @[Switch.scala 41:38:@26561.4]
  assign _T_65404 = select_11 == 6'h17; // @[Switch.scala 41:52:@26563.4]
  assign output_23_11 = io_outValid_11 & _T_65404; // @[Switch.scala 41:38:@26564.4]
  assign _T_65407 = select_12 == 6'h17; // @[Switch.scala 41:52:@26566.4]
  assign output_23_12 = io_outValid_12 & _T_65407; // @[Switch.scala 41:38:@26567.4]
  assign _T_65410 = select_13 == 6'h17; // @[Switch.scala 41:52:@26569.4]
  assign output_23_13 = io_outValid_13 & _T_65410; // @[Switch.scala 41:38:@26570.4]
  assign _T_65413 = select_14 == 6'h17; // @[Switch.scala 41:52:@26572.4]
  assign output_23_14 = io_outValid_14 & _T_65413; // @[Switch.scala 41:38:@26573.4]
  assign _T_65416 = select_15 == 6'h17; // @[Switch.scala 41:52:@26575.4]
  assign output_23_15 = io_outValid_15 & _T_65416; // @[Switch.scala 41:38:@26576.4]
  assign _T_65419 = select_16 == 6'h17; // @[Switch.scala 41:52:@26578.4]
  assign output_23_16 = io_outValid_16 & _T_65419; // @[Switch.scala 41:38:@26579.4]
  assign _T_65422 = select_17 == 6'h17; // @[Switch.scala 41:52:@26581.4]
  assign output_23_17 = io_outValid_17 & _T_65422; // @[Switch.scala 41:38:@26582.4]
  assign _T_65425 = select_18 == 6'h17; // @[Switch.scala 41:52:@26584.4]
  assign output_23_18 = io_outValid_18 & _T_65425; // @[Switch.scala 41:38:@26585.4]
  assign _T_65428 = select_19 == 6'h17; // @[Switch.scala 41:52:@26587.4]
  assign output_23_19 = io_outValid_19 & _T_65428; // @[Switch.scala 41:38:@26588.4]
  assign _T_65431 = select_20 == 6'h17; // @[Switch.scala 41:52:@26590.4]
  assign output_23_20 = io_outValid_20 & _T_65431; // @[Switch.scala 41:38:@26591.4]
  assign _T_65434 = select_21 == 6'h17; // @[Switch.scala 41:52:@26593.4]
  assign output_23_21 = io_outValid_21 & _T_65434; // @[Switch.scala 41:38:@26594.4]
  assign _T_65437 = select_22 == 6'h17; // @[Switch.scala 41:52:@26596.4]
  assign output_23_22 = io_outValid_22 & _T_65437; // @[Switch.scala 41:38:@26597.4]
  assign _T_65440 = select_23 == 6'h17; // @[Switch.scala 41:52:@26599.4]
  assign output_23_23 = io_outValid_23 & _T_65440; // @[Switch.scala 41:38:@26600.4]
  assign _T_65443 = select_24 == 6'h17; // @[Switch.scala 41:52:@26602.4]
  assign output_23_24 = io_outValid_24 & _T_65443; // @[Switch.scala 41:38:@26603.4]
  assign _T_65446 = select_25 == 6'h17; // @[Switch.scala 41:52:@26605.4]
  assign output_23_25 = io_outValid_25 & _T_65446; // @[Switch.scala 41:38:@26606.4]
  assign _T_65449 = select_26 == 6'h17; // @[Switch.scala 41:52:@26608.4]
  assign output_23_26 = io_outValid_26 & _T_65449; // @[Switch.scala 41:38:@26609.4]
  assign _T_65452 = select_27 == 6'h17; // @[Switch.scala 41:52:@26611.4]
  assign output_23_27 = io_outValid_27 & _T_65452; // @[Switch.scala 41:38:@26612.4]
  assign _T_65455 = select_28 == 6'h17; // @[Switch.scala 41:52:@26614.4]
  assign output_23_28 = io_outValid_28 & _T_65455; // @[Switch.scala 41:38:@26615.4]
  assign _T_65458 = select_29 == 6'h17; // @[Switch.scala 41:52:@26617.4]
  assign output_23_29 = io_outValid_29 & _T_65458; // @[Switch.scala 41:38:@26618.4]
  assign _T_65461 = select_30 == 6'h17; // @[Switch.scala 41:52:@26620.4]
  assign output_23_30 = io_outValid_30 & _T_65461; // @[Switch.scala 41:38:@26621.4]
  assign _T_65464 = select_31 == 6'h17; // @[Switch.scala 41:52:@26623.4]
  assign output_23_31 = io_outValid_31 & _T_65464; // @[Switch.scala 41:38:@26624.4]
  assign _T_65467 = select_32 == 6'h17; // @[Switch.scala 41:52:@26626.4]
  assign output_23_32 = io_outValid_32 & _T_65467; // @[Switch.scala 41:38:@26627.4]
  assign _T_65470 = select_33 == 6'h17; // @[Switch.scala 41:52:@26629.4]
  assign output_23_33 = io_outValid_33 & _T_65470; // @[Switch.scala 41:38:@26630.4]
  assign _T_65473 = select_34 == 6'h17; // @[Switch.scala 41:52:@26632.4]
  assign output_23_34 = io_outValid_34 & _T_65473; // @[Switch.scala 41:38:@26633.4]
  assign _T_65476 = select_35 == 6'h17; // @[Switch.scala 41:52:@26635.4]
  assign output_23_35 = io_outValid_35 & _T_65476; // @[Switch.scala 41:38:@26636.4]
  assign _T_65479 = select_36 == 6'h17; // @[Switch.scala 41:52:@26638.4]
  assign output_23_36 = io_outValid_36 & _T_65479; // @[Switch.scala 41:38:@26639.4]
  assign _T_65482 = select_37 == 6'h17; // @[Switch.scala 41:52:@26641.4]
  assign output_23_37 = io_outValid_37 & _T_65482; // @[Switch.scala 41:38:@26642.4]
  assign _T_65485 = select_38 == 6'h17; // @[Switch.scala 41:52:@26644.4]
  assign output_23_38 = io_outValid_38 & _T_65485; // @[Switch.scala 41:38:@26645.4]
  assign _T_65488 = select_39 == 6'h17; // @[Switch.scala 41:52:@26647.4]
  assign output_23_39 = io_outValid_39 & _T_65488; // @[Switch.scala 41:38:@26648.4]
  assign _T_65491 = select_40 == 6'h17; // @[Switch.scala 41:52:@26650.4]
  assign output_23_40 = io_outValid_40 & _T_65491; // @[Switch.scala 41:38:@26651.4]
  assign _T_65494 = select_41 == 6'h17; // @[Switch.scala 41:52:@26653.4]
  assign output_23_41 = io_outValid_41 & _T_65494; // @[Switch.scala 41:38:@26654.4]
  assign _T_65497 = select_42 == 6'h17; // @[Switch.scala 41:52:@26656.4]
  assign output_23_42 = io_outValid_42 & _T_65497; // @[Switch.scala 41:38:@26657.4]
  assign _T_65500 = select_43 == 6'h17; // @[Switch.scala 41:52:@26659.4]
  assign output_23_43 = io_outValid_43 & _T_65500; // @[Switch.scala 41:38:@26660.4]
  assign _T_65503 = select_44 == 6'h17; // @[Switch.scala 41:52:@26662.4]
  assign output_23_44 = io_outValid_44 & _T_65503; // @[Switch.scala 41:38:@26663.4]
  assign _T_65506 = select_45 == 6'h17; // @[Switch.scala 41:52:@26665.4]
  assign output_23_45 = io_outValid_45 & _T_65506; // @[Switch.scala 41:38:@26666.4]
  assign _T_65509 = select_46 == 6'h17; // @[Switch.scala 41:52:@26668.4]
  assign output_23_46 = io_outValid_46 & _T_65509; // @[Switch.scala 41:38:@26669.4]
  assign _T_65512 = select_47 == 6'h17; // @[Switch.scala 41:52:@26671.4]
  assign output_23_47 = io_outValid_47 & _T_65512; // @[Switch.scala 41:38:@26672.4]
  assign _T_65515 = select_48 == 6'h17; // @[Switch.scala 41:52:@26674.4]
  assign output_23_48 = io_outValid_48 & _T_65515; // @[Switch.scala 41:38:@26675.4]
  assign _T_65518 = select_49 == 6'h17; // @[Switch.scala 41:52:@26677.4]
  assign output_23_49 = io_outValid_49 & _T_65518; // @[Switch.scala 41:38:@26678.4]
  assign _T_65521 = select_50 == 6'h17; // @[Switch.scala 41:52:@26680.4]
  assign output_23_50 = io_outValid_50 & _T_65521; // @[Switch.scala 41:38:@26681.4]
  assign _T_65524 = select_51 == 6'h17; // @[Switch.scala 41:52:@26683.4]
  assign output_23_51 = io_outValid_51 & _T_65524; // @[Switch.scala 41:38:@26684.4]
  assign _T_65527 = select_52 == 6'h17; // @[Switch.scala 41:52:@26686.4]
  assign output_23_52 = io_outValid_52 & _T_65527; // @[Switch.scala 41:38:@26687.4]
  assign _T_65530 = select_53 == 6'h17; // @[Switch.scala 41:52:@26689.4]
  assign output_23_53 = io_outValid_53 & _T_65530; // @[Switch.scala 41:38:@26690.4]
  assign _T_65533 = select_54 == 6'h17; // @[Switch.scala 41:52:@26692.4]
  assign output_23_54 = io_outValid_54 & _T_65533; // @[Switch.scala 41:38:@26693.4]
  assign _T_65536 = select_55 == 6'h17; // @[Switch.scala 41:52:@26695.4]
  assign output_23_55 = io_outValid_55 & _T_65536; // @[Switch.scala 41:38:@26696.4]
  assign _T_65539 = select_56 == 6'h17; // @[Switch.scala 41:52:@26698.4]
  assign output_23_56 = io_outValid_56 & _T_65539; // @[Switch.scala 41:38:@26699.4]
  assign _T_65542 = select_57 == 6'h17; // @[Switch.scala 41:52:@26701.4]
  assign output_23_57 = io_outValid_57 & _T_65542; // @[Switch.scala 41:38:@26702.4]
  assign _T_65545 = select_58 == 6'h17; // @[Switch.scala 41:52:@26704.4]
  assign output_23_58 = io_outValid_58 & _T_65545; // @[Switch.scala 41:38:@26705.4]
  assign _T_65548 = select_59 == 6'h17; // @[Switch.scala 41:52:@26707.4]
  assign output_23_59 = io_outValid_59 & _T_65548; // @[Switch.scala 41:38:@26708.4]
  assign _T_65551 = select_60 == 6'h17; // @[Switch.scala 41:52:@26710.4]
  assign output_23_60 = io_outValid_60 & _T_65551; // @[Switch.scala 41:38:@26711.4]
  assign _T_65554 = select_61 == 6'h17; // @[Switch.scala 41:52:@26713.4]
  assign output_23_61 = io_outValid_61 & _T_65554; // @[Switch.scala 41:38:@26714.4]
  assign _T_65557 = select_62 == 6'h17; // @[Switch.scala 41:52:@26716.4]
  assign output_23_62 = io_outValid_62 & _T_65557; // @[Switch.scala 41:38:@26717.4]
  assign _T_65560 = select_63 == 6'h17; // @[Switch.scala 41:52:@26719.4]
  assign output_23_63 = io_outValid_63 & _T_65560; // @[Switch.scala 41:38:@26720.4]
  assign _T_65568 = {output_23_7,output_23_6,output_23_5,output_23_4,output_23_3,output_23_2,output_23_1,output_23_0}; // @[Switch.scala 43:31:@26728.4]
  assign _T_65576 = {output_23_15,output_23_14,output_23_13,output_23_12,output_23_11,output_23_10,output_23_9,output_23_8,_T_65568}; // @[Switch.scala 43:31:@26736.4]
  assign _T_65583 = {output_23_23,output_23_22,output_23_21,output_23_20,output_23_19,output_23_18,output_23_17,output_23_16}; // @[Switch.scala 43:31:@26743.4]
  assign _T_65592 = {output_23_31,output_23_30,output_23_29,output_23_28,output_23_27,output_23_26,output_23_25,output_23_24,_T_65583,_T_65576}; // @[Switch.scala 43:31:@26752.4]
  assign _T_65599 = {output_23_39,output_23_38,output_23_37,output_23_36,output_23_35,output_23_34,output_23_33,output_23_32}; // @[Switch.scala 43:31:@26759.4]
  assign _T_65607 = {output_23_47,output_23_46,output_23_45,output_23_44,output_23_43,output_23_42,output_23_41,output_23_40,_T_65599}; // @[Switch.scala 43:31:@26767.4]
  assign _T_65614 = {output_23_55,output_23_54,output_23_53,output_23_52,output_23_51,output_23_50,output_23_49,output_23_48}; // @[Switch.scala 43:31:@26774.4]
  assign _T_65623 = {output_23_63,output_23_62,output_23_61,output_23_60,output_23_59,output_23_58,output_23_57,output_23_56,_T_65614,_T_65607}; // @[Switch.scala 43:31:@26783.4]
  assign _T_65624 = {_T_65623,_T_65592}; // @[Switch.scala 43:31:@26784.4]
  assign _T_65628 = select_0 == 6'h18; // @[Switch.scala 41:52:@26787.4]
  assign output_24_0 = io_outValid_0 & _T_65628; // @[Switch.scala 41:38:@26788.4]
  assign _T_65631 = select_1 == 6'h18; // @[Switch.scala 41:52:@26790.4]
  assign output_24_1 = io_outValid_1 & _T_65631; // @[Switch.scala 41:38:@26791.4]
  assign _T_65634 = select_2 == 6'h18; // @[Switch.scala 41:52:@26793.4]
  assign output_24_2 = io_outValid_2 & _T_65634; // @[Switch.scala 41:38:@26794.4]
  assign _T_65637 = select_3 == 6'h18; // @[Switch.scala 41:52:@26796.4]
  assign output_24_3 = io_outValid_3 & _T_65637; // @[Switch.scala 41:38:@26797.4]
  assign _T_65640 = select_4 == 6'h18; // @[Switch.scala 41:52:@26799.4]
  assign output_24_4 = io_outValid_4 & _T_65640; // @[Switch.scala 41:38:@26800.4]
  assign _T_65643 = select_5 == 6'h18; // @[Switch.scala 41:52:@26802.4]
  assign output_24_5 = io_outValid_5 & _T_65643; // @[Switch.scala 41:38:@26803.4]
  assign _T_65646 = select_6 == 6'h18; // @[Switch.scala 41:52:@26805.4]
  assign output_24_6 = io_outValid_6 & _T_65646; // @[Switch.scala 41:38:@26806.4]
  assign _T_65649 = select_7 == 6'h18; // @[Switch.scala 41:52:@26808.4]
  assign output_24_7 = io_outValid_7 & _T_65649; // @[Switch.scala 41:38:@26809.4]
  assign _T_65652 = select_8 == 6'h18; // @[Switch.scala 41:52:@26811.4]
  assign output_24_8 = io_outValid_8 & _T_65652; // @[Switch.scala 41:38:@26812.4]
  assign _T_65655 = select_9 == 6'h18; // @[Switch.scala 41:52:@26814.4]
  assign output_24_9 = io_outValid_9 & _T_65655; // @[Switch.scala 41:38:@26815.4]
  assign _T_65658 = select_10 == 6'h18; // @[Switch.scala 41:52:@26817.4]
  assign output_24_10 = io_outValid_10 & _T_65658; // @[Switch.scala 41:38:@26818.4]
  assign _T_65661 = select_11 == 6'h18; // @[Switch.scala 41:52:@26820.4]
  assign output_24_11 = io_outValid_11 & _T_65661; // @[Switch.scala 41:38:@26821.4]
  assign _T_65664 = select_12 == 6'h18; // @[Switch.scala 41:52:@26823.4]
  assign output_24_12 = io_outValid_12 & _T_65664; // @[Switch.scala 41:38:@26824.4]
  assign _T_65667 = select_13 == 6'h18; // @[Switch.scala 41:52:@26826.4]
  assign output_24_13 = io_outValid_13 & _T_65667; // @[Switch.scala 41:38:@26827.4]
  assign _T_65670 = select_14 == 6'h18; // @[Switch.scala 41:52:@26829.4]
  assign output_24_14 = io_outValid_14 & _T_65670; // @[Switch.scala 41:38:@26830.4]
  assign _T_65673 = select_15 == 6'h18; // @[Switch.scala 41:52:@26832.4]
  assign output_24_15 = io_outValid_15 & _T_65673; // @[Switch.scala 41:38:@26833.4]
  assign _T_65676 = select_16 == 6'h18; // @[Switch.scala 41:52:@26835.4]
  assign output_24_16 = io_outValid_16 & _T_65676; // @[Switch.scala 41:38:@26836.4]
  assign _T_65679 = select_17 == 6'h18; // @[Switch.scala 41:52:@26838.4]
  assign output_24_17 = io_outValid_17 & _T_65679; // @[Switch.scala 41:38:@26839.4]
  assign _T_65682 = select_18 == 6'h18; // @[Switch.scala 41:52:@26841.4]
  assign output_24_18 = io_outValid_18 & _T_65682; // @[Switch.scala 41:38:@26842.4]
  assign _T_65685 = select_19 == 6'h18; // @[Switch.scala 41:52:@26844.4]
  assign output_24_19 = io_outValid_19 & _T_65685; // @[Switch.scala 41:38:@26845.4]
  assign _T_65688 = select_20 == 6'h18; // @[Switch.scala 41:52:@26847.4]
  assign output_24_20 = io_outValid_20 & _T_65688; // @[Switch.scala 41:38:@26848.4]
  assign _T_65691 = select_21 == 6'h18; // @[Switch.scala 41:52:@26850.4]
  assign output_24_21 = io_outValid_21 & _T_65691; // @[Switch.scala 41:38:@26851.4]
  assign _T_65694 = select_22 == 6'h18; // @[Switch.scala 41:52:@26853.4]
  assign output_24_22 = io_outValid_22 & _T_65694; // @[Switch.scala 41:38:@26854.4]
  assign _T_65697 = select_23 == 6'h18; // @[Switch.scala 41:52:@26856.4]
  assign output_24_23 = io_outValid_23 & _T_65697; // @[Switch.scala 41:38:@26857.4]
  assign _T_65700 = select_24 == 6'h18; // @[Switch.scala 41:52:@26859.4]
  assign output_24_24 = io_outValid_24 & _T_65700; // @[Switch.scala 41:38:@26860.4]
  assign _T_65703 = select_25 == 6'h18; // @[Switch.scala 41:52:@26862.4]
  assign output_24_25 = io_outValid_25 & _T_65703; // @[Switch.scala 41:38:@26863.4]
  assign _T_65706 = select_26 == 6'h18; // @[Switch.scala 41:52:@26865.4]
  assign output_24_26 = io_outValid_26 & _T_65706; // @[Switch.scala 41:38:@26866.4]
  assign _T_65709 = select_27 == 6'h18; // @[Switch.scala 41:52:@26868.4]
  assign output_24_27 = io_outValid_27 & _T_65709; // @[Switch.scala 41:38:@26869.4]
  assign _T_65712 = select_28 == 6'h18; // @[Switch.scala 41:52:@26871.4]
  assign output_24_28 = io_outValid_28 & _T_65712; // @[Switch.scala 41:38:@26872.4]
  assign _T_65715 = select_29 == 6'h18; // @[Switch.scala 41:52:@26874.4]
  assign output_24_29 = io_outValid_29 & _T_65715; // @[Switch.scala 41:38:@26875.4]
  assign _T_65718 = select_30 == 6'h18; // @[Switch.scala 41:52:@26877.4]
  assign output_24_30 = io_outValid_30 & _T_65718; // @[Switch.scala 41:38:@26878.4]
  assign _T_65721 = select_31 == 6'h18; // @[Switch.scala 41:52:@26880.4]
  assign output_24_31 = io_outValid_31 & _T_65721; // @[Switch.scala 41:38:@26881.4]
  assign _T_65724 = select_32 == 6'h18; // @[Switch.scala 41:52:@26883.4]
  assign output_24_32 = io_outValid_32 & _T_65724; // @[Switch.scala 41:38:@26884.4]
  assign _T_65727 = select_33 == 6'h18; // @[Switch.scala 41:52:@26886.4]
  assign output_24_33 = io_outValid_33 & _T_65727; // @[Switch.scala 41:38:@26887.4]
  assign _T_65730 = select_34 == 6'h18; // @[Switch.scala 41:52:@26889.4]
  assign output_24_34 = io_outValid_34 & _T_65730; // @[Switch.scala 41:38:@26890.4]
  assign _T_65733 = select_35 == 6'h18; // @[Switch.scala 41:52:@26892.4]
  assign output_24_35 = io_outValid_35 & _T_65733; // @[Switch.scala 41:38:@26893.4]
  assign _T_65736 = select_36 == 6'h18; // @[Switch.scala 41:52:@26895.4]
  assign output_24_36 = io_outValid_36 & _T_65736; // @[Switch.scala 41:38:@26896.4]
  assign _T_65739 = select_37 == 6'h18; // @[Switch.scala 41:52:@26898.4]
  assign output_24_37 = io_outValid_37 & _T_65739; // @[Switch.scala 41:38:@26899.4]
  assign _T_65742 = select_38 == 6'h18; // @[Switch.scala 41:52:@26901.4]
  assign output_24_38 = io_outValid_38 & _T_65742; // @[Switch.scala 41:38:@26902.4]
  assign _T_65745 = select_39 == 6'h18; // @[Switch.scala 41:52:@26904.4]
  assign output_24_39 = io_outValid_39 & _T_65745; // @[Switch.scala 41:38:@26905.4]
  assign _T_65748 = select_40 == 6'h18; // @[Switch.scala 41:52:@26907.4]
  assign output_24_40 = io_outValid_40 & _T_65748; // @[Switch.scala 41:38:@26908.4]
  assign _T_65751 = select_41 == 6'h18; // @[Switch.scala 41:52:@26910.4]
  assign output_24_41 = io_outValid_41 & _T_65751; // @[Switch.scala 41:38:@26911.4]
  assign _T_65754 = select_42 == 6'h18; // @[Switch.scala 41:52:@26913.4]
  assign output_24_42 = io_outValid_42 & _T_65754; // @[Switch.scala 41:38:@26914.4]
  assign _T_65757 = select_43 == 6'h18; // @[Switch.scala 41:52:@26916.4]
  assign output_24_43 = io_outValid_43 & _T_65757; // @[Switch.scala 41:38:@26917.4]
  assign _T_65760 = select_44 == 6'h18; // @[Switch.scala 41:52:@26919.4]
  assign output_24_44 = io_outValid_44 & _T_65760; // @[Switch.scala 41:38:@26920.4]
  assign _T_65763 = select_45 == 6'h18; // @[Switch.scala 41:52:@26922.4]
  assign output_24_45 = io_outValid_45 & _T_65763; // @[Switch.scala 41:38:@26923.4]
  assign _T_65766 = select_46 == 6'h18; // @[Switch.scala 41:52:@26925.4]
  assign output_24_46 = io_outValid_46 & _T_65766; // @[Switch.scala 41:38:@26926.4]
  assign _T_65769 = select_47 == 6'h18; // @[Switch.scala 41:52:@26928.4]
  assign output_24_47 = io_outValid_47 & _T_65769; // @[Switch.scala 41:38:@26929.4]
  assign _T_65772 = select_48 == 6'h18; // @[Switch.scala 41:52:@26931.4]
  assign output_24_48 = io_outValid_48 & _T_65772; // @[Switch.scala 41:38:@26932.4]
  assign _T_65775 = select_49 == 6'h18; // @[Switch.scala 41:52:@26934.4]
  assign output_24_49 = io_outValid_49 & _T_65775; // @[Switch.scala 41:38:@26935.4]
  assign _T_65778 = select_50 == 6'h18; // @[Switch.scala 41:52:@26937.4]
  assign output_24_50 = io_outValid_50 & _T_65778; // @[Switch.scala 41:38:@26938.4]
  assign _T_65781 = select_51 == 6'h18; // @[Switch.scala 41:52:@26940.4]
  assign output_24_51 = io_outValid_51 & _T_65781; // @[Switch.scala 41:38:@26941.4]
  assign _T_65784 = select_52 == 6'h18; // @[Switch.scala 41:52:@26943.4]
  assign output_24_52 = io_outValid_52 & _T_65784; // @[Switch.scala 41:38:@26944.4]
  assign _T_65787 = select_53 == 6'h18; // @[Switch.scala 41:52:@26946.4]
  assign output_24_53 = io_outValid_53 & _T_65787; // @[Switch.scala 41:38:@26947.4]
  assign _T_65790 = select_54 == 6'h18; // @[Switch.scala 41:52:@26949.4]
  assign output_24_54 = io_outValid_54 & _T_65790; // @[Switch.scala 41:38:@26950.4]
  assign _T_65793 = select_55 == 6'h18; // @[Switch.scala 41:52:@26952.4]
  assign output_24_55 = io_outValid_55 & _T_65793; // @[Switch.scala 41:38:@26953.4]
  assign _T_65796 = select_56 == 6'h18; // @[Switch.scala 41:52:@26955.4]
  assign output_24_56 = io_outValid_56 & _T_65796; // @[Switch.scala 41:38:@26956.4]
  assign _T_65799 = select_57 == 6'h18; // @[Switch.scala 41:52:@26958.4]
  assign output_24_57 = io_outValid_57 & _T_65799; // @[Switch.scala 41:38:@26959.4]
  assign _T_65802 = select_58 == 6'h18; // @[Switch.scala 41:52:@26961.4]
  assign output_24_58 = io_outValid_58 & _T_65802; // @[Switch.scala 41:38:@26962.4]
  assign _T_65805 = select_59 == 6'h18; // @[Switch.scala 41:52:@26964.4]
  assign output_24_59 = io_outValid_59 & _T_65805; // @[Switch.scala 41:38:@26965.4]
  assign _T_65808 = select_60 == 6'h18; // @[Switch.scala 41:52:@26967.4]
  assign output_24_60 = io_outValid_60 & _T_65808; // @[Switch.scala 41:38:@26968.4]
  assign _T_65811 = select_61 == 6'h18; // @[Switch.scala 41:52:@26970.4]
  assign output_24_61 = io_outValid_61 & _T_65811; // @[Switch.scala 41:38:@26971.4]
  assign _T_65814 = select_62 == 6'h18; // @[Switch.scala 41:52:@26973.4]
  assign output_24_62 = io_outValid_62 & _T_65814; // @[Switch.scala 41:38:@26974.4]
  assign _T_65817 = select_63 == 6'h18; // @[Switch.scala 41:52:@26976.4]
  assign output_24_63 = io_outValid_63 & _T_65817; // @[Switch.scala 41:38:@26977.4]
  assign _T_65825 = {output_24_7,output_24_6,output_24_5,output_24_4,output_24_3,output_24_2,output_24_1,output_24_0}; // @[Switch.scala 43:31:@26985.4]
  assign _T_65833 = {output_24_15,output_24_14,output_24_13,output_24_12,output_24_11,output_24_10,output_24_9,output_24_8,_T_65825}; // @[Switch.scala 43:31:@26993.4]
  assign _T_65840 = {output_24_23,output_24_22,output_24_21,output_24_20,output_24_19,output_24_18,output_24_17,output_24_16}; // @[Switch.scala 43:31:@27000.4]
  assign _T_65849 = {output_24_31,output_24_30,output_24_29,output_24_28,output_24_27,output_24_26,output_24_25,output_24_24,_T_65840,_T_65833}; // @[Switch.scala 43:31:@27009.4]
  assign _T_65856 = {output_24_39,output_24_38,output_24_37,output_24_36,output_24_35,output_24_34,output_24_33,output_24_32}; // @[Switch.scala 43:31:@27016.4]
  assign _T_65864 = {output_24_47,output_24_46,output_24_45,output_24_44,output_24_43,output_24_42,output_24_41,output_24_40,_T_65856}; // @[Switch.scala 43:31:@27024.4]
  assign _T_65871 = {output_24_55,output_24_54,output_24_53,output_24_52,output_24_51,output_24_50,output_24_49,output_24_48}; // @[Switch.scala 43:31:@27031.4]
  assign _T_65880 = {output_24_63,output_24_62,output_24_61,output_24_60,output_24_59,output_24_58,output_24_57,output_24_56,_T_65871,_T_65864}; // @[Switch.scala 43:31:@27040.4]
  assign _T_65881 = {_T_65880,_T_65849}; // @[Switch.scala 43:31:@27041.4]
  assign _T_65885 = select_0 == 6'h19; // @[Switch.scala 41:52:@27044.4]
  assign output_25_0 = io_outValid_0 & _T_65885; // @[Switch.scala 41:38:@27045.4]
  assign _T_65888 = select_1 == 6'h19; // @[Switch.scala 41:52:@27047.4]
  assign output_25_1 = io_outValid_1 & _T_65888; // @[Switch.scala 41:38:@27048.4]
  assign _T_65891 = select_2 == 6'h19; // @[Switch.scala 41:52:@27050.4]
  assign output_25_2 = io_outValid_2 & _T_65891; // @[Switch.scala 41:38:@27051.4]
  assign _T_65894 = select_3 == 6'h19; // @[Switch.scala 41:52:@27053.4]
  assign output_25_3 = io_outValid_3 & _T_65894; // @[Switch.scala 41:38:@27054.4]
  assign _T_65897 = select_4 == 6'h19; // @[Switch.scala 41:52:@27056.4]
  assign output_25_4 = io_outValid_4 & _T_65897; // @[Switch.scala 41:38:@27057.4]
  assign _T_65900 = select_5 == 6'h19; // @[Switch.scala 41:52:@27059.4]
  assign output_25_5 = io_outValid_5 & _T_65900; // @[Switch.scala 41:38:@27060.4]
  assign _T_65903 = select_6 == 6'h19; // @[Switch.scala 41:52:@27062.4]
  assign output_25_6 = io_outValid_6 & _T_65903; // @[Switch.scala 41:38:@27063.4]
  assign _T_65906 = select_7 == 6'h19; // @[Switch.scala 41:52:@27065.4]
  assign output_25_7 = io_outValid_7 & _T_65906; // @[Switch.scala 41:38:@27066.4]
  assign _T_65909 = select_8 == 6'h19; // @[Switch.scala 41:52:@27068.4]
  assign output_25_8 = io_outValid_8 & _T_65909; // @[Switch.scala 41:38:@27069.4]
  assign _T_65912 = select_9 == 6'h19; // @[Switch.scala 41:52:@27071.4]
  assign output_25_9 = io_outValid_9 & _T_65912; // @[Switch.scala 41:38:@27072.4]
  assign _T_65915 = select_10 == 6'h19; // @[Switch.scala 41:52:@27074.4]
  assign output_25_10 = io_outValid_10 & _T_65915; // @[Switch.scala 41:38:@27075.4]
  assign _T_65918 = select_11 == 6'h19; // @[Switch.scala 41:52:@27077.4]
  assign output_25_11 = io_outValid_11 & _T_65918; // @[Switch.scala 41:38:@27078.4]
  assign _T_65921 = select_12 == 6'h19; // @[Switch.scala 41:52:@27080.4]
  assign output_25_12 = io_outValid_12 & _T_65921; // @[Switch.scala 41:38:@27081.4]
  assign _T_65924 = select_13 == 6'h19; // @[Switch.scala 41:52:@27083.4]
  assign output_25_13 = io_outValid_13 & _T_65924; // @[Switch.scala 41:38:@27084.4]
  assign _T_65927 = select_14 == 6'h19; // @[Switch.scala 41:52:@27086.4]
  assign output_25_14 = io_outValid_14 & _T_65927; // @[Switch.scala 41:38:@27087.4]
  assign _T_65930 = select_15 == 6'h19; // @[Switch.scala 41:52:@27089.4]
  assign output_25_15 = io_outValid_15 & _T_65930; // @[Switch.scala 41:38:@27090.4]
  assign _T_65933 = select_16 == 6'h19; // @[Switch.scala 41:52:@27092.4]
  assign output_25_16 = io_outValid_16 & _T_65933; // @[Switch.scala 41:38:@27093.4]
  assign _T_65936 = select_17 == 6'h19; // @[Switch.scala 41:52:@27095.4]
  assign output_25_17 = io_outValid_17 & _T_65936; // @[Switch.scala 41:38:@27096.4]
  assign _T_65939 = select_18 == 6'h19; // @[Switch.scala 41:52:@27098.4]
  assign output_25_18 = io_outValid_18 & _T_65939; // @[Switch.scala 41:38:@27099.4]
  assign _T_65942 = select_19 == 6'h19; // @[Switch.scala 41:52:@27101.4]
  assign output_25_19 = io_outValid_19 & _T_65942; // @[Switch.scala 41:38:@27102.4]
  assign _T_65945 = select_20 == 6'h19; // @[Switch.scala 41:52:@27104.4]
  assign output_25_20 = io_outValid_20 & _T_65945; // @[Switch.scala 41:38:@27105.4]
  assign _T_65948 = select_21 == 6'h19; // @[Switch.scala 41:52:@27107.4]
  assign output_25_21 = io_outValid_21 & _T_65948; // @[Switch.scala 41:38:@27108.4]
  assign _T_65951 = select_22 == 6'h19; // @[Switch.scala 41:52:@27110.4]
  assign output_25_22 = io_outValid_22 & _T_65951; // @[Switch.scala 41:38:@27111.4]
  assign _T_65954 = select_23 == 6'h19; // @[Switch.scala 41:52:@27113.4]
  assign output_25_23 = io_outValid_23 & _T_65954; // @[Switch.scala 41:38:@27114.4]
  assign _T_65957 = select_24 == 6'h19; // @[Switch.scala 41:52:@27116.4]
  assign output_25_24 = io_outValid_24 & _T_65957; // @[Switch.scala 41:38:@27117.4]
  assign _T_65960 = select_25 == 6'h19; // @[Switch.scala 41:52:@27119.4]
  assign output_25_25 = io_outValid_25 & _T_65960; // @[Switch.scala 41:38:@27120.4]
  assign _T_65963 = select_26 == 6'h19; // @[Switch.scala 41:52:@27122.4]
  assign output_25_26 = io_outValid_26 & _T_65963; // @[Switch.scala 41:38:@27123.4]
  assign _T_65966 = select_27 == 6'h19; // @[Switch.scala 41:52:@27125.4]
  assign output_25_27 = io_outValid_27 & _T_65966; // @[Switch.scala 41:38:@27126.4]
  assign _T_65969 = select_28 == 6'h19; // @[Switch.scala 41:52:@27128.4]
  assign output_25_28 = io_outValid_28 & _T_65969; // @[Switch.scala 41:38:@27129.4]
  assign _T_65972 = select_29 == 6'h19; // @[Switch.scala 41:52:@27131.4]
  assign output_25_29 = io_outValid_29 & _T_65972; // @[Switch.scala 41:38:@27132.4]
  assign _T_65975 = select_30 == 6'h19; // @[Switch.scala 41:52:@27134.4]
  assign output_25_30 = io_outValid_30 & _T_65975; // @[Switch.scala 41:38:@27135.4]
  assign _T_65978 = select_31 == 6'h19; // @[Switch.scala 41:52:@27137.4]
  assign output_25_31 = io_outValid_31 & _T_65978; // @[Switch.scala 41:38:@27138.4]
  assign _T_65981 = select_32 == 6'h19; // @[Switch.scala 41:52:@27140.4]
  assign output_25_32 = io_outValid_32 & _T_65981; // @[Switch.scala 41:38:@27141.4]
  assign _T_65984 = select_33 == 6'h19; // @[Switch.scala 41:52:@27143.4]
  assign output_25_33 = io_outValid_33 & _T_65984; // @[Switch.scala 41:38:@27144.4]
  assign _T_65987 = select_34 == 6'h19; // @[Switch.scala 41:52:@27146.4]
  assign output_25_34 = io_outValid_34 & _T_65987; // @[Switch.scala 41:38:@27147.4]
  assign _T_65990 = select_35 == 6'h19; // @[Switch.scala 41:52:@27149.4]
  assign output_25_35 = io_outValid_35 & _T_65990; // @[Switch.scala 41:38:@27150.4]
  assign _T_65993 = select_36 == 6'h19; // @[Switch.scala 41:52:@27152.4]
  assign output_25_36 = io_outValid_36 & _T_65993; // @[Switch.scala 41:38:@27153.4]
  assign _T_65996 = select_37 == 6'h19; // @[Switch.scala 41:52:@27155.4]
  assign output_25_37 = io_outValid_37 & _T_65996; // @[Switch.scala 41:38:@27156.4]
  assign _T_65999 = select_38 == 6'h19; // @[Switch.scala 41:52:@27158.4]
  assign output_25_38 = io_outValid_38 & _T_65999; // @[Switch.scala 41:38:@27159.4]
  assign _T_66002 = select_39 == 6'h19; // @[Switch.scala 41:52:@27161.4]
  assign output_25_39 = io_outValid_39 & _T_66002; // @[Switch.scala 41:38:@27162.4]
  assign _T_66005 = select_40 == 6'h19; // @[Switch.scala 41:52:@27164.4]
  assign output_25_40 = io_outValid_40 & _T_66005; // @[Switch.scala 41:38:@27165.4]
  assign _T_66008 = select_41 == 6'h19; // @[Switch.scala 41:52:@27167.4]
  assign output_25_41 = io_outValid_41 & _T_66008; // @[Switch.scala 41:38:@27168.4]
  assign _T_66011 = select_42 == 6'h19; // @[Switch.scala 41:52:@27170.4]
  assign output_25_42 = io_outValid_42 & _T_66011; // @[Switch.scala 41:38:@27171.4]
  assign _T_66014 = select_43 == 6'h19; // @[Switch.scala 41:52:@27173.4]
  assign output_25_43 = io_outValid_43 & _T_66014; // @[Switch.scala 41:38:@27174.4]
  assign _T_66017 = select_44 == 6'h19; // @[Switch.scala 41:52:@27176.4]
  assign output_25_44 = io_outValid_44 & _T_66017; // @[Switch.scala 41:38:@27177.4]
  assign _T_66020 = select_45 == 6'h19; // @[Switch.scala 41:52:@27179.4]
  assign output_25_45 = io_outValid_45 & _T_66020; // @[Switch.scala 41:38:@27180.4]
  assign _T_66023 = select_46 == 6'h19; // @[Switch.scala 41:52:@27182.4]
  assign output_25_46 = io_outValid_46 & _T_66023; // @[Switch.scala 41:38:@27183.4]
  assign _T_66026 = select_47 == 6'h19; // @[Switch.scala 41:52:@27185.4]
  assign output_25_47 = io_outValid_47 & _T_66026; // @[Switch.scala 41:38:@27186.4]
  assign _T_66029 = select_48 == 6'h19; // @[Switch.scala 41:52:@27188.4]
  assign output_25_48 = io_outValid_48 & _T_66029; // @[Switch.scala 41:38:@27189.4]
  assign _T_66032 = select_49 == 6'h19; // @[Switch.scala 41:52:@27191.4]
  assign output_25_49 = io_outValid_49 & _T_66032; // @[Switch.scala 41:38:@27192.4]
  assign _T_66035 = select_50 == 6'h19; // @[Switch.scala 41:52:@27194.4]
  assign output_25_50 = io_outValid_50 & _T_66035; // @[Switch.scala 41:38:@27195.4]
  assign _T_66038 = select_51 == 6'h19; // @[Switch.scala 41:52:@27197.4]
  assign output_25_51 = io_outValid_51 & _T_66038; // @[Switch.scala 41:38:@27198.4]
  assign _T_66041 = select_52 == 6'h19; // @[Switch.scala 41:52:@27200.4]
  assign output_25_52 = io_outValid_52 & _T_66041; // @[Switch.scala 41:38:@27201.4]
  assign _T_66044 = select_53 == 6'h19; // @[Switch.scala 41:52:@27203.4]
  assign output_25_53 = io_outValid_53 & _T_66044; // @[Switch.scala 41:38:@27204.4]
  assign _T_66047 = select_54 == 6'h19; // @[Switch.scala 41:52:@27206.4]
  assign output_25_54 = io_outValid_54 & _T_66047; // @[Switch.scala 41:38:@27207.4]
  assign _T_66050 = select_55 == 6'h19; // @[Switch.scala 41:52:@27209.4]
  assign output_25_55 = io_outValid_55 & _T_66050; // @[Switch.scala 41:38:@27210.4]
  assign _T_66053 = select_56 == 6'h19; // @[Switch.scala 41:52:@27212.4]
  assign output_25_56 = io_outValid_56 & _T_66053; // @[Switch.scala 41:38:@27213.4]
  assign _T_66056 = select_57 == 6'h19; // @[Switch.scala 41:52:@27215.4]
  assign output_25_57 = io_outValid_57 & _T_66056; // @[Switch.scala 41:38:@27216.4]
  assign _T_66059 = select_58 == 6'h19; // @[Switch.scala 41:52:@27218.4]
  assign output_25_58 = io_outValid_58 & _T_66059; // @[Switch.scala 41:38:@27219.4]
  assign _T_66062 = select_59 == 6'h19; // @[Switch.scala 41:52:@27221.4]
  assign output_25_59 = io_outValid_59 & _T_66062; // @[Switch.scala 41:38:@27222.4]
  assign _T_66065 = select_60 == 6'h19; // @[Switch.scala 41:52:@27224.4]
  assign output_25_60 = io_outValid_60 & _T_66065; // @[Switch.scala 41:38:@27225.4]
  assign _T_66068 = select_61 == 6'h19; // @[Switch.scala 41:52:@27227.4]
  assign output_25_61 = io_outValid_61 & _T_66068; // @[Switch.scala 41:38:@27228.4]
  assign _T_66071 = select_62 == 6'h19; // @[Switch.scala 41:52:@27230.4]
  assign output_25_62 = io_outValid_62 & _T_66071; // @[Switch.scala 41:38:@27231.4]
  assign _T_66074 = select_63 == 6'h19; // @[Switch.scala 41:52:@27233.4]
  assign output_25_63 = io_outValid_63 & _T_66074; // @[Switch.scala 41:38:@27234.4]
  assign _T_66082 = {output_25_7,output_25_6,output_25_5,output_25_4,output_25_3,output_25_2,output_25_1,output_25_0}; // @[Switch.scala 43:31:@27242.4]
  assign _T_66090 = {output_25_15,output_25_14,output_25_13,output_25_12,output_25_11,output_25_10,output_25_9,output_25_8,_T_66082}; // @[Switch.scala 43:31:@27250.4]
  assign _T_66097 = {output_25_23,output_25_22,output_25_21,output_25_20,output_25_19,output_25_18,output_25_17,output_25_16}; // @[Switch.scala 43:31:@27257.4]
  assign _T_66106 = {output_25_31,output_25_30,output_25_29,output_25_28,output_25_27,output_25_26,output_25_25,output_25_24,_T_66097,_T_66090}; // @[Switch.scala 43:31:@27266.4]
  assign _T_66113 = {output_25_39,output_25_38,output_25_37,output_25_36,output_25_35,output_25_34,output_25_33,output_25_32}; // @[Switch.scala 43:31:@27273.4]
  assign _T_66121 = {output_25_47,output_25_46,output_25_45,output_25_44,output_25_43,output_25_42,output_25_41,output_25_40,_T_66113}; // @[Switch.scala 43:31:@27281.4]
  assign _T_66128 = {output_25_55,output_25_54,output_25_53,output_25_52,output_25_51,output_25_50,output_25_49,output_25_48}; // @[Switch.scala 43:31:@27288.4]
  assign _T_66137 = {output_25_63,output_25_62,output_25_61,output_25_60,output_25_59,output_25_58,output_25_57,output_25_56,_T_66128,_T_66121}; // @[Switch.scala 43:31:@27297.4]
  assign _T_66138 = {_T_66137,_T_66106}; // @[Switch.scala 43:31:@27298.4]
  assign _T_66142 = select_0 == 6'h1a; // @[Switch.scala 41:52:@27301.4]
  assign output_26_0 = io_outValid_0 & _T_66142; // @[Switch.scala 41:38:@27302.4]
  assign _T_66145 = select_1 == 6'h1a; // @[Switch.scala 41:52:@27304.4]
  assign output_26_1 = io_outValid_1 & _T_66145; // @[Switch.scala 41:38:@27305.4]
  assign _T_66148 = select_2 == 6'h1a; // @[Switch.scala 41:52:@27307.4]
  assign output_26_2 = io_outValid_2 & _T_66148; // @[Switch.scala 41:38:@27308.4]
  assign _T_66151 = select_3 == 6'h1a; // @[Switch.scala 41:52:@27310.4]
  assign output_26_3 = io_outValid_3 & _T_66151; // @[Switch.scala 41:38:@27311.4]
  assign _T_66154 = select_4 == 6'h1a; // @[Switch.scala 41:52:@27313.4]
  assign output_26_4 = io_outValid_4 & _T_66154; // @[Switch.scala 41:38:@27314.4]
  assign _T_66157 = select_5 == 6'h1a; // @[Switch.scala 41:52:@27316.4]
  assign output_26_5 = io_outValid_5 & _T_66157; // @[Switch.scala 41:38:@27317.4]
  assign _T_66160 = select_6 == 6'h1a; // @[Switch.scala 41:52:@27319.4]
  assign output_26_6 = io_outValid_6 & _T_66160; // @[Switch.scala 41:38:@27320.4]
  assign _T_66163 = select_7 == 6'h1a; // @[Switch.scala 41:52:@27322.4]
  assign output_26_7 = io_outValid_7 & _T_66163; // @[Switch.scala 41:38:@27323.4]
  assign _T_66166 = select_8 == 6'h1a; // @[Switch.scala 41:52:@27325.4]
  assign output_26_8 = io_outValid_8 & _T_66166; // @[Switch.scala 41:38:@27326.4]
  assign _T_66169 = select_9 == 6'h1a; // @[Switch.scala 41:52:@27328.4]
  assign output_26_9 = io_outValid_9 & _T_66169; // @[Switch.scala 41:38:@27329.4]
  assign _T_66172 = select_10 == 6'h1a; // @[Switch.scala 41:52:@27331.4]
  assign output_26_10 = io_outValid_10 & _T_66172; // @[Switch.scala 41:38:@27332.4]
  assign _T_66175 = select_11 == 6'h1a; // @[Switch.scala 41:52:@27334.4]
  assign output_26_11 = io_outValid_11 & _T_66175; // @[Switch.scala 41:38:@27335.4]
  assign _T_66178 = select_12 == 6'h1a; // @[Switch.scala 41:52:@27337.4]
  assign output_26_12 = io_outValid_12 & _T_66178; // @[Switch.scala 41:38:@27338.4]
  assign _T_66181 = select_13 == 6'h1a; // @[Switch.scala 41:52:@27340.4]
  assign output_26_13 = io_outValid_13 & _T_66181; // @[Switch.scala 41:38:@27341.4]
  assign _T_66184 = select_14 == 6'h1a; // @[Switch.scala 41:52:@27343.4]
  assign output_26_14 = io_outValid_14 & _T_66184; // @[Switch.scala 41:38:@27344.4]
  assign _T_66187 = select_15 == 6'h1a; // @[Switch.scala 41:52:@27346.4]
  assign output_26_15 = io_outValid_15 & _T_66187; // @[Switch.scala 41:38:@27347.4]
  assign _T_66190 = select_16 == 6'h1a; // @[Switch.scala 41:52:@27349.4]
  assign output_26_16 = io_outValid_16 & _T_66190; // @[Switch.scala 41:38:@27350.4]
  assign _T_66193 = select_17 == 6'h1a; // @[Switch.scala 41:52:@27352.4]
  assign output_26_17 = io_outValid_17 & _T_66193; // @[Switch.scala 41:38:@27353.4]
  assign _T_66196 = select_18 == 6'h1a; // @[Switch.scala 41:52:@27355.4]
  assign output_26_18 = io_outValid_18 & _T_66196; // @[Switch.scala 41:38:@27356.4]
  assign _T_66199 = select_19 == 6'h1a; // @[Switch.scala 41:52:@27358.4]
  assign output_26_19 = io_outValid_19 & _T_66199; // @[Switch.scala 41:38:@27359.4]
  assign _T_66202 = select_20 == 6'h1a; // @[Switch.scala 41:52:@27361.4]
  assign output_26_20 = io_outValid_20 & _T_66202; // @[Switch.scala 41:38:@27362.4]
  assign _T_66205 = select_21 == 6'h1a; // @[Switch.scala 41:52:@27364.4]
  assign output_26_21 = io_outValid_21 & _T_66205; // @[Switch.scala 41:38:@27365.4]
  assign _T_66208 = select_22 == 6'h1a; // @[Switch.scala 41:52:@27367.4]
  assign output_26_22 = io_outValid_22 & _T_66208; // @[Switch.scala 41:38:@27368.4]
  assign _T_66211 = select_23 == 6'h1a; // @[Switch.scala 41:52:@27370.4]
  assign output_26_23 = io_outValid_23 & _T_66211; // @[Switch.scala 41:38:@27371.4]
  assign _T_66214 = select_24 == 6'h1a; // @[Switch.scala 41:52:@27373.4]
  assign output_26_24 = io_outValid_24 & _T_66214; // @[Switch.scala 41:38:@27374.4]
  assign _T_66217 = select_25 == 6'h1a; // @[Switch.scala 41:52:@27376.4]
  assign output_26_25 = io_outValid_25 & _T_66217; // @[Switch.scala 41:38:@27377.4]
  assign _T_66220 = select_26 == 6'h1a; // @[Switch.scala 41:52:@27379.4]
  assign output_26_26 = io_outValid_26 & _T_66220; // @[Switch.scala 41:38:@27380.4]
  assign _T_66223 = select_27 == 6'h1a; // @[Switch.scala 41:52:@27382.4]
  assign output_26_27 = io_outValid_27 & _T_66223; // @[Switch.scala 41:38:@27383.4]
  assign _T_66226 = select_28 == 6'h1a; // @[Switch.scala 41:52:@27385.4]
  assign output_26_28 = io_outValid_28 & _T_66226; // @[Switch.scala 41:38:@27386.4]
  assign _T_66229 = select_29 == 6'h1a; // @[Switch.scala 41:52:@27388.4]
  assign output_26_29 = io_outValid_29 & _T_66229; // @[Switch.scala 41:38:@27389.4]
  assign _T_66232 = select_30 == 6'h1a; // @[Switch.scala 41:52:@27391.4]
  assign output_26_30 = io_outValid_30 & _T_66232; // @[Switch.scala 41:38:@27392.4]
  assign _T_66235 = select_31 == 6'h1a; // @[Switch.scala 41:52:@27394.4]
  assign output_26_31 = io_outValid_31 & _T_66235; // @[Switch.scala 41:38:@27395.4]
  assign _T_66238 = select_32 == 6'h1a; // @[Switch.scala 41:52:@27397.4]
  assign output_26_32 = io_outValid_32 & _T_66238; // @[Switch.scala 41:38:@27398.4]
  assign _T_66241 = select_33 == 6'h1a; // @[Switch.scala 41:52:@27400.4]
  assign output_26_33 = io_outValid_33 & _T_66241; // @[Switch.scala 41:38:@27401.4]
  assign _T_66244 = select_34 == 6'h1a; // @[Switch.scala 41:52:@27403.4]
  assign output_26_34 = io_outValid_34 & _T_66244; // @[Switch.scala 41:38:@27404.4]
  assign _T_66247 = select_35 == 6'h1a; // @[Switch.scala 41:52:@27406.4]
  assign output_26_35 = io_outValid_35 & _T_66247; // @[Switch.scala 41:38:@27407.4]
  assign _T_66250 = select_36 == 6'h1a; // @[Switch.scala 41:52:@27409.4]
  assign output_26_36 = io_outValid_36 & _T_66250; // @[Switch.scala 41:38:@27410.4]
  assign _T_66253 = select_37 == 6'h1a; // @[Switch.scala 41:52:@27412.4]
  assign output_26_37 = io_outValid_37 & _T_66253; // @[Switch.scala 41:38:@27413.4]
  assign _T_66256 = select_38 == 6'h1a; // @[Switch.scala 41:52:@27415.4]
  assign output_26_38 = io_outValid_38 & _T_66256; // @[Switch.scala 41:38:@27416.4]
  assign _T_66259 = select_39 == 6'h1a; // @[Switch.scala 41:52:@27418.4]
  assign output_26_39 = io_outValid_39 & _T_66259; // @[Switch.scala 41:38:@27419.4]
  assign _T_66262 = select_40 == 6'h1a; // @[Switch.scala 41:52:@27421.4]
  assign output_26_40 = io_outValid_40 & _T_66262; // @[Switch.scala 41:38:@27422.4]
  assign _T_66265 = select_41 == 6'h1a; // @[Switch.scala 41:52:@27424.4]
  assign output_26_41 = io_outValid_41 & _T_66265; // @[Switch.scala 41:38:@27425.4]
  assign _T_66268 = select_42 == 6'h1a; // @[Switch.scala 41:52:@27427.4]
  assign output_26_42 = io_outValid_42 & _T_66268; // @[Switch.scala 41:38:@27428.4]
  assign _T_66271 = select_43 == 6'h1a; // @[Switch.scala 41:52:@27430.4]
  assign output_26_43 = io_outValid_43 & _T_66271; // @[Switch.scala 41:38:@27431.4]
  assign _T_66274 = select_44 == 6'h1a; // @[Switch.scala 41:52:@27433.4]
  assign output_26_44 = io_outValid_44 & _T_66274; // @[Switch.scala 41:38:@27434.4]
  assign _T_66277 = select_45 == 6'h1a; // @[Switch.scala 41:52:@27436.4]
  assign output_26_45 = io_outValid_45 & _T_66277; // @[Switch.scala 41:38:@27437.4]
  assign _T_66280 = select_46 == 6'h1a; // @[Switch.scala 41:52:@27439.4]
  assign output_26_46 = io_outValid_46 & _T_66280; // @[Switch.scala 41:38:@27440.4]
  assign _T_66283 = select_47 == 6'h1a; // @[Switch.scala 41:52:@27442.4]
  assign output_26_47 = io_outValid_47 & _T_66283; // @[Switch.scala 41:38:@27443.4]
  assign _T_66286 = select_48 == 6'h1a; // @[Switch.scala 41:52:@27445.4]
  assign output_26_48 = io_outValid_48 & _T_66286; // @[Switch.scala 41:38:@27446.4]
  assign _T_66289 = select_49 == 6'h1a; // @[Switch.scala 41:52:@27448.4]
  assign output_26_49 = io_outValid_49 & _T_66289; // @[Switch.scala 41:38:@27449.4]
  assign _T_66292 = select_50 == 6'h1a; // @[Switch.scala 41:52:@27451.4]
  assign output_26_50 = io_outValid_50 & _T_66292; // @[Switch.scala 41:38:@27452.4]
  assign _T_66295 = select_51 == 6'h1a; // @[Switch.scala 41:52:@27454.4]
  assign output_26_51 = io_outValid_51 & _T_66295; // @[Switch.scala 41:38:@27455.4]
  assign _T_66298 = select_52 == 6'h1a; // @[Switch.scala 41:52:@27457.4]
  assign output_26_52 = io_outValid_52 & _T_66298; // @[Switch.scala 41:38:@27458.4]
  assign _T_66301 = select_53 == 6'h1a; // @[Switch.scala 41:52:@27460.4]
  assign output_26_53 = io_outValid_53 & _T_66301; // @[Switch.scala 41:38:@27461.4]
  assign _T_66304 = select_54 == 6'h1a; // @[Switch.scala 41:52:@27463.4]
  assign output_26_54 = io_outValid_54 & _T_66304; // @[Switch.scala 41:38:@27464.4]
  assign _T_66307 = select_55 == 6'h1a; // @[Switch.scala 41:52:@27466.4]
  assign output_26_55 = io_outValid_55 & _T_66307; // @[Switch.scala 41:38:@27467.4]
  assign _T_66310 = select_56 == 6'h1a; // @[Switch.scala 41:52:@27469.4]
  assign output_26_56 = io_outValid_56 & _T_66310; // @[Switch.scala 41:38:@27470.4]
  assign _T_66313 = select_57 == 6'h1a; // @[Switch.scala 41:52:@27472.4]
  assign output_26_57 = io_outValid_57 & _T_66313; // @[Switch.scala 41:38:@27473.4]
  assign _T_66316 = select_58 == 6'h1a; // @[Switch.scala 41:52:@27475.4]
  assign output_26_58 = io_outValid_58 & _T_66316; // @[Switch.scala 41:38:@27476.4]
  assign _T_66319 = select_59 == 6'h1a; // @[Switch.scala 41:52:@27478.4]
  assign output_26_59 = io_outValid_59 & _T_66319; // @[Switch.scala 41:38:@27479.4]
  assign _T_66322 = select_60 == 6'h1a; // @[Switch.scala 41:52:@27481.4]
  assign output_26_60 = io_outValid_60 & _T_66322; // @[Switch.scala 41:38:@27482.4]
  assign _T_66325 = select_61 == 6'h1a; // @[Switch.scala 41:52:@27484.4]
  assign output_26_61 = io_outValid_61 & _T_66325; // @[Switch.scala 41:38:@27485.4]
  assign _T_66328 = select_62 == 6'h1a; // @[Switch.scala 41:52:@27487.4]
  assign output_26_62 = io_outValid_62 & _T_66328; // @[Switch.scala 41:38:@27488.4]
  assign _T_66331 = select_63 == 6'h1a; // @[Switch.scala 41:52:@27490.4]
  assign output_26_63 = io_outValid_63 & _T_66331; // @[Switch.scala 41:38:@27491.4]
  assign _T_66339 = {output_26_7,output_26_6,output_26_5,output_26_4,output_26_3,output_26_2,output_26_1,output_26_0}; // @[Switch.scala 43:31:@27499.4]
  assign _T_66347 = {output_26_15,output_26_14,output_26_13,output_26_12,output_26_11,output_26_10,output_26_9,output_26_8,_T_66339}; // @[Switch.scala 43:31:@27507.4]
  assign _T_66354 = {output_26_23,output_26_22,output_26_21,output_26_20,output_26_19,output_26_18,output_26_17,output_26_16}; // @[Switch.scala 43:31:@27514.4]
  assign _T_66363 = {output_26_31,output_26_30,output_26_29,output_26_28,output_26_27,output_26_26,output_26_25,output_26_24,_T_66354,_T_66347}; // @[Switch.scala 43:31:@27523.4]
  assign _T_66370 = {output_26_39,output_26_38,output_26_37,output_26_36,output_26_35,output_26_34,output_26_33,output_26_32}; // @[Switch.scala 43:31:@27530.4]
  assign _T_66378 = {output_26_47,output_26_46,output_26_45,output_26_44,output_26_43,output_26_42,output_26_41,output_26_40,_T_66370}; // @[Switch.scala 43:31:@27538.4]
  assign _T_66385 = {output_26_55,output_26_54,output_26_53,output_26_52,output_26_51,output_26_50,output_26_49,output_26_48}; // @[Switch.scala 43:31:@27545.4]
  assign _T_66394 = {output_26_63,output_26_62,output_26_61,output_26_60,output_26_59,output_26_58,output_26_57,output_26_56,_T_66385,_T_66378}; // @[Switch.scala 43:31:@27554.4]
  assign _T_66395 = {_T_66394,_T_66363}; // @[Switch.scala 43:31:@27555.4]
  assign _T_66399 = select_0 == 6'h1b; // @[Switch.scala 41:52:@27558.4]
  assign output_27_0 = io_outValid_0 & _T_66399; // @[Switch.scala 41:38:@27559.4]
  assign _T_66402 = select_1 == 6'h1b; // @[Switch.scala 41:52:@27561.4]
  assign output_27_1 = io_outValid_1 & _T_66402; // @[Switch.scala 41:38:@27562.4]
  assign _T_66405 = select_2 == 6'h1b; // @[Switch.scala 41:52:@27564.4]
  assign output_27_2 = io_outValid_2 & _T_66405; // @[Switch.scala 41:38:@27565.4]
  assign _T_66408 = select_3 == 6'h1b; // @[Switch.scala 41:52:@27567.4]
  assign output_27_3 = io_outValid_3 & _T_66408; // @[Switch.scala 41:38:@27568.4]
  assign _T_66411 = select_4 == 6'h1b; // @[Switch.scala 41:52:@27570.4]
  assign output_27_4 = io_outValid_4 & _T_66411; // @[Switch.scala 41:38:@27571.4]
  assign _T_66414 = select_5 == 6'h1b; // @[Switch.scala 41:52:@27573.4]
  assign output_27_5 = io_outValid_5 & _T_66414; // @[Switch.scala 41:38:@27574.4]
  assign _T_66417 = select_6 == 6'h1b; // @[Switch.scala 41:52:@27576.4]
  assign output_27_6 = io_outValid_6 & _T_66417; // @[Switch.scala 41:38:@27577.4]
  assign _T_66420 = select_7 == 6'h1b; // @[Switch.scala 41:52:@27579.4]
  assign output_27_7 = io_outValid_7 & _T_66420; // @[Switch.scala 41:38:@27580.4]
  assign _T_66423 = select_8 == 6'h1b; // @[Switch.scala 41:52:@27582.4]
  assign output_27_8 = io_outValid_8 & _T_66423; // @[Switch.scala 41:38:@27583.4]
  assign _T_66426 = select_9 == 6'h1b; // @[Switch.scala 41:52:@27585.4]
  assign output_27_9 = io_outValid_9 & _T_66426; // @[Switch.scala 41:38:@27586.4]
  assign _T_66429 = select_10 == 6'h1b; // @[Switch.scala 41:52:@27588.4]
  assign output_27_10 = io_outValid_10 & _T_66429; // @[Switch.scala 41:38:@27589.4]
  assign _T_66432 = select_11 == 6'h1b; // @[Switch.scala 41:52:@27591.4]
  assign output_27_11 = io_outValid_11 & _T_66432; // @[Switch.scala 41:38:@27592.4]
  assign _T_66435 = select_12 == 6'h1b; // @[Switch.scala 41:52:@27594.4]
  assign output_27_12 = io_outValid_12 & _T_66435; // @[Switch.scala 41:38:@27595.4]
  assign _T_66438 = select_13 == 6'h1b; // @[Switch.scala 41:52:@27597.4]
  assign output_27_13 = io_outValid_13 & _T_66438; // @[Switch.scala 41:38:@27598.4]
  assign _T_66441 = select_14 == 6'h1b; // @[Switch.scala 41:52:@27600.4]
  assign output_27_14 = io_outValid_14 & _T_66441; // @[Switch.scala 41:38:@27601.4]
  assign _T_66444 = select_15 == 6'h1b; // @[Switch.scala 41:52:@27603.4]
  assign output_27_15 = io_outValid_15 & _T_66444; // @[Switch.scala 41:38:@27604.4]
  assign _T_66447 = select_16 == 6'h1b; // @[Switch.scala 41:52:@27606.4]
  assign output_27_16 = io_outValid_16 & _T_66447; // @[Switch.scala 41:38:@27607.4]
  assign _T_66450 = select_17 == 6'h1b; // @[Switch.scala 41:52:@27609.4]
  assign output_27_17 = io_outValid_17 & _T_66450; // @[Switch.scala 41:38:@27610.4]
  assign _T_66453 = select_18 == 6'h1b; // @[Switch.scala 41:52:@27612.4]
  assign output_27_18 = io_outValid_18 & _T_66453; // @[Switch.scala 41:38:@27613.4]
  assign _T_66456 = select_19 == 6'h1b; // @[Switch.scala 41:52:@27615.4]
  assign output_27_19 = io_outValid_19 & _T_66456; // @[Switch.scala 41:38:@27616.4]
  assign _T_66459 = select_20 == 6'h1b; // @[Switch.scala 41:52:@27618.4]
  assign output_27_20 = io_outValid_20 & _T_66459; // @[Switch.scala 41:38:@27619.4]
  assign _T_66462 = select_21 == 6'h1b; // @[Switch.scala 41:52:@27621.4]
  assign output_27_21 = io_outValid_21 & _T_66462; // @[Switch.scala 41:38:@27622.4]
  assign _T_66465 = select_22 == 6'h1b; // @[Switch.scala 41:52:@27624.4]
  assign output_27_22 = io_outValid_22 & _T_66465; // @[Switch.scala 41:38:@27625.4]
  assign _T_66468 = select_23 == 6'h1b; // @[Switch.scala 41:52:@27627.4]
  assign output_27_23 = io_outValid_23 & _T_66468; // @[Switch.scala 41:38:@27628.4]
  assign _T_66471 = select_24 == 6'h1b; // @[Switch.scala 41:52:@27630.4]
  assign output_27_24 = io_outValid_24 & _T_66471; // @[Switch.scala 41:38:@27631.4]
  assign _T_66474 = select_25 == 6'h1b; // @[Switch.scala 41:52:@27633.4]
  assign output_27_25 = io_outValid_25 & _T_66474; // @[Switch.scala 41:38:@27634.4]
  assign _T_66477 = select_26 == 6'h1b; // @[Switch.scala 41:52:@27636.4]
  assign output_27_26 = io_outValid_26 & _T_66477; // @[Switch.scala 41:38:@27637.4]
  assign _T_66480 = select_27 == 6'h1b; // @[Switch.scala 41:52:@27639.4]
  assign output_27_27 = io_outValid_27 & _T_66480; // @[Switch.scala 41:38:@27640.4]
  assign _T_66483 = select_28 == 6'h1b; // @[Switch.scala 41:52:@27642.4]
  assign output_27_28 = io_outValid_28 & _T_66483; // @[Switch.scala 41:38:@27643.4]
  assign _T_66486 = select_29 == 6'h1b; // @[Switch.scala 41:52:@27645.4]
  assign output_27_29 = io_outValid_29 & _T_66486; // @[Switch.scala 41:38:@27646.4]
  assign _T_66489 = select_30 == 6'h1b; // @[Switch.scala 41:52:@27648.4]
  assign output_27_30 = io_outValid_30 & _T_66489; // @[Switch.scala 41:38:@27649.4]
  assign _T_66492 = select_31 == 6'h1b; // @[Switch.scala 41:52:@27651.4]
  assign output_27_31 = io_outValid_31 & _T_66492; // @[Switch.scala 41:38:@27652.4]
  assign _T_66495 = select_32 == 6'h1b; // @[Switch.scala 41:52:@27654.4]
  assign output_27_32 = io_outValid_32 & _T_66495; // @[Switch.scala 41:38:@27655.4]
  assign _T_66498 = select_33 == 6'h1b; // @[Switch.scala 41:52:@27657.4]
  assign output_27_33 = io_outValid_33 & _T_66498; // @[Switch.scala 41:38:@27658.4]
  assign _T_66501 = select_34 == 6'h1b; // @[Switch.scala 41:52:@27660.4]
  assign output_27_34 = io_outValid_34 & _T_66501; // @[Switch.scala 41:38:@27661.4]
  assign _T_66504 = select_35 == 6'h1b; // @[Switch.scala 41:52:@27663.4]
  assign output_27_35 = io_outValid_35 & _T_66504; // @[Switch.scala 41:38:@27664.4]
  assign _T_66507 = select_36 == 6'h1b; // @[Switch.scala 41:52:@27666.4]
  assign output_27_36 = io_outValid_36 & _T_66507; // @[Switch.scala 41:38:@27667.4]
  assign _T_66510 = select_37 == 6'h1b; // @[Switch.scala 41:52:@27669.4]
  assign output_27_37 = io_outValid_37 & _T_66510; // @[Switch.scala 41:38:@27670.4]
  assign _T_66513 = select_38 == 6'h1b; // @[Switch.scala 41:52:@27672.4]
  assign output_27_38 = io_outValid_38 & _T_66513; // @[Switch.scala 41:38:@27673.4]
  assign _T_66516 = select_39 == 6'h1b; // @[Switch.scala 41:52:@27675.4]
  assign output_27_39 = io_outValid_39 & _T_66516; // @[Switch.scala 41:38:@27676.4]
  assign _T_66519 = select_40 == 6'h1b; // @[Switch.scala 41:52:@27678.4]
  assign output_27_40 = io_outValid_40 & _T_66519; // @[Switch.scala 41:38:@27679.4]
  assign _T_66522 = select_41 == 6'h1b; // @[Switch.scala 41:52:@27681.4]
  assign output_27_41 = io_outValid_41 & _T_66522; // @[Switch.scala 41:38:@27682.4]
  assign _T_66525 = select_42 == 6'h1b; // @[Switch.scala 41:52:@27684.4]
  assign output_27_42 = io_outValid_42 & _T_66525; // @[Switch.scala 41:38:@27685.4]
  assign _T_66528 = select_43 == 6'h1b; // @[Switch.scala 41:52:@27687.4]
  assign output_27_43 = io_outValid_43 & _T_66528; // @[Switch.scala 41:38:@27688.4]
  assign _T_66531 = select_44 == 6'h1b; // @[Switch.scala 41:52:@27690.4]
  assign output_27_44 = io_outValid_44 & _T_66531; // @[Switch.scala 41:38:@27691.4]
  assign _T_66534 = select_45 == 6'h1b; // @[Switch.scala 41:52:@27693.4]
  assign output_27_45 = io_outValid_45 & _T_66534; // @[Switch.scala 41:38:@27694.4]
  assign _T_66537 = select_46 == 6'h1b; // @[Switch.scala 41:52:@27696.4]
  assign output_27_46 = io_outValid_46 & _T_66537; // @[Switch.scala 41:38:@27697.4]
  assign _T_66540 = select_47 == 6'h1b; // @[Switch.scala 41:52:@27699.4]
  assign output_27_47 = io_outValid_47 & _T_66540; // @[Switch.scala 41:38:@27700.4]
  assign _T_66543 = select_48 == 6'h1b; // @[Switch.scala 41:52:@27702.4]
  assign output_27_48 = io_outValid_48 & _T_66543; // @[Switch.scala 41:38:@27703.4]
  assign _T_66546 = select_49 == 6'h1b; // @[Switch.scala 41:52:@27705.4]
  assign output_27_49 = io_outValid_49 & _T_66546; // @[Switch.scala 41:38:@27706.4]
  assign _T_66549 = select_50 == 6'h1b; // @[Switch.scala 41:52:@27708.4]
  assign output_27_50 = io_outValid_50 & _T_66549; // @[Switch.scala 41:38:@27709.4]
  assign _T_66552 = select_51 == 6'h1b; // @[Switch.scala 41:52:@27711.4]
  assign output_27_51 = io_outValid_51 & _T_66552; // @[Switch.scala 41:38:@27712.4]
  assign _T_66555 = select_52 == 6'h1b; // @[Switch.scala 41:52:@27714.4]
  assign output_27_52 = io_outValid_52 & _T_66555; // @[Switch.scala 41:38:@27715.4]
  assign _T_66558 = select_53 == 6'h1b; // @[Switch.scala 41:52:@27717.4]
  assign output_27_53 = io_outValid_53 & _T_66558; // @[Switch.scala 41:38:@27718.4]
  assign _T_66561 = select_54 == 6'h1b; // @[Switch.scala 41:52:@27720.4]
  assign output_27_54 = io_outValid_54 & _T_66561; // @[Switch.scala 41:38:@27721.4]
  assign _T_66564 = select_55 == 6'h1b; // @[Switch.scala 41:52:@27723.4]
  assign output_27_55 = io_outValid_55 & _T_66564; // @[Switch.scala 41:38:@27724.4]
  assign _T_66567 = select_56 == 6'h1b; // @[Switch.scala 41:52:@27726.4]
  assign output_27_56 = io_outValid_56 & _T_66567; // @[Switch.scala 41:38:@27727.4]
  assign _T_66570 = select_57 == 6'h1b; // @[Switch.scala 41:52:@27729.4]
  assign output_27_57 = io_outValid_57 & _T_66570; // @[Switch.scala 41:38:@27730.4]
  assign _T_66573 = select_58 == 6'h1b; // @[Switch.scala 41:52:@27732.4]
  assign output_27_58 = io_outValid_58 & _T_66573; // @[Switch.scala 41:38:@27733.4]
  assign _T_66576 = select_59 == 6'h1b; // @[Switch.scala 41:52:@27735.4]
  assign output_27_59 = io_outValid_59 & _T_66576; // @[Switch.scala 41:38:@27736.4]
  assign _T_66579 = select_60 == 6'h1b; // @[Switch.scala 41:52:@27738.4]
  assign output_27_60 = io_outValid_60 & _T_66579; // @[Switch.scala 41:38:@27739.4]
  assign _T_66582 = select_61 == 6'h1b; // @[Switch.scala 41:52:@27741.4]
  assign output_27_61 = io_outValid_61 & _T_66582; // @[Switch.scala 41:38:@27742.4]
  assign _T_66585 = select_62 == 6'h1b; // @[Switch.scala 41:52:@27744.4]
  assign output_27_62 = io_outValid_62 & _T_66585; // @[Switch.scala 41:38:@27745.4]
  assign _T_66588 = select_63 == 6'h1b; // @[Switch.scala 41:52:@27747.4]
  assign output_27_63 = io_outValid_63 & _T_66588; // @[Switch.scala 41:38:@27748.4]
  assign _T_66596 = {output_27_7,output_27_6,output_27_5,output_27_4,output_27_3,output_27_2,output_27_1,output_27_0}; // @[Switch.scala 43:31:@27756.4]
  assign _T_66604 = {output_27_15,output_27_14,output_27_13,output_27_12,output_27_11,output_27_10,output_27_9,output_27_8,_T_66596}; // @[Switch.scala 43:31:@27764.4]
  assign _T_66611 = {output_27_23,output_27_22,output_27_21,output_27_20,output_27_19,output_27_18,output_27_17,output_27_16}; // @[Switch.scala 43:31:@27771.4]
  assign _T_66620 = {output_27_31,output_27_30,output_27_29,output_27_28,output_27_27,output_27_26,output_27_25,output_27_24,_T_66611,_T_66604}; // @[Switch.scala 43:31:@27780.4]
  assign _T_66627 = {output_27_39,output_27_38,output_27_37,output_27_36,output_27_35,output_27_34,output_27_33,output_27_32}; // @[Switch.scala 43:31:@27787.4]
  assign _T_66635 = {output_27_47,output_27_46,output_27_45,output_27_44,output_27_43,output_27_42,output_27_41,output_27_40,_T_66627}; // @[Switch.scala 43:31:@27795.4]
  assign _T_66642 = {output_27_55,output_27_54,output_27_53,output_27_52,output_27_51,output_27_50,output_27_49,output_27_48}; // @[Switch.scala 43:31:@27802.4]
  assign _T_66651 = {output_27_63,output_27_62,output_27_61,output_27_60,output_27_59,output_27_58,output_27_57,output_27_56,_T_66642,_T_66635}; // @[Switch.scala 43:31:@27811.4]
  assign _T_66652 = {_T_66651,_T_66620}; // @[Switch.scala 43:31:@27812.4]
  assign _T_66656 = select_0 == 6'h1c; // @[Switch.scala 41:52:@27815.4]
  assign output_28_0 = io_outValid_0 & _T_66656; // @[Switch.scala 41:38:@27816.4]
  assign _T_66659 = select_1 == 6'h1c; // @[Switch.scala 41:52:@27818.4]
  assign output_28_1 = io_outValid_1 & _T_66659; // @[Switch.scala 41:38:@27819.4]
  assign _T_66662 = select_2 == 6'h1c; // @[Switch.scala 41:52:@27821.4]
  assign output_28_2 = io_outValid_2 & _T_66662; // @[Switch.scala 41:38:@27822.4]
  assign _T_66665 = select_3 == 6'h1c; // @[Switch.scala 41:52:@27824.4]
  assign output_28_3 = io_outValid_3 & _T_66665; // @[Switch.scala 41:38:@27825.4]
  assign _T_66668 = select_4 == 6'h1c; // @[Switch.scala 41:52:@27827.4]
  assign output_28_4 = io_outValid_4 & _T_66668; // @[Switch.scala 41:38:@27828.4]
  assign _T_66671 = select_5 == 6'h1c; // @[Switch.scala 41:52:@27830.4]
  assign output_28_5 = io_outValid_5 & _T_66671; // @[Switch.scala 41:38:@27831.4]
  assign _T_66674 = select_6 == 6'h1c; // @[Switch.scala 41:52:@27833.4]
  assign output_28_6 = io_outValid_6 & _T_66674; // @[Switch.scala 41:38:@27834.4]
  assign _T_66677 = select_7 == 6'h1c; // @[Switch.scala 41:52:@27836.4]
  assign output_28_7 = io_outValid_7 & _T_66677; // @[Switch.scala 41:38:@27837.4]
  assign _T_66680 = select_8 == 6'h1c; // @[Switch.scala 41:52:@27839.4]
  assign output_28_8 = io_outValid_8 & _T_66680; // @[Switch.scala 41:38:@27840.4]
  assign _T_66683 = select_9 == 6'h1c; // @[Switch.scala 41:52:@27842.4]
  assign output_28_9 = io_outValid_9 & _T_66683; // @[Switch.scala 41:38:@27843.4]
  assign _T_66686 = select_10 == 6'h1c; // @[Switch.scala 41:52:@27845.4]
  assign output_28_10 = io_outValid_10 & _T_66686; // @[Switch.scala 41:38:@27846.4]
  assign _T_66689 = select_11 == 6'h1c; // @[Switch.scala 41:52:@27848.4]
  assign output_28_11 = io_outValid_11 & _T_66689; // @[Switch.scala 41:38:@27849.4]
  assign _T_66692 = select_12 == 6'h1c; // @[Switch.scala 41:52:@27851.4]
  assign output_28_12 = io_outValid_12 & _T_66692; // @[Switch.scala 41:38:@27852.4]
  assign _T_66695 = select_13 == 6'h1c; // @[Switch.scala 41:52:@27854.4]
  assign output_28_13 = io_outValid_13 & _T_66695; // @[Switch.scala 41:38:@27855.4]
  assign _T_66698 = select_14 == 6'h1c; // @[Switch.scala 41:52:@27857.4]
  assign output_28_14 = io_outValid_14 & _T_66698; // @[Switch.scala 41:38:@27858.4]
  assign _T_66701 = select_15 == 6'h1c; // @[Switch.scala 41:52:@27860.4]
  assign output_28_15 = io_outValid_15 & _T_66701; // @[Switch.scala 41:38:@27861.4]
  assign _T_66704 = select_16 == 6'h1c; // @[Switch.scala 41:52:@27863.4]
  assign output_28_16 = io_outValid_16 & _T_66704; // @[Switch.scala 41:38:@27864.4]
  assign _T_66707 = select_17 == 6'h1c; // @[Switch.scala 41:52:@27866.4]
  assign output_28_17 = io_outValid_17 & _T_66707; // @[Switch.scala 41:38:@27867.4]
  assign _T_66710 = select_18 == 6'h1c; // @[Switch.scala 41:52:@27869.4]
  assign output_28_18 = io_outValid_18 & _T_66710; // @[Switch.scala 41:38:@27870.4]
  assign _T_66713 = select_19 == 6'h1c; // @[Switch.scala 41:52:@27872.4]
  assign output_28_19 = io_outValid_19 & _T_66713; // @[Switch.scala 41:38:@27873.4]
  assign _T_66716 = select_20 == 6'h1c; // @[Switch.scala 41:52:@27875.4]
  assign output_28_20 = io_outValid_20 & _T_66716; // @[Switch.scala 41:38:@27876.4]
  assign _T_66719 = select_21 == 6'h1c; // @[Switch.scala 41:52:@27878.4]
  assign output_28_21 = io_outValid_21 & _T_66719; // @[Switch.scala 41:38:@27879.4]
  assign _T_66722 = select_22 == 6'h1c; // @[Switch.scala 41:52:@27881.4]
  assign output_28_22 = io_outValid_22 & _T_66722; // @[Switch.scala 41:38:@27882.4]
  assign _T_66725 = select_23 == 6'h1c; // @[Switch.scala 41:52:@27884.4]
  assign output_28_23 = io_outValid_23 & _T_66725; // @[Switch.scala 41:38:@27885.4]
  assign _T_66728 = select_24 == 6'h1c; // @[Switch.scala 41:52:@27887.4]
  assign output_28_24 = io_outValid_24 & _T_66728; // @[Switch.scala 41:38:@27888.4]
  assign _T_66731 = select_25 == 6'h1c; // @[Switch.scala 41:52:@27890.4]
  assign output_28_25 = io_outValid_25 & _T_66731; // @[Switch.scala 41:38:@27891.4]
  assign _T_66734 = select_26 == 6'h1c; // @[Switch.scala 41:52:@27893.4]
  assign output_28_26 = io_outValid_26 & _T_66734; // @[Switch.scala 41:38:@27894.4]
  assign _T_66737 = select_27 == 6'h1c; // @[Switch.scala 41:52:@27896.4]
  assign output_28_27 = io_outValid_27 & _T_66737; // @[Switch.scala 41:38:@27897.4]
  assign _T_66740 = select_28 == 6'h1c; // @[Switch.scala 41:52:@27899.4]
  assign output_28_28 = io_outValid_28 & _T_66740; // @[Switch.scala 41:38:@27900.4]
  assign _T_66743 = select_29 == 6'h1c; // @[Switch.scala 41:52:@27902.4]
  assign output_28_29 = io_outValid_29 & _T_66743; // @[Switch.scala 41:38:@27903.4]
  assign _T_66746 = select_30 == 6'h1c; // @[Switch.scala 41:52:@27905.4]
  assign output_28_30 = io_outValid_30 & _T_66746; // @[Switch.scala 41:38:@27906.4]
  assign _T_66749 = select_31 == 6'h1c; // @[Switch.scala 41:52:@27908.4]
  assign output_28_31 = io_outValid_31 & _T_66749; // @[Switch.scala 41:38:@27909.4]
  assign _T_66752 = select_32 == 6'h1c; // @[Switch.scala 41:52:@27911.4]
  assign output_28_32 = io_outValid_32 & _T_66752; // @[Switch.scala 41:38:@27912.4]
  assign _T_66755 = select_33 == 6'h1c; // @[Switch.scala 41:52:@27914.4]
  assign output_28_33 = io_outValid_33 & _T_66755; // @[Switch.scala 41:38:@27915.4]
  assign _T_66758 = select_34 == 6'h1c; // @[Switch.scala 41:52:@27917.4]
  assign output_28_34 = io_outValid_34 & _T_66758; // @[Switch.scala 41:38:@27918.4]
  assign _T_66761 = select_35 == 6'h1c; // @[Switch.scala 41:52:@27920.4]
  assign output_28_35 = io_outValid_35 & _T_66761; // @[Switch.scala 41:38:@27921.4]
  assign _T_66764 = select_36 == 6'h1c; // @[Switch.scala 41:52:@27923.4]
  assign output_28_36 = io_outValid_36 & _T_66764; // @[Switch.scala 41:38:@27924.4]
  assign _T_66767 = select_37 == 6'h1c; // @[Switch.scala 41:52:@27926.4]
  assign output_28_37 = io_outValid_37 & _T_66767; // @[Switch.scala 41:38:@27927.4]
  assign _T_66770 = select_38 == 6'h1c; // @[Switch.scala 41:52:@27929.4]
  assign output_28_38 = io_outValid_38 & _T_66770; // @[Switch.scala 41:38:@27930.4]
  assign _T_66773 = select_39 == 6'h1c; // @[Switch.scala 41:52:@27932.4]
  assign output_28_39 = io_outValid_39 & _T_66773; // @[Switch.scala 41:38:@27933.4]
  assign _T_66776 = select_40 == 6'h1c; // @[Switch.scala 41:52:@27935.4]
  assign output_28_40 = io_outValid_40 & _T_66776; // @[Switch.scala 41:38:@27936.4]
  assign _T_66779 = select_41 == 6'h1c; // @[Switch.scala 41:52:@27938.4]
  assign output_28_41 = io_outValid_41 & _T_66779; // @[Switch.scala 41:38:@27939.4]
  assign _T_66782 = select_42 == 6'h1c; // @[Switch.scala 41:52:@27941.4]
  assign output_28_42 = io_outValid_42 & _T_66782; // @[Switch.scala 41:38:@27942.4]
  assign _T_66785 = select_43 == 6'h1c; // @[Switch.scala 41:52:@27944.4]
  assign output_28_43 = io_outValid_43 & _T_66785; // @[Switch.scala 41:38:@27945.4]
  assign _T_66788 = select_44 == 6'h1c; // @[Switch.scala 41:52:@27947.4]
  assign output_28_44 = io_outValid_44 & _T_66788; // @[Switch.scala 41:38:@27948.4]
  assign _T_66791 = select_45 == 6'h1c; // @[Switch.scala 41:52:@27950.4]
  assign output_28_45 = io_outValid_45 & _T_66791; // @[Switch.scala 41:38:@27951.4]
  assign _T_66794 = select_46 == 6'h1c; // @[Switch.scala 41:52:@27953.4]
  assign output_28_46 = io_outValid_46 & _T_66794; // @[Switch.scala 41:38:@27954.4]
  assign _T_66797 = select_47 == 6'h1c; // @[Switch.scala 41:52:@27956.4]
  assign output_28_47 = io_outValid_47 & _T_66797; // @[Switch.scala 41:38:@27957.4]
  assign _T_66800 = select_48 == 6'h1c; // @[Switch.scala 41:52:@27959.4]
  assign output_28_48 = io_outValid_48 & _T_66800; // @[Switch.scala 41:38:@27960.4]
  assign _T_66803 = select_49 == 6'h1c; // @[Switch.scala 41:52:@27962.4]
  assign output_28_49 = io_outValid_49 & _T_66803; // @[Switch.scala 41:38:@27963.4]
  assign _T_66806 = select_50 == 6'h1c; // @[Switch.scala 41:52:@27965.4]
  assign output_28_50 = io_outValid_50 & _T_66806; // @[Switch.scala 41:38:@27966.4]
  assign _T_66809 = select_51 == 6'h1c; // @[Switch.scala 41:52:@27968.4]
  assign output_28_51 = io_outValid_51 & _T_66809; // @[Switch.scala 41:38:@27969.4]
  assign _T_66812 = select_52 == 6'h1c; // @[Switch.scala 41:52:@27971.4]
  assign output_28_52 = io_outValid_52 & _T_66812; // @[Switch.scala 41:38:@27972.4]
  assign _T_66815 = select_53 == 6'h1c; // @[Switch.scala 41:52:@27974.4]
  assign output_28_53 = io_outValid_53 & _T_66815; // @[Switch.scala 41:38:@27975.4]
  assign _T_66818 = select_54 == 6'h1c; // @[Switch.scala 41:52:@27977.4]
  assign output_28_54 = io_outValid_54 & _T_66818; // @[Switch.scala 41:38:@27978.4]
  assign _T_66821 = select_55 == 6'h1c; // @[Switch.scala 41:52:@27980.4]
  assign output_28_55 = io_outValid_55 & _T_66821; // @[Switch.scala 41:38:@27981.4]
  assign _T_66824 = select_56 == 6'h1c; // @[Switch.scala 41:52:@27983.4]
  assign output_28_56 = io_outValid_56 & _T_66824; // @[Switch.scala 41:38:@27984.4]
  assign _T_66827 = select_57 == 6'h1c; // @[Switch.scala 41:52:@27986.4]
  assign output_28_57 = io_outValid_57 & _T_66827; // @[Switch.scala 41:38:@27987.4]
  assign _T_66830 = select_58 == 6'h1c; // @[Switch.scala 41:52:@27989.4]
  assign output_28_58 = io_outValid_58 & _T_66830; // @[Switch.scala 41:38:@27990.4]
  assign _T_66833 = select_59 == 6'h1c; // @[Switch.scala 41:52:@27992.4]
  assign output_28_59 = io_outValid_59 & _T_66833; // @[Switch.scala 41:38:@27993.4]
  assign _T_66836 = select_60 == 6'h1c; // @[Switch.scala 41:52:@27995.4]
  assign output_28_60 = io_outValid_60 & _T_66836; // @[Switch.scala 41:38:@27996.4]
  assign _T_66839 = select_61 == 6'h1c; // @[Switch.scala 41:52:@27998.4]
  assign output_28_61 = io_outValid_61 & _T_66839; // @[Switch.scala 41:38:@27999.4]
  assign _T_66842 = select_62 == 6'h1c; // @[Switch.scala 41:52:@28001.4]
  assign output_28_62 = io_outValid_62 & _T_66842; // @[Switch.scala 41:38:@28002.4]
  assign _T_66845 = select_63 == 6'h1c; // @[Switch.scala 41:52:@28004.4]
  assign output_28_63 = io_outValid_63 & _T_66845; // @[Switch.scala 41:38:@28005.4]
  assign _T_66853 = {output_28_7,output_28_6,output_28_5,output_28_4,output_28_3,output_28_2,output_28_1,output_28_0}; // @[Switch.scala 43:31:@28013.4]
  assign _T_66861 = {output_28_15,output_28_14,output_28_13,output_28_12,output_28_11,output_28_10,output_28_9,output_28_8,_T_66853}; // @[Switch.scala 43:31:@28021.4]
  assign _T_66868 = {output_28_23,output_28_22,output_28_21,output_28_20,output_28_19,output_28_18,output_28_17,output_28_16}; // @[Switch.scala 43:31:@28028.4]
  assign _T_66877 = {output_28_31,output_28_30,output_28_29,output_28_28,output_28_27,output_28_26,output_28_25,output_28_24,_T_66868,_T_66861}; // @[Switch.scala 43:31:@28037.4]
  assign _T_66884 = {output_28_39,output_28_38,output_28_37,output_28_36,output_28_35,output_28_34,output_28_33,output_28_32}; // @[Switch.scala 43:31:@28044.4]
  assign _T_66892 = {output_28_47,output_28_46,output_28_45,output_28_44,output_28_43,output_28_42,output_28_41,output_28_40,_T_66884}; // @[Switch.scala 43:31:@28052.4]
  assign _T_66899 = {output_28_55,output_28_54,output_28_53,output_28_52,output_28_51,output_28_50,output_28_49,output_28_48}; // @[Switch.scala 43:31:@28059.4]
  assign _T_66908 = {output_28_63,output_28_62,output_28_61,output_28_60,output_28_59,output_28_58,output_28_57,output_28_56,_T_66899,_T_66892}; // @[Switch.scala 43:31:@28068.4]
  assign _T_66909 = {_T_66908,_T_66877}; // @[Switch.scala 43:31:@28069.4]
  assign _T_66913 = select_0 == 6'h1d; // @[Switch.scala 41:52:@28072.4]
  assign output_29_0 = io_outValid_0 & _T_66913; // @[Switch.scala 41:38:@28073.4]
  assign _T_66916 = select_1 == 6'h1d; // @[Switch.scala 41:52:@28075.4]
  assign output_29_1 = io_outValid_1 & _T_66916; // @[Switch.scala 41:38:@28076.4]
  assign _T_66919 = select_2 == 6'h1d; // @[Switch.scala 41:52:@28078.4]
  assign output_29_2 = io_outValid_2 & _T_66919; // @[Switch.scala 41:38:@28079.4]
  assign _T_66922 = select_3 == 6'h1d; // @[Switch.scala 41:52:@28081.4]
  assign output_29_3 = io_outValid_3 & _T_66922; // @[Switch.scala 41:38:@28082.4]
  assign _T_66925 = select_4 == 6'h1d; // @[Switch.scala 41:52:@28084.4]
  assign output_29_4 = io_outValid_4 & _T_66925; // @[Switch.scala 41:38:@28085.4]
  assign _T_66928 = select_5 == 6'h1d; // @[Switch.scala 41:52:@28087.4]
  assign output_29_5 = io_outValid_5 & _T_66928; // @[Switch.scala 41:38:@28088.4]
  assign _T_66931 = select_6 == 6'h1d; // @[Switch.scala 41:52:@28090.4]
  assign output_29_6 = io_outValid_6 & _T_66931; // @[Switch.scala 41:38:@28091.4]
  assign _T_66934 = select_7 == 6'h1d; // @[Switch.scala 41:52:@28093.4]
  assign output_29_7 = io_outValid_7 & _T_66934; // @[Switch.scala 41:38:@28094.4]
  assign _T_66937 = select_8 == 6'h1d; // @[Switch.scala 41:52:@28096.4]
  assign output_29_8 = io_outValid_8 & _T_66937; // @[Switch.scala 41:38:@28097.4]
  assign _T_66940 = select_9 == 6'h1d; // @[Switch.scala 41:52:@28099.4]
  assign output_29_9 = io_outValid_9 & _T_66940; // @[Switch.scala 41:38:@28100.4]
  assign _T_66943 = select_10 == 6'h1d; // @[Switch.scala 41:52:@28102.4]
  assign output_29_10 = io_outValid_10 & _T_66943; // @[Switch.scala 41:38:@28103.4]
  assign _T_66946 = select_11 == 6'h1d; // @[Switch.scala 41:52:@28105.4]
  assign output_29_11 = io_outValid_11 & _T_66946; // @[Switch.scala 41:38:@28106.4]
  assign _T_66949 = select_12 == 6'h1d; // @[Switch.scala 41:52:@28108.4]
  assign output_29_12 = io_outValid_12 & _T_66949; // @[Switch.scala 41:38:@28109.4]
  assign _T_66952 = select_13 == 6'h1d; // @[Switch.scala 41:52:@28111.4]
  assign output_29_13 = io_outValid_13 & _T_66952; // @[Switch.scala 41:38:@28112.4]
  assign _T_66955 = select_14 == 6'h1d; // @[Switch.scala 41:52:@28114.4]
  assign output_29_14 = io_outValid_14 & _T_66955; // @[Switch.scala 41:38:@28115.4]
  assign _T_66958 = select_15 == 6'h1d; // @[Switch.scala 41:52:@28117.4]
  assign output_29_15 = io_outValid_15 & _T_66958; // @[Switch.scala 41:38:@28118.4]
  assign _T_66961 = select_16 == 6'h1d; // @[Switch.scala 41:52:@28120.4]
  assign output_29_16 = io_outValid_16 & _T_66961; // @[Switch.scala 41:38:@28121.4]
  assign _T_66964 = select_17 == 6'h1d; // @[Switch.scala 41:52:@28123.4]
  assign output_29_17 = io_outValid_17 & _T_66964; // @[Switch.scala 41:38:@28124.4]
  assign _T_66967 = select_18 == 6'h1d; // @[Switch.scala 41:52:@28126.4]
  assign output_29_18 = io_outValid_18 & _T_66967; // @[Switch.scala 41:38:@28127.4]
  assign _T_66970 = select_19 == 6'h1d; // @[Switch.scala 41:52:@28129.4]
  assign output_29_19 = io_outValid_19 & _T_66970; // @[Switch.scala 41:38:@28130.4]
  assign _T_66973 = select_20 == 6'h1d; // @[Switch.scala 41:52:@28132.4]
  assign output_29_20 = io_outValid_20 & _T_66973; // @[Switch.scala 41:38:@28133.4]
  assign _T_66976 = select_21 == 6'h1d; // @[Switch.scala 41:52:@28135.4]
  assign output_29_21 = io_outValid_21 & _T_66976; // @[Switch.scala 41:38:@28136.4]
  assign _T_66979 = select_22 == 6'h1d; // @[Switch.scala 41:52:@28138.4]
  assign output_29_22 = io_outValid_22 & _T_66979; // @[Switch.scala 41:38:@28139.4]
  assign _T_66982 = select_23 == 6'h1d; // @[Switch.scala 41:52:@28141.4]
  assign output_29_23 = io_outValid_23 & _T_66982; // @[Switch.scala 41:38:@28142.4]
  assign _T_66985 = select_24 == 6'h1d; // @[Switch.scala 41:52:@28144.4]
  assign output_29_24 = io_outValid_24 & _T_66985; // @[Switch.scala 41:38:@28145.4]
  assign _T_66988 = select_25 == 6'h1d; // @[Switch.scala 41:52:@28147.4]
  assign output_29_25 = io_outValid_25 & _T_66988; // @[Switch.scala 41:38:@28148.4]
  assign _T_66991 = select_26 == 6'h1d; // @[Switch.scala 41:52:@28150.4]
  assign output_29_26 = io_outValid_26 & _T_66991; // @[Switch.scala 41:38:@28151.4]
  assign _T_66994 = select_27 == 6'h1d; // @[Switch.scala 41:52:@28153.4]
  assign output_29_27 = io_outValid_27 & _T_66994; // @[Switch.scala 41:38:@28154.4]
  assign _T_66997 = select_28 == 6'h1d; // @[Switch.scala 41:52:@28156.4]
  assign output_29_28 = io_outValid_28 & _T_66997; // @[Switch.scala 41:38:@28157.4]
  assign _T_67000 = select_29 == 6'h1d; // @[Switch.scala 41:52:@28159.4]
  assign output_29_29 = io_outValid_29 & _T_67000; // @[Switch.scala 41:38:@28160.4]
  assign _T_67003 = select_30 == 6'h1d; // @[Switch.scala 41:52:@28162.4]
  assign output_29_30 = io_outValid_30 & _T_67003; // @[Switch.scala 41:38:@28163.4]
  assign _T_67006 = select_31 == 6'h1d; // @[Switch.scala 41:52:@28165.4]
  assign output_29_31 = io_outValid_31 & _T_67006; // @[Switch.scala 41:38:@28166.4]
  assign _T_67009 = select_32 == 6'h1d; // @[Switch.scala 41:52:@28168.4]
  assign output_29_32 = io_outValid_32 & _T_67009; // @[Switch.scala 41:38:@28169.4]
  assign _T_67012 = select_33 == 6'h1d; // @[Switch.scala 41:52:@28171.4]
  assign output_29_33 = io_outValid_33 & _T_67012; // @[Switch.scala 41:38:@28172.4]
  assign _T_67015 = select_34 == 6'h1d; // @[Switch.scala 41:52:@28174.4]
  assign output_29_34 = io_outValid_34 & _T_67015; // @[Switch.scala 41:38:@28175.4]
  assign _T_67018 = select_35 == 6'h1d; // @[Switch.scala 41:52:@28177.4]
  assign output_29_35 = io_outValid_35 & _T_67018; // @[Switch.scala 41:38:@28178.4]
  assign _T_67021 = select_36 == 6'h1d; // @[Switch.scala 41:52:@28180.4]
  assign output_29_36 = io_outValid_36 & _T_67021; // @[Switch.scala 41:38:@28181.4]
  assign _T_67024 = select_37 == 6'h1d; // @[Switch.scala 41:52:@28183.4]
  assign output_29_37 = io_outValid_37 & _T_67024; // @[Switch.scala 41:38:@28184.4]
  assign _T_67027 = select_38 == 6'h1d; // @[Switch.scala 41:52:@28186.4]
  assign output_29_38 = io_outValid_38 & _T_67027; // @[Switch.scala 41:38:@28187.4]
  assign _T_67030 = select_39 == 6'h1d; // @[Switch.scala 41:52:@28189.4]
  assign output_29_39 = io_outValid_39 & _T_67030; // @[Switch.scala 41:38:@28190.4]
  assign _T_67033 = select_40 == 6'h1d; // @[Switch.scala 41:52:@28192.4]
  assign output_29_40 = io_outValid_40 & _T_67033; // @[Switch.scala 41:38:@28193.4]
  assign _T_67036 = select_41 == 6'h1d; // @[Switch.scala 41:52:@28195.4]
  assign output_29_41 = io_outValid_41 & _T_67036; // @[Switch.scala 41:38:@28196.4]
  assign _T_67039 = select_42 == 6'h1d; // @[Switch.scala 41:52:@28198.4]
  assign output_29_42 = io_outValid_42 & _T_67039; // @[Switch.scala 41:38:@28199.4]
  assign _T_67042 = select_43 == 6'h1d; // @[Switch.scala 41:52:@28201.4]
  assign output_29_43 = io_outValid_43 & _T_67042; // @[Switch.scala 41:38:@28202.4]
  assign _T_67045 = select_44 == 6'h1d; // @[Switch.scala 41:52:@28204.4]
  assign output_29_44 = io_outValid_44 & _T_67045; // @[Switch.scala 41:38:@28205.4]
  assign _T_67048 = select_45 == 6'h1d; // @[Switch.scala 41:52:@28207.4]
  assign output_29_45 = io_outValid_45 & _T_67048; // @[Switch.scala 41:38:@28208.4]
  assign _T_67051 = select_46 == 6'h1d; // @[Switch.scala 41:52:@28210.4]
  assign output_29_46 = io_outValid_46 & _T_67051; // @[Switch.scala 41:38:@28211.4]
  assign _T_67054 = select_47 == 6'h1d; // @[Switch.scala 41:52:@28213.4]
  assign output_29_47 = io_outValid_47 & _T_67054; // @[Switch.scala 41:38:@28214.4]
  assign _T_67057 = select_48 == 6'h1d; // @[Switch.scala 41:52:@28216.4]
  assign output_29_48 = io_outValid_48 & _T_67057; // @[Switch.scala 41:38:@28217.4]
  assign _T_67060 = select_49 == 6'h1d; // @[Switch.scala 41:52:@28219.4]
  assign output_29_49 = io_outValid_49 & _T_67060; // @[Switch.scala 41:38:@28220.4]
  assign _T_67063 = select_50 == 6'h1d; // @[Switch.scala 41:52:@28222.4]
  assign output_29_50 = io_outValid_50 & _T_67063; // @[Switch.scala 41:38:@28223.4]
  assign _T_67066 = select_51 == 6'h1d; // @[Switch.scala 41:52:@28225.4]
  assign output_29_51 = io_outValid_51 & _T_67066; // @[Switch.scala 41:38:@28226.4]
  assign _T_67069 = select_52 == 6'h1d; // @[Switch.scala 41:52:@28228.4]
  assign output_29_52 = io_outValid_52 & _T_67069; // @[Switch.scala 41:38:@28229.4]
  assign _T_67072 = select_53 == 6'h1d; // @[Switch.scala 41:52:@28231.4]
  assign output_29_53 = io_outValid_53 & _T_67072; // @[Switch.scala 41:38:@28232.4]
  assign _T_67075 = select_54 == 6'h1d; // @[Switch.scala 41:52:@28234.4]
  assign output_29_54 = io_outValid_54 & _T_67075; // @[Switch.scala 41:38:@28235.4]
  assign _T_67078 = select_55 == 6'h1d; // @[Switch.scala 41:52:@28237.4]
  assign output_29_55 = io_outValid_55 & _T_67078; // @[Switch.scala 41:38:@28238.4]
  assign _T_67081 = select_56 == 6'h1d; // @[Switch.scala 41:52:@28240.4]
  assign output_29_56 = io_outValid_56 & _T_67081; // @[Switch.scala 41:38:@28241.4]
  assign _T_67084 = select_57 == 6'h1d; // @[Switch.scala 41:52:@28243.4]
  assign output_29_57 = io_outValid_57 & _T_67084; // @[Switch.scala 41:38:@28244.4]
  assign _T_67087 = select_58 == 6'h1d; // @[Switch.scala 41:52:@28246.4]
  assign output_29_58 = io_outValid_58 & _T_67087; // @[Switch.scala 41:38:@28247.4]
  assign _T_67090 = select_59 == 6'h1d; // @[Switch.scala 41:52:@28249.4]
  assign output_29_59 = io_outValid_59 & _T_67090; // @[Switch.scala 41:38:@28250.4]
  assign _T_67093 = select_60 == 6'h1d; // @[Switch.scala 41:52:@28252.4]
  assign output_29_60 = io_outValid_60 & _T_67093; // @[Switch.scala 41:38:@28253.4]
  assign _T_67096 = select_61 == 6'h1d; // @[Switch.scala 41:52:@28255.4]
  assign output_29_61 = io_outValid_61 & _T_67096; // @[Switch.scala 41:38:@28256.4]
  assign _T_67099 = select_62 == 6'h1d; // @[Switch.scala 41:52:@28258.4]
  assign output_29_62 = io_outValid_62 & _T_67099; // @[Switch.scala 41:38:@28259.4]
  assign _T_67102 = select_63 == 6'h1d; // @[Switch.scala 41:52:@28261.4]
  assign output_29_63 = io_outValid_63 & _T_67102; // @[Switch.scala 41:38:@28262.4]
  assign _T_67110 = {output_29_7,output_29_6,output_29_5,output_29_4,output_29_3,output_29_2,output_29_1,output_29_0}; // @[Switch.scala 43:31:@28270.4]
  assign _T_67118 = {output_29_15,output_29_14,output_29_13,output_29_12,output_29_11,output_29_10,output_29_9,output_29_8,_T_67110}; // @[Switch.scala 43:31:@28278.4]
  assign _T_67125 = {output_29_23,output_29_22,output_29_21,output_29_20,output_29_19,output_29_18,output_29_17,output_29_16}; // @[Switch.scala 43:31:@28285.4]
  assign _T_67134 = {output_29_31,output_29_30,output_29_29,output_29_28,output_29_27,output_29_26,output_29_25,output_29_24,_T_67125,_T_67118}; // @[Switch.scala 43:31:@28294.4]
  assign _T_67141 = {output_29_39,output_29_38,output_29_37,output_29_36,output_29_35,output_29_34,output_29_33,output_29_32}; // @[Switch.scala 43:31:@28301.4]
  assign _T_67149 = {output_29_47,output_29_46,output_29_45,output_29_44,output_29_43,output_29_42,output_29_41,output_29_40,_T_67141}; // @[Switch.scala 43:31:@28309.4]
  assign _T_67156 = {output_29_55,output_29_54,output_29_53,output_29_52,output_29_51,output_29_50,output_29_49,output_29_48}; // @[Switch.scala 43:31:@28316.4]
  assign _T_67165 = {output_29_63,output_29_62,output_29_61,output_29_60,output_29_59,output_29_58,output_29_57,output_29_56,_T_67156,_T_67149}; // @[Switch.scala 43:31:@28325.4]
  assign _T_67166 = {_T_67165,_T_67134}; // @[Switch.scala 43:31:@28326.4]
  assign _T_67170 = select_0 == 6'h1e; // @[Switch.scala 41:52:@28329.4]
  assign output_30_0 = io_outValid_0 & _T_67170; // @[Switch.scala 41:38:@28330.4]
  assign _T_67173 = select_1 == 6'h1e; // @[Switch.scala 41:52:@28332.4]
  assign output_30_1 = io_outValid_1 & _T_67173; // @[Switch.scala 41:38:@28333.4]
  assign _T_67176 = select_2 == 6'h1e; // @[Switch.scala 41:52:@28335.4]
  assign output_30_2 = io_outValid_2 & _T_67176; // @[Switch.scala 41:38:@28336.4]
  assign _T_67179 = select_3 == 6'h1e; // @[Switch.scala 41:52:@28338.4]
  assign output_30_3 = io_outValid_3 & _T_67179; // @[Switch.scala 41:38:@28339.4]
  assign _T_67182 = select_4 == 6'h1e; // @[Switch.scala 41:52:@28341.4]
  assign output_30_4 = io_outValid_4 & _T_67182; // @[Switch.scala 41:38:@28342.4]
  assign _T_67185 = select_5 == 6'h1e; // @[Switch.scala 41:52:@28344.4]
  assign output_30_5 = io_outValid_5 & _T_67185; // @[Switch.scala 41:38:@28345.4]
  assign _T_67188 = select_6 == 6'h1e; // @[Switch.scala 41:52:@28347.4]
  assign output_30_6 = io_outValid_6 & _T_67188; // @[Switch.scala 41:38:@28348.4]
  assign _T_67191 = select_7 == 6'h1e; // @[Switch.scala 41:52:@28350.4]
  assign output_30_7 = io_outValid_7 & _T_67191; // @[Switch.scala 41:38:@28351.4]
  assign _T_67194 = select_8 == 6'h1e; // @[Switch.scala 41:52:@28353.4]
  assign output_30_8 = io_outValid_8 & _T_67194; // @[Switch.scala 41:38:@28354.4]
  assign _T_67197 = select_9 == 6'h1e; // @[Switch.scala 41:52:@28356.4]
  assign output_30_9 = io_outValid_9 & _T_67197; // @[Switch.scala 41:38:@28357.4]
  assign _T_67200 = select_10 == 6'h1e; // @[Switch.scala 41:52:@28359.4]
  assign output_30_10 = io_outValid_10 & _T_67200; // @[Switch.scala 41:38:@28360.4]
  assign _T_67203 = select_11 == 6'h1e; // @[Switch.scala 41:52:@28362.4]
  assign output_30_11 = io_outValid_11 & _T_67203; // @[Switch.scala 41:38:@28363.4]
  assign _T_67206 = select_12 == 6'h1e; // @[Switch.scala 41:52:@28365.4]
  assign output_30_12 = io_outValid_12 & _T_67206; // @[Switch.scala 41:38:@28366.4]
  assign _T_67209 = select_13 == 6'h1e; // @[Switch.scala 41:52:@28368.4]
  assign output_30_13 = io_outValid_13 & _T_67209; // @[Switch.scala 41:38:@28369.4]
  assign _T_67212 = select_14 == 6'h1e; // @[Switch.scala 41:52:@28371.4]
  assign output_30_14 = io_outValid_14 & _T_67212; // @[Switch.scala 41:38:@28372.4]
  assign _T_67215 = select_15 == 6'h1e; // @[Switch.scala 41:52:@28374.4]
  assign output_30_15 = io_outValid_15 & _T_67215; // @[Switch.scala 41:38:@28375.4]
  assign _T_67218 = select_16 == 6'h1e; // @[Switch.scala 41:52:@28377.4]
  assign output_30_16 = io_outValid_16 & _T_67218; // @[Switch.scala 41:38:@28378.4]
  assign _T_67221 = select_17 == 6'h1e; // @[Switch.scala 41:52:@28380.4]
  assign output_30_17 = io_outValid_17 & _T_67221; // @[Switch.scala 41:38:@28381.4]
  assign _T_67224 = select_18 == 6'h1e; // @[Switch.scala 41:52:@28383.4]
  assign output_30_18 = io_outValid_18 & _T_67224; // @[Switch.scala 41:38:@28384.4]
  assign _T_67227 = select_19 == 6'h1e; // @[Switch.scala 41:52:@28386.4]
  assign output_30_19 = io_outValid_19 & _T_67227; // @[Switch.scala 41:38:@28387.4]
  assign _T_67230 = select_20 == 6'h1e; // @[Switch.scala 41:52:@28389.4]
  assign output_30_20 = io_outValid_20 & _T_67230; // @[Switch.scala 41:38:@28390.4]
  assign _T_67233 = select_21 == 6'h1e; // @[Switch.scala 41:52:@28392.4]
  assign output_30_21 = io_outValid_21 & _T_67233; // @[Switch.scala 41:38:@28393.4]
  assign _T_67236 = select_22 == 6'h1e; // @[Switch.scala 41:52:@28395.4]
  assign output_30_22 = io_outValid_22 & _T_67236; // @[Switch.scala 41:38:@28396.4]
  assign _T_67239 = select_23 == 6'h1e; // @[Switch.scala 41:52:@28398.4]
  assign output_30_23 = io_outValid_23 & _T_67239; // @[Switch.scala 41:38:@28399.4]
  assign _T_67242 = select_24 == 6'h1e; // @[Switch.scala 41:52:@28401.4]
  assign output_30_24 = io_outValid_24 & _T_67242; // @[Switch.scala 41:38:@28402.4]
  assign _T_67245 = select_25 == 6'h1e; // @[Switch.scala 41:52:@28404.4]
  assign output_30_25 = io_outValid_25 & _T_67245; // @[Switch.scala 41:38:@28405.4]
  assign _T_67248 = select_26 == 6'h1e; // @[Switch.scala 41:52:@28407.4]
  assign output_30_26 = io_outValid_26 & _T_67248; // @[Switch.scala 41:38:@28408.4]
  assign _T_67251 = select_27 == 6'h1e; // @[Switch.scala 41:52:@28410.4]
  assign output_30_27 = io_outValid_27 & _T_67251; // @[Switch.scala 41:38:@28411.4]
  assign _T_67254 = select_28 == 6'h1e; // @[Switch.scala 41:52:@28413.4]
  assign output_30_28 = io_outValid_28 & _T_67254; // @[Switch.scala 41:38:@28414.4]
  assign _T_67257 = select_29 == 6'h1e; // @[Switch.scala 41:52:@28416.4]
  assign output_30_29 = io_outValid_29 & _T_67257; // @[Switch.scala 41:38:@28417.4]
  assign _T_67260 = select_30 == 6'h1e; // @[Switch.scala 41:52:@28419.4]
  assign output_30_30 = io_outValid_30 & _T_67260; // @[Switch.scala 41:38:@28420.4]
  assign _T_67263 = select_31 == 6'h1e; // @[Switch.scala 41:52:@28422.4]
  assign output_30_31 = io_outValid_31 & _T_67263; // @[Switch.scala 41:38:@28423.4]
  assign _T_67266 = select_32 == 6'h1e; // @[Switch.scala 41:52:@28425.4]
  assign output_30_32 = io_outValid_32 & _T_67266; // @[Switch.scala 41:38:@28426.4]
  assign _T_67269 = select_33 == 6'h1e; // @[Switch.scala 41:52:@28428.4]
  assign output_30_33 = io_outValid_33 & _T_67269; // @[Switch.scala 41:38:@28429.4]
  assign _T_67272 = select_34 == 6'h1e; // @[Switch.scala 41:52:@28431.4]
  assign output_30_34 = io_outValid_34 & _T_67272; // @[Switch.scala 41:38:@28432.4]
  assign _T_67275 = select_35 == 6'h1e; // @[Switch.scala 41:52:@28434.4]
  assign output_30_35 = io_outValid_35 & _T_67275; // @[Switch.scala 41:38:@28435.4]
  assign _T_67278 = select_36 == 6'h1e; // @[Switch.scala 41:52:@28437.4]
  assign output_30_36 = io_outValid_36 & _T_67278; // @[Switch.scala 41:38:@28438.4]
  assign _T_67281 = select_37 == 6'h1e; // @[Switch.scala 41:52:@28440.4]
  assign output_30_37 = io_outValid_37 & _T_67281; // @[Switch.scala 41:38:@28441.4]
  assign _T_67284 = select_38 == 6'h1e; // @[Switch.scala 41:52:@28443.4]
  assign output_30_38 = io_outValid_38 & _T_67284; // @[Switch.scala 41:38:@28444.4]
  assign _T_67287 = select_39 == 6'h1e; // @[Switch.scala 41:52:@28446.4]
  assign output_30_39 = io_outValid_39 & _T_67287; // @[Switch.scala 41:38:@28447.4]
  assign _T_67290 = select_40 == 6'h1e; // @[Switch.scala 41:52:@28449.4]
  assign output_30_40 = io_outValid_40 & _T_67290; // @[Switch.scala 41:38:@28450.4]
  assign _T_67293 = select_41 == 6'h1e; // @[Switch.scala 41:52:@28452.4]
  assign output_30_41 = io_outValid_41 & _T_67293; // @[Switch.scala 41:38:@28453.4]
  assign _T_67296 = select_42 == 6'h1e; // @[Switch.scala 41:52:@28455.4]
  assign output_30_42 = io_outValid_42 & _T_67296; // @[Switch.scala 41:38:@28456.4]
  assign _T_67299 = select_43 == 6'h1e; // @[Switch.scala 41:52:@28458.4]
  assign output_30_43 = io_outValid_43 & _T_67299; // @[Switch.scala 41:38:@28459.4]
  assign _T_67302 = select_44 == 6'h1e; // @[Switch.scala 41:52:@28461.4]
  assign output_30_44 = io_outValid_44 & _T_67302; // @[Switch.scala 41:38:@28462.4]
  assign _T_67305 = select_45 == 6'h1e; // @[Switch.scala 41:52:@28464.4]
  assign output_30_45 = io_outValid_45 & _T_67305; // @[Switch.scala 41:38:@28465.4]
  assign _T_67308 = select_46 == 6'h1e; // @[Switch.scala 41:52:@28467.4]
  assign output_30_46 = io_outValid_46 & _T_67308; // @[Switch.scala 41:38:@28468.4]
  assign _T_67311 = select_47 == 6'h1e; // @[Switch.scala 41:52:@28470.4]
  assign output_30_47 = io_outValid_47 & _T_67311; // @[Switch.scala 41:38:@28471.4]
  assign _T_67314 = select_48 == 6'h1e; // @[Switch.scala 41:52:@28473.4]
  assign output_30_48 = io_outValid_48 & _T_67314; // @[Switch.scala 41:38:@28474.4]
  assign _T_67317 = select_49 == 6'h1e; // @[Switch.scala 41:52:@28476.4]
  assign output_30_49 = io_outValid_49 & _T_67317; // @[Switch.scala 41:38:@28477.4]
  assign _T_67320 = select_50 == 6'h1e; // @[Switch.scala 41:52:@28479.4]
  assign output_30_50 = io_outValid_50 & _T_67320; // @[Switch.scala 41:38:@28480.4]
  assign _T_67323 = select_51 == 6'h1e; // @[Switch.scala 41:52:@28482.4]
  assign output_30_51 = io_outValid_51 & _T_67323; // @[Switch.scala 41:38:@28483.4]
  assign _T_67326 = select_52 == 6'h1e; // @[Switch.scala 41:52:@28485.4]
  assign output_30_52 = io_outValid_52 & _T_67326; // @[Switch.scala 41:38:@28486.4]
  assign _T_67329 = select_53 == 6'h1e; // @[Switch.scala 41:52:@28488.4]
  assign output_30_53 = io_outValid_53 & _T_67329; // @[Switch.scala 41:38:@28489.4]
  assign _T_67332 = select_54 == 6'h1e; // @[Switch.scala 41:52:@28491.4]
  assign output_30_54 = io_outValid_54 & _T_67332; // @[Switch.scala 41:38:@28492.4]
  assign _T_67335 = select_55 == 6'h1e; // @[Switch.scala 41:52:@28494.4]
  assign output_30_55 = io_outValid_55 & _T_67335; // @[Switch.scala 41:38:@28495.4]
  assign _T_67338 = select_56 == 6'h1e; // @[Switch.scala 41:52:@28497.4]
  assign output_30_56 = io_outValid_56 & _T_67338; // @[Switch.scala 41:38:@28498.4]
  assign _T_67341 = select_57 == 6'h1e; // @[Switch.scala 41:52:@28500.4]
  assign output_30_57 = io_outValid_57 & _T_67341; // @[Switch.scala 41:38:@28501.4]
  assign _T_67344 = select_58 == 6'h1e; // @[Switch.scala 41:52:@28503.4]
  assign output_30_58 = io_outValid_58 & _T_67344; // @[Switch.scala 41:38:@28504.4]
  assign _T_67347 = select_59 == 6'h1e; // @[Switch.scala 41:52:@28506.4]
  assign output_30_59 = io_outValid_59 & _T_67347; // @[Switch.scala 41:38:@28507.4]
  assign _T_67350 = select_60 == 6'h1e; // @[Switch.scala 41:52:@28509.4]
  assign output_30_60 = io_outValid_60 & _T_67350; // @[Switch.scala 41:38:@28510.4]
  assign _T_67353 = select_61 == 6'h1e; // @[Switch.scala 41:52:@28512.4]
  assign output_30_61 = io_outValid_61 & _T_67353; // @[Switch.scala 41:38:@28513.4]
  assign _T_67356 = select_62 == 6'h1e; // @[Switch.scala 41:52:@28515.4]
  assign output_30_62 = io_outValid_62 & _T_67356; // @[Switch.scala 41:38:@28516.4]
  assign _T_67359 = select_63 == 6'h1e; // @[Switch.scala 41:52:@28518.4]
  assign output_30_63 = io_outValid_63 & _T_67359; // @[Switch.scala 41:38:@28519.4]
  assign _T_67367 = {output_30_7,output_30_6,output_30_5,output_30_4,output_30_3,output_30_2,output_30_1,output_30_0}; // @[Switch.scala 43:31:@28527.4]
  assign _T_67375 = {output_30_15,output_30_14,output_30_13,output_30_12,output_30_11,output_30_10,output_30_9,output_30_8,_T_67367}; // @[Switch.scala 43:31:@28535.4]
  assign _T_67382 = {output_30_23,output_30_22,output_30_21,output_30_20,output_30_19,output_30_18,output_30_17,output_30_16}; // @[Switch.scala 43:31:@28542.4]
  assign _T_67391 = {output_30_31,output_30_30,output_30_29,output_30_28,output_30_27,output_30_26,output_30_25,output_30_24,_T_67382,_T_67375}; // @[Switch.scala 43:31:@28551.4]
  assign _T_67398 = {output_30_39,output_30_38,output_30_37,output_30_36,output_30_35,output_30_34,output_30_33,output_30_32}; // @[Switch.scala 43:31:@28558.4]
  assign _T_67406 = {output_30_47,output_30_46,output_30_45,output_30_44,output_30_43,output_30_42,output_30_41,output_30_40,_T_67398}; // @[Switch.scala 43:31:@28566.4]
  assign _T_67413 = {output_30_55,output_30_54,output_30_53,output_30_52,output_30_51,output_30_50,output_30_49,output_30_48}; // @[Switch.scala 43:31:@28573.4]
  assign _T_67422 = {output_30_63,output_30_62,output_30_61,output_30_60,output_30_59,output_30_58,output_30_57,output_30_56,_T_67413,_T_67406}; // @[Switch.scala 43:31:@28582.4]
  assign _T_67423 = {_T_67422,_T_67391}; // @[Switch.scala 43:31:@28583.4]
  assign _T_67427 = select_0 == 6'h1f; // @[Switch.scala 41:52:@28586.4]
  assign output_31_0 = io_outValid_0 & _T_67427; // @[Switch.scala 41:38:@28587.4]
  assign _T_67430 = select_1 == 6'h1f; // @[Switch.scala 41:52:@28589.4]
  assign output_31_1 = io_outValid_1 & _T_67430; // @[Switch.scala 41:38:@28590.4]
  assign _T_67433 = select_2 == 6'h1f; // @[Switch.scala 41:52:@28592.4]
  assign output_31_2 = io_outValid_2 & _T_67433; // @[Switch.scala 41:38:@28593.4]
  assign _T_67436 = select_3 == 6'h1f; // @[Switch.scala 41:52:@28595.4]
  assign output_31_3 = io_outValid_3 & _T_67436; // @[Switch.scala 41:38:@28596.4]
  assign _T_67439 = select_4 == 6'h1f; // @[Switch.scala 41:52:@28598.4]
  assign output_31_4 = io_outValid_4 & _T_67439; // @[Switch.scala 41:38:@28599.4]
  assign _T_67442 = select_5 == 6'h1f; // @[Switch.scala 41:52:@28601.4]
  assign output_31_5 = io_outValid_5 & _T_67442; // @[Switch.scala 41:38:@28602.4]
  assign _T_67445 = select_6 == 6'h1f; // @[Switch.scala 41:52:@28604.4]
  assign output_31_6 = io_outValid_6 & _T_67445; // @[Switch.scala 41:38:@28605.4]
  assign _T_67448 = select_7 == 6'h1f; // @[Switch.scala 41:52:@28607.4]
  assign output_31_7 = io_outValid_7 & _T_67448; // @[Switch.scala 41:38:@28608.4]
  assign _T_67451 = select_8 == 6'h1f; // @[Switch.scala 41:52:@28610.4]
  assign output_31_8 = io_outValid_8 & _T_67451; // @[Switch.scala 41:38:@28611.4]
  assign _T_67454 = select_9 == 6'h1f; // @[Switch.scala 41:52:@28613.4]
  assign output_31_9 = io_outValid_9 & _T_67454; // @[Switch.scala 41:38:@28614.4]
  assign _T_67457 = select_10 == 6'h1f; // @[Switch.scala 41:52:@28616.4]
  assign output_31_10 = io_outValid_10 & _T_67457; // @[Switch.scala 41:38:@28617.4]
  assign _T_67460 = select_11 == 6'h1f; // @[Switch.scala 41:52:@28619.4]
  assign output_31_11 = io_outValid_11 & _T_67460; // @[Switch.scala 41:38:@28620.4]
  assign _T_67463 = select_12 == 6'h1f; // @[Switch.scala 41:52:@28622.4]
  assign output_31_12 = io_outValid_12 & _T_67463; // @[Switch.scala 41:38:@28623.4]
  assign _T_67466 = select_13 == 6'h1f; // @[Switch.scala 41:52:@28625.4]
  assign output_31_13 = io_outValid_13 & _T_67466; // @[Switch.scala 41:38:@28626.4]
  assign _T_67469 = select_14 == 6'h1f; // @[Switch.scala 41:52:@28628.4]
  assign output_31_14 = io_outValid_14 & _T_67469; // @[Switch.scala 41:38:@28629.4]
  assign _T_67472 = select_15 == 6'h1f; // @[Switch.scala 41:52:@28631.4]
  assign output_31_15 = io_outValid_15 & _T_67472; // @[Switch.scala 41:38:@28632.4]
  assign _T_67475 = select_16 == 6'h1f; // @[Switch.scala 41:52:@28634.4]
  assign output_31_16 = io_outValid_16 & _T_67475; // @[Switch.scala 41:38:@28635.4]
  assign _T_67478 = select_17 == 6'h1f; // @[Switch.scala 41:52:@28637.4]
  assign output_31_17 = io_outValid_17 & _T_67478; // @[Switch.scala 41:38:@28638.4]
  assign _T_67481 = select_18 == 6'h1f; // @[Switch.scala 41:52:@28640.4]
  assign output_31_18 = io_outValid_18 & _T_67481; // @[Switch.scala 41:38:@28641.4]
  assign _T_67484 = select_19 == 6'h1f; // @[Switch.scala 41:52:@28643.4]
  assign output_31_19 = io_outValid_19 & _T_67484; // @[Switch.scala 41:38:@28644.4]
  assign _T_67487 = select_20 == 6'h1f; // @[Switch.scala 41:52:@28646.4]
  assign output_31_20 = io_outValid_20 & _T_67487; // @[Switch.scala 41:38:@28647.4]
  assign _T_67490 = select_21 == 6'h1f; // @[Switch.scala 41:52:@28649.4]
  assign output_31_21 = io_outValid_21 & _T_67490; // @[Switch.scala 41:38:@28650.4]
  assign _T_67493 = select_22 == 6'h1f; // @[Switch.scala 41:52:@28652.4]
  assign output_31_22 = io_outValid_22 & _T_67493; // @[Switch.scala 41:38:@28653.4]
  assign _T_67496 = select_23 == 6'h1f; // @[Switch.scala 41:52:@28655.4]
  assign output_31_23 = io_outValid_23 & _T_67496; // @[Switch.scala 41:38:@28656.4]
  assign _T_67499 = select_24 == 6'h1f; // @[Switch.scala 41:52:@28658.4]
  assign output_31_24 = io_outValid_24 & _T_67499; // @[Switch.scala 41:38:@28659.4]
  assign _T_67502 = select_25 == 6'h1f; // @[Switch.scala 41:52:@28661.4]
  assign output_31_25 = io_outValid_25 & _T_67502; // @[Switch.scala 41:38:@28662.4]
  assign _T_67505 = select_26 == 6'h1f; // @[Switch.scala 41:52:@28664.4]
  assign output_31_26 = io_outValid_26 & _T_67505; // @[Switch.scala 41:38:@28665.4]
  assign _T_67508 = select_27 == 6'h1f; // @[Switch.scala 41:52:@28667.4]
  assign output_31_27 = io_outValid_27 & _T_67508; // @[Switch.scala 41:38:@28668.4]
  assign _T_67511 = select_28 == 6'h1f; // @[Switch.scala 41:52:@28670.4]
  assign output_31_28 = io_outValid_28 & _T_67511; // @[Switch.scala 41:38:@28671.4]
  assign _T_67514 = select_29 == 6'h1f; // @[Switch.scala 41:52:@28673.4]
  assign output_31_29 = io_outValid_29 & _T_67514; // @[Switch.scala 41:38:@28674.4]
  assign _T_67517 = select_30 == 6'h1f; // @[Switch.scala 41:52:@28676.4]
  assign output_31_30 = io_outValid_30 & _T_67517; // @[Switch.scala 41:38:@28677.4]
  assign _T_67520 = select_31 == 6'h1f; // @[Switch.scala 41:52:@28679.4]
  assign output_31_31 = io_outValid_31 & _T_67520; // @[Switch.scala 41:38:@28680.4]
  assign _T_67523 = select_32 == 6'h1f; // @[Switch.scala 41:52:@28682.4]
  assign output_31_32 = io_outValid_32 & _T_67523; // @[Switch.scala 41:38:@28683.4]
  assign _T_67526 = select_33 == 6'h1f; // @[Switch.scala 41:52:@28685.4]
  assign output_31_33 = io_outValid_33 & _T_67526; // @[Switch.scala 41:38:@28686.4]
  assign _T_67529 = select_34 == 6'h1f; // @[Switch.scala 41:52:@28688.4]
  assign output_31_34 = io_outValid_34 & _T_67529; // @[Switch.scala 41:38:@28689.4]
  assign _T_67532 = select_35 == 6'h1f; // @[Switch.scala 41:52:@28691.4]
  assign output_31_35 = io_outValid_35 & _T_67532; // @[Switch.scala 41:38:@28692.4]
  assign _T_67535 = select_36 == 6'h1f; // @[Switch.scala 41:52:@28694.4]
  assign output_31_36 = io_outValid_36 & _T_67535; // @[Switch.scala 41:38:@28695.4]
  assign _T_67538 = select_37 == 6'h1f; // @[Switch.scala 41:52:@28697.4]
  assign output_31_37 = io_outValid_37 & _T_67538; // @[Switch.scala 41:38:@28698.4]
  assign _T_67541 = select_38 == 6'h1f; // @[Switch.scala 41:52:@28700.4]
  assign output_31_38 = io_outValid_38 & _T_67541; // @[Switch.scala 41:38:@28701.4]
  assign _T_67544 = select_39 == 6'h1f; // @[Switch.scala 41:52:@28703.4]
  assign output_31_39 = io_outValid_39 & _T_67544; // @[Switch.scala 41:38:@28704.4]
  assign _T_67547 = select_40 == 6'h1f; // @[Switch.scala 41:52:@28706.4]
  assign output_31_40 = io_outValid_40 & _T_67547; // @[Switch.scala 41:38:@28707.4]
  assign _T_67550 = select_41 == 6'h1f; // @[Switch.scala 41:52:@28709.4]
  assign output_31_41 = io_outValid_41 & _T_67550; // @[Switch.scala 41:38:@28710.4]
  assign _T_67553 = select_42 == 6'h1f; // @[Switch.scala 41:52:@28712.4]
  assign output_31_42 = io_outValid_42 & _T_67553; // @[Switch.scala 41:38:@28713.4]
  assign _T_67556 = select_43 == 6'h1f; // @[Switch.scala 41:52:@28715.4]
  assign output_31_43 = io_outValid_43 & _T_67556; // @[Switch.scala 41:38:@28716.4]
  assign _T_67559 = select_44 == 6'h1f; // @[Switch.scala 41:52:@28718.4]
  assign output_31_44 = io_outValid_44 & _T_67559; // @[Switch.scala 41:38:@28719.4]
  assign _T_67562 = select_45 == 6'h1f; // @[Switch.scala 41:52:@28721.4]
  assign output_31_45 = io_outValid_45 & _T_67562; // @[Switch.scala 41:38:@28722.4]
  assign _T_67565 = select_46 == 6'h1f; // @[Switch.scala 41:52:@28724.4]
  assign output_31_46 = io_outValid_46 & _T_67565; // @[Switch.scala 41:38:@28725.4]
  assign _T_67568 = select_47 == 6'h1f; // @[Switch.scala 41:52:@28727.4]
  assign output_31_47 = io_outValid_47 & _T_67568; // @[Switch.scala 41:38:@28728.4]
  assign _T_67571 = select_48 == 6'h1f; // @[Switch.scala 41:52:@28730.4]
  assign output_31_48 = io_outValid_48 & _T_67571; // @[Switch.scala 41:38:@28731.4]
  assign _T_67574 = select_49 == 6'h1f; // @[Switch.scala 41:52:@28733.4]
  assign output_31_49 = io_outValid_49 & _T_67574; // @[Switch.scala 41:38:@28734.4]
  assign _T_67577 = select_50 == 6'h1f; // @[Switch.scala 41:52:@28736.4]
  assign output_31_50 = io_outValid_50 & _T_67577; // @[Switch.scala 41:38:@28737.4]
  assign _T_67580 = select_51 == 6'h1f; // @[Switch.scala 41:52:@28739.4]
  assign output_31_51 = io_outValid_51 & _T_67580; // @[Switch.scala 41:38:@28740.4]
  assign _T_67583 = select_52 == 6'h1f; // @[Switch.scala 41:52:@28742.4]
  assign output_31_52 = io_outValid_52 & _T_67583; // @[Switch.scala 41:38:@28743.4]
  assign _T_67586 = select_53 == 6'h1f; // @[Switch.scala 41:52:@28745.4]
  assign output_31_53 = io_outValid_53 & _T_67586; // @[Switch.scala 41:38:@28746.4]
  assign _T_67589 = select_54 == 6'h1f; // @[Switch.scala 41:52:@28748.4]
  assign output_31_54 = io_outValid_54 & _T_67589; // @[Switch.scala 41:38:@28749.4]
  assign _T_67592 = select_55 == 6'h1f; // @[Switch.scala 41:52:@28751.4]
  assign output_31_55 = io_outValid_55 & _T_67592; // @[Switch.scala 41:38:@28752.4]
  assign _T_67595 = select_56 == 6'h1f; // @[Switch.scala 41:52:@28754.4]
  assign output_31_56 = io_outValid_56 & _T_67595; // @[Switch.scala 41:38:@28755.4]
  assign _T_67598 = select_57 == 6'h1f; // @[Switch.scala 41:52:@28757.4]
  assign output_31_57 = io_outValid_57 & _T_67598; // @[Switch.scala 41:38:@28758.4]
  assign _T_67601 = select_58 == 6'h1f; // @[Switch.scala 41:52:@28760.4]
  assign output_31_58 = io_outValid_58 & _T_67601; // @[Switch.scala 41:38:@28761.4]
  assign _T_67604 = select_59 == 6'h1f; // @[Switch.scala 41:52:@28763.4]
  assign output_31_59 = io_outValid_59 & _T_67604; // @[Switch.scala 41:38:@28764.4]
  assign _T_67607 = select_60 == 6'h1f; // @[Switch.scala 41:52:@28766.4]
  assign output_31_60 = io_outValid_60 & _T_67607; // @[Switch.scala 41:38:@28767.4]
  assign _T_67610 = select_61 == 6'h1f; // @[Switch.scala 41:52:@28769.4]
  assign output_31_61 = io_outValid_61 & _T_67610; // @[Switch.scala 41:38:@28770.4]
  assign _T_67613 = select_62 == 6'h1f; // @[Switch.scala 41:52:@28772.4]
  assign output_31_62 = io_outValid_62 & _T_67613; // @[Switch.scala 41:38:@28773.4]
  assign _T_67616 = select_63 == 6'h1f; // @[Switch.scala 41:52:@28775.4]
  assign output_31_63 = io_outValid_63 & _T_67616; // @[Switch.scala 41:38:@28776.4]
  assign _T_67624 = {output_31_7,output_31_6,output_31_5,output_31_4,output_31_3,output_31_2,output_31_1,output_31_0}; // @[Switch.scala 43:31:@28784.4]
  assign _T_67632 = {output_31_15,output_31_14,output_31_13,output_31_12,output_31_11,output_31_10,output_31_9,output_31_8,_T_67624}; // @[Switch.scala 43:31:@28792.4]
  assign _T_67639 = {output_31_23,output_31_22,output_31_21,output_31_20,output_31_19,output_31_18,output_31_17,output_31_16}; // @[Switch.scala 43:31:@28799.4]
  assign _T_67648 = {output_31_31,output_31_30,output_31_29,output_31_28,output_31_27,output_31_26,output_31_25,output_31_24,_T_67639,_T_67632}; // @[Switch.scala 43:31:@28808.4]
  assign _T_67655 = {output_31_39,output_31_38,output_31_37,output_31_36,output_31_35,output_31_34,output_31_33,output_31_32}; // @[Switch.scala 43:31:@28815.4]
  assign _T_67663 = {output_31_47,output_31_46,output_31_45,output_31_44,output_31_43,output_31_42,output_31_41,output_31_40,_T_67655}; // @[Switch.scala 43:31:@28823.4]
  assign _T_67670 = {output_31_55,output_31_54,output_31_53,output_31_52,output_31_51,output_31_50,output_31_49,output_31_48}; // @[Switch.scala 43:31:@28830.4]
  assign _T_67679 = {output_31_63,output_31_62,output_31_61,output_31_60,output_31_59,output_31_58,output_31_57,output_31_56,_T_67670,_T_67663}; // @[Switch.scala 43:31:@28839.4]
  assign _T_67680 = {_T_67679,_T_67648}; // @[Switch.scala 43:31:@28840.4]
  assign _T_67684 = select_0 == 6'h20; // @[Switch.scala 41:52:@28843.4]
  assign output_32_0 = io_outValid_0 & _T_67684; // @[Switch.scala 41:38:@28844.4]
  assign _T_67687 = select_1 == 6'h20; // @[Switch.scala 41:52:@28846.4]
  assign output_32_1 = io_outValid_1 & _T_67687; // @[Switch.scala 41:38:@28847.4]
  assign _T_67690 = select_2 == 6'h20; // @[Switch.scala 41:52:@28849.4]
  assign output_32_2 = io_outValid_2 & _T_67690; // @[Switch.scala 41:38:@28850.4]
  assign _T_67693 = select_3 == 6'h20; // @[Switch.scala 41:52:@28852.4]
  assign output_32_3 = io_outValid_3 & _T_67693; // @[Switch.scala 41:38:@28853.4]
  assign _T_67696 = select_4 == 6'h20; // @[Switch.scala 41:52:@28855.4]
  assign output_32_4 = io_outValid_4 & _T_67696; // @[Switch.scala 41:38:@28856.4]
  assign _T_67699 = select_5 == 6'h20; // @[Switch.scala 41:52:@28858.4]
  assign output_32_5 = io_outValid_5 & _T_67699; // @[Switch.scala 41:38:@28859.4]
  assign _T_67702 = select_6 == 6'h20; // @[Switch.scala 41:52:@28861.4]
  assign output_32_6 = io_outValid_6 & _T_67702; // @[Switch.scala 41:38:@28862.4]
  assign _T_67705 = select_7 == 6'h20; // @[Switch.scala 41:52:@28864.4]
  assign output_32_7 = io_outValid_7 & _T_67705; // @[Switch.scala 41:38:@28865.4]
  assign _T_67708 = select_8 == 6'h20; // @[Switch.scala 41:52:@28867.4]
  assign output_32_8 = io_outValid_8 & _T_67708; // @[Switch.scala 41:38:@28868.4]
  assign _T_67711 = select_9 == 6'h20; // @[Switch.scala 41:52:@28870.4]
  assign output_32_9 = io_outValid_9 & _T_67711; // @[Switch.scala 41:38:@28871.4]
  assign _T_67714 = select_10 == 6'h20; // @[Switch.scala 41:52:@28873.4]
  assign output_32_10 = io_outValid_10 & _T_67714; // @[Switch.scala 41:38:@28874.4]
  assign _T_67717 = select_11 == 6'h20; // @[Switch.scala 41:52:@28876.4]
  assign output_32_11 = io_outValid_11 & _T_67717; // @[Switch.scala 41:38:@28877.4]
  assign _T_67720 = select_12 == 6'h20; // @[Switch.scala 41:52:@28879.4]
  assign output_32_12 = io_outValid_12 & _T_67720; // @[Switch.scala 41:38:@28880.4]
  assign _T_67723 = select_13 == 6'h20; // @[Switch.scala 41:52:@28882.4]
  assign output_32_13 = io_outValid_13 & _T_67723; // @[Switch.scala 41:38:@28883.4]
  assign _T_67726 = select_14 == 6'h20; // @[Switch.scala 41:52:@28885.4]
  assign output_32_14 = io_outValid_14 & _T_67726; // @[Switch.scala 41:38:@28886.4]
  assign _T_67729 = select_15 == 6'h20; // @[Switch.scala 41:52:@28888.4]
  assign output_32_15 = io_outValid_15 & _T_67729; // @[Switch.scala 41:38:@28889.4]
  assign _T_67732 = select_16 == 6'h20; // @[Switch.scala 41:52:@28891.4]
  assign output_32_16 = io_outValid_16 & _T_67732; // @[Switch.scala 41:38:@28892.4]
  assign _T_67735 = select_17 == 6'h20; // @[Switch.scala 41:52:@28894.4]
  assign output_32_17 = io_outValid_17 & _T_67735; // @[Switch.scala 41:38:@28895.4]
  assign _T_67738 = select_18 == 6'h20; // @[Switch.scala 41:52:@28897.4]
  assign output_32_18 = io_outValid_18 & _T_67738; // @[Switch.scala 41:38:@28898.4]
  assign _T_67741 = select_19 == 6'h20; // @[Switch.scala 41:52:@28900.4]
  assign output_32_19 = io_outValid_19 & _T_67741; // @[Switch.scala 41:38:@28901.4]
  assign _T_67744 = select_20 == 6'h20; // @[Switch.scala 41:52:@28903.4]
  assign output_32_20 = io_outValid_20 & _T_67744; // @[Switch.scala 41:38:@28904.4]
  assign _T_67747 = select_21 == 6'h20; // @[Switch.scala 41:52:@28906.4]
  assign output_32_21 = io_outValid_21 & _T_67747; // @[Switch.scala 41:38:@28907.4]
  assign _T_67750 = select_22 == 6'h20; // @[Switch.scala 41:52:@28909.4]
  assign output_32_22 = io_outValid_22 & _T_67750; // @[Switch.scala 41:38:@28910.4]
  assign _T_67753 = select_23 == 6'h20; // @[Switch.scala 41:52:@28912.4]
  assign output_32_23 = io_outValid_23 & _T_67753; // @[Switch.scala 41:38:@28913.4]
  assign _T_67756 = select_24 == 6'h20; // @[Switch.scala 41:52:@28915.4]
  assign output_32_24 = io_outValid_24 & _T_67756; // @[Switch.scala 41:38:@28916.4]
  assign _T_67759 = select_25 == 6'h20; // @[Switch.scala 41:52:@28918.4]
  assign output_32_25 = io_outValid_25 & _T_67759; // @[Switch.scala 41:38:@28919.4]
  assign _T_67762 = select_26 == 6'h20; // @[Switch.scala 41:52:@28921.4]
  assign output_32_26 = io_outValid_26 & _T_67762; // @[Switch.scala 41:38:@28922.4]
  assign _T_67765 = select_27 == 6'h20; // @[Switch.scala 41:52:@28924.4]
  assign output_32_27 = io_outValid_27 & _T_67765; // @[Switch.scala 41:38:@28925.4]
  assign _T_67768 = select_28 == 6'h20; // @[Switch.scala 41:52:@28927.4]
  assign output_32_28 = io_outValid_28 & _T_67768; // @[Switch.scala 41:38:@28928.4]
  assign _T_67771 = select_29 == 6'h20; // @[Switch.scala 41:52:@28930.4]
  assign output_32_29 = io_outValid_29 & _T_67771; // @[Switch.scala 41:38:@28931.4]
  assign _T_67774 = select_30 == 6'h20; // @[Switch.scala 41:52:@28933.4]
  assign output_32_30 = io_outValid_30 & _T_67774; // @[Switch.scala 41:38:@28934.4]
  assign _T_67777 = select_31 == 6'h20; // @[Switch.scala 41:52:@28936.4]
  assign output_32_31 = io_outValid_31 & _T_67777; // @[Switch.scala 41:38:@28937.4]
  assign _T_67780 = select_32 == 6'h20; // @[Switch.scala 41:52:@28939.4]
  assign output_32_32 = io_outValid_32 & _T_67780; // @[Switch.scala 41:38:@28940.4]
  assign _T_67783 = select_33 == 6'h20; // @[Switch.scala 41:52:@28942.4]
  assign output_32_33 = io_outValid_33 & _T_67783; // @[Switch.scala 41:38:@28943.4]
  assign _T_67786 = select_34 == 6'h20; // @[Switch.scala 41:52:@28945.4]
  assign output_32_34 = io_outValid_34 & _T_67786; // @[Switch.scala 41:38:@28946.4]
  assign _T_67789 = select_35 == 6'h20; // @[Switch.scala 41:52:@28948.4]
  assign output_32_35 = io_outValid_35 & _T_67789; // @[Switch.scala 41:38:@28949.4]
  assign _T_67792 = select_36 == 6'h20; // @[Switch.scala 41:52:@28951.4]
  assign output_32_36 = io_outValid_36 & _T_67792; // @[Switch.scala 41:38:@28952.4]
  assign _T_67795 = select_37 == 6'h20; // @[Switch.scala 41:52:@28954.4]
  assign output_32_37 = io_outValid_37 & _T_67795; // @[Switch.scala 41:38:@28955.4]
  assign _T_67798 = select_38 == 6'h20; // @[Switch.scala 41:52:@28957.4]
  assign output_32_38 = io_outValid_38 & _T_67798; // @[Switch.scala 41:38:@28958.4]
  assign _T_67801 = select_39 == 6'h20; // @[Switch.scala 41:52:@28960.4]
  assign output_32_39 = io_outValid_39 & _T_67801; // @[Switch.scala 41:38:@28961.4]
  assign _T_67804 = select_40 == 6'h20; // @[Switch.scala 41:52:@28963.4]
  assign output_32_40 = io_outValid_40 & _T_67804; // @[Switch.scala 41:38:@28964.4]
  assign _T_67807 = select_41 == 6'h20; // @[Switch.scala 41:52:@28966.4]
  assign output_32_41 = io_outValid_41 & _T_67807; // @[Switch.scala 41:38:@28967.4]
  assign _T_67810 = select_42 == 6'h20; // @[Switch.scala 41:52:@28969.4]
  assign output_32_42 = io_outValid_42 & _T_67810; // @[Switch.scala 41:38:@28970.4]
  assign _T_67813 = select_43 == 6'h20; // @[Switch.scala 41:52:@28972.4]
  assign output_32_43 = io_outValid_43 & _T_67813; // @[Switch.scala 41:38:@28973.4]
  assign _T_67816 = select_44 == 6'h20; // @[Switch.scala 41:52:@28975.4]
  assign output_32_44 = io_outValid_44 & _T_67816; // @[Switch.scala 41:38:@28976.4]
  assign _T_67819 = select_45 == 6'h20; // @[Switch.scala 41:52:@28978.4]
  assign output_32_45 = io_outValid_45 & _T_67819; // @[Switch.scala 41:38:@28979.4]
  assign _T_67822 = select_46 == 6'h20; // @[Switch.scala 41:52:@28981.4]
  assign output_32_46 = io_outValid_46 & _T_67822; // @[Switch.scala 41:38:@28982.4]
  assign _T_67825 = select_47 == 6'h20; // @[Switch.scala 41:52:@28984.4]
  assign output_32_47 = io_outValid_47 & _T_67825; // @[Switch.scala 41:38:@28985.4]
  assign _T_67828 = select_48 == 6'h20; // @[Switch.scala 41:52:@28987.4]
  assign output_32_48 = io_outValid_48 & _T_67828; // @[Switch.scala 41:38:@28988.4]
  assign _T_67831 = select_49 == 6'h20; // @[Switch.scala 41:52:@28990.4]
  assign output_32_49 = io_outValid_49 & _T_67831; // @[Switch.scala 41:38:@28991.4]
  assign _T_67834 = select_50 == 6'h20; // @[Switch.scala 41:52:@28993.4]
  assign output_32_50 = io_outValid_50 & _T_67834; // @[Switch.scala 41:38:@28994.4]
  assign _T_67837 = select_51 == 6'h20; // @[Switch.scala 41:52:@28996.4]
  assign output_32_51 = io_outValid_51 & _T_67837; // @[Switch.scala 41:38:@28997.4]
  assign _T_67840 = select_52 == 6'h20; // @[Switch.scala 41:52:@28999.4]
  assign output_32_52 = io_outValid_52 & _T_67840; // @[Switch.scala 41:38:@29000.4]
  assign _T_67843 = select_53 == 6'h20; // @[Switch.scala 41:52:@29002.4]
  assign output_32_53 = io_outValid_53 & _T_67843; // @[Switch.scala 41:38:@29003.4]
  assign _T_67846 = select_54 == 6'h20; // @[Switch.scala 41:52:@29005.4]
  assign output_32_54 = io_outValid_54 & _T_67846; // @[Switch.scala 41:38:@29006.4]
  assign _T_67849 = select_55 == 6'h20; // @[Switch.scala 41:52:@29008.4]
  assign output_32_55 = io_outValid_55 & _T_67849; // @[Switch.scala 41:38:@29009.4]
  assign _T_67852 = select_56 == 6'h20; // @[Switch.scala 41:52:@29011.4]
  assign output_32_56 = io_outValid_56 & _T_67852; // @[Switch.scala 41:38:@29012.4]
  assign _T_67855 = select_57 == 6'h20; // @[Switch.scala 41:52:@29014.4]
  assign output_32_57 = io_outValid_57 & _T_67855; // @[Switch.scala 41:38:@29015.4]
  assign _T_67858 = select_58 == 6'h20; // @[Switch.scala 41:52:@29017.4]
  assign output_32_58 = io_outValid_58 & _T_67858; // @[Switch.scala 41:38:@29018.4]
  assign _T_67861 = select_59 == 6'h20; // @[Switch.scala 41:52:@29020.4]
  assign output_32_59 = io_outValid_59 & _T_67861; // @[Switch.scala 41:38:@29021.4]
  assign _T_67864 = select_60 == 6'h20; // @[Switch.scala 41:52:@29023.4]
  assign output_32_60 = io_outValid_60 & _T_67864; // @[Switch.scala 41:38:@29024.4]
  assign _T_67867 = select_61 == 6'h20; // @[Switch.scala 41:52:@29026.4]
  assign output_32_61 = io_outValid_61 & _T_67867; // @[Switch.scala 41:38:@29027.4]
  assign _T_67870 = select_62 == 6'h20; // @[Switch.scala 41:52:@29029.4]
  assign output_32_62 = io_outValid_62 & _T_67870; // @[Switch.scala 41:38:@29030.4]
  assign _T_67873 = select_63 == 6'h20; // @[Switch.scala 41:52:@29032.4]
  assign output_32_63 = io_outValid_63 & _T_67873; // @[Switch.scala 41:38:@29033.4]
  assign _T_67881 = {output_32_7,output_32_6,output_32_5,output_32_4,output_32_3,output_32_2,output_32_1,output_32_0}; // @[Switch.scala 43:31:@29041.4]
  assign _T_67889 = {output_32_15,output_32_14,output_32_13,output_32_12,output_32_11,output_32_10,output_32_9,output_32_8,_T_67881}; // @[Switch.scala 43:31:@29049.4]
  assign _T_67896 = {output_32_23,output_32_22,output_32_21,output_32_20,output_32_19,output_32_18,output_32_17,output_32_16}; // @[Switch.scala 43:31:@29056.4]
  assign _T_67905 = {output_32_31,output_32_30,output_32_29,output_32_28,output_32_27,output_32_26,output_32_25,output_32_24,_T_67896,_T_67889}; // @[Switch.scala 43:31:@29065.4]
  assign _T_67912 = {output_32_39,output_32_38,output_32_37,output_32_36,output_32_35,output_32_34,output_32_33,output_32_32}; // @[Switch.scala 43:31:@29072.4]
  assign _T_67920 = {output_32_47,output_32_46,output_32_45,output_32_44,output_32_43,output_32_42,output_32_41,output_32_40,_T_67912}; // @[Switch.scala 43:31:@29080.4]
  assign _T_67927 = {output_32_55,output_32_54,output_32_53,output_32_52,output_32_51,output_32_50,output_32_49,output_32_48}; // @[Switch.scala 43:31:@29087.4]
  assign _T_67936 = {output_32_63,output_32_62,output_32_61,output_32_60,output_32_59,output_32_58,output_32_57,output_32_56,_T_67927,_T_67920}; // @[Switch.scala 43:31:@29096.4]
  assign _T_67937 = {_T_67936,_T_67905}; // @[Switch.scala 43:31:@29097.4]
  assign _T_67941 = select_0 == 6'h21; // @[Switch.scala 41:52:@29100.4]
  assign output_33_0 = io_outValid_0 & _T_67941; // @[Switch.scala 41:38:@29101.4]
  assign _T_67944 = select_1 == 6'h21; // @[Switch.scala 41:52:@29103.4]
  assign output_33_1 = io_outValid_1 & _T_67944; // @[Switch.scala 41:38:@29104.4]
  assign _T_67947 = select_2 == 6'h21; // @[Switch.scala 41:52:@29106.4]
  assign output_33_2 = io_outValid_2 & _T_67947; // @[Switch.scala 41:38:@29107.4]
  assign _T_67950 = select_3 == 6'h21; // @[Switch.scala 41:52:@29109.4]
  assign output_33_3 = io_outValid_3 & _T_67950; // @[Switch.scala 41:38:@29110.4]
  assign _T_67953 = select_4 == 6'h21; // @[Switch.scala 41:52:@29112.4]
  assign output_33_4 = io_outValid_4 & _T_67953; // @[Switch.scala 41:38:@29113.4]
  assign _T_67956 = select_5 == 6'h21; // @[Switch.scala 41:52:@29115.4]
  assign output_33_5 = io_outValid_5 & _T_67956; // @[Switch.scala 41:38:@29116.4]
  assign _T_67959 = select_6 == 6'h21; // @[Switch.scala 41:52:@29118.4]
  assign output_33_6 = io_outValid_6 & _T_67959; // @[Switch.scala 41:38:@29119.4]
  assign _T_67962 = select_7 == 6'h21; // @[Switch.scala 41:52:@29121.4]
  assign output_33_7 = io_outValid_7 & _T_67962; // @[Switch.scala 41:38:@29122.4]
  assign _T_67965 = select_8 == 6'h21; // @[Switch.scala 41:52:@29124.4]
  assign output_33_8 = io_outValid_8 & _T_67965; // @[Switch.scala 41:38:@29125.4]
  assign _T_67968 = select_9 == 6'h21; // @[Switch.scala 41:52:@29127.4]
  assign output_33_9 = io_outValid_9 & _T_67968; // @[Switch.scala 41:38:@29128.4]
  assign _T_67971 = select_10 == 6'h21; // @[Switch.scala 41:52:@29130.4]
  assign output_33_10 = io_outValid_10 & _T_67971; // @[Switch.scala 41:38:@29131.4]
  assign _T_67974 = select_11 == 6'h21; // @[Switch.scala 41:52:@29133.4]
  assign output_33_11 = io_outValid_11 & _T_67974; // @[Switch.scala 41:38:@29134.4]
  assign _T_67977 = select_12 == 6'h21; // @[Switch.scala 41:52:@29136.4]
  assign output_33_12 = io_outValid_12 & _T_67977; // @[Switch.scala 41:38:@29137.4]
  assign _T_67980 = select_13 == 6'h21; // @[Switch.scala 41:52:@29139.4]
  assign output_33_13 = io_outValid_13 & _T_67980; // @[Switch.scala 41:38:@29140.4]
  assign _T_67983 = select_14 == 6'h21; // @[Switch.scala 41:52:@29142.4]
  assign output_33_14 = io_outValid_14 & _T_67983; // @[Switch.scala 41:38:@29143.4]
  assign _T_67986 = select_15 == 6'h21; // @[Switch.scala 41:52:@29145.4]
  assign output_33_15 = io_outValid_15 & _T_67986; // @[Switch.scala 41:38:@29146.4]
  assign _T_67989 = select_16 == 6'h21; // @[Switch.scala 41:52:@29148.4]
  assign output_33_16 = io_outValid_16 & _T_67989; // @[Switch.scala 41:38:@29149.4]
  assign _T_67992 = select_17 == 6'h21; // @[Switch.scala 41:52:@29151.4]
  assign output_33_17 = io_outValid_17 & _T_67992; // @[Switch.scala 41:38:@29152.4]
  assign _T_67995 = select_18 == 6'h21; // @[Switch.scala 41:52:@29154.4]
  assign output_33_18 = io_outValid_18 & _T_67995; // @[Switch.scala 41:38:@29155.4]
  assign _T_67998 = select_19 == 6'h21; // @[Switch.scala 41:52:@29157.4]
  assign output_33_19 = io_outValid_19 & _T_67998; // @[Switch.scala 41:38:@29158.4]
  assign _T_68001 = select_20 == 6'h21; // @[Switch.scala 41:52:@29160.4]
  assign output_33_20 = io_outValid_20 & _T_68001; // @[Switch.scala 41:38:@29161.4]
  assign _T_68004 = select_21 == 6'h21; // @[Switch.scala 41:52:@29163.4]
  assign output_33_21 = io_outValid_21 & _T_68004; // @[Switch.scala 41:38:@29164.4]
  assign _T_68007 = select_22 == 6'h21; // @[Switch.scala 41:52:@29166.4]
  assign output_33_22 = io_outValid_22 & _T_68007; // @[Switch.scala 41:38:@29167.4]
  assign _T_68010 = select_23 == 6'h21; // @[Switch.scala 41:52:@29169.4]
  assign output_33_23 = io_outValid_23 & _T_68010; // @[Switch.scala 41:38:@29170.4]
  assign _T_68013 = select_24 == 6'h21; // @[Switch.scala 41:52:@29172.4]
  assign output_33_24 = io_outValid_24 & _T_68013; // @[Switch.scala 41:38:@29173.4]
  assign _T_68016 = select_25 == 6'h21; // @[Switch.scala 41:52:@29175.4]
  assign output_33_25 = io_outValid_25 & _T_68016; // @[Switch.scala 41:38:@29176.4]
  assign _T_68019 = select_26 == 6'h21; // @[Switch.scala 41:52:@29178.4]
  assign output_33_26 = io_outValid_26 & _T_68019; // @[Switch.scala 41:38:@29179.4]
  assign _T_68022 = select_27 == 6'h21; // @[Switch.scala 41:52:@29181.4]
  assign output_33_27 = io_outValid_27 & _T_68022; // @[Switch.scala 41:38:@29182.4]
  assign _T_68025 = select_28 == 6'h21; // @[Switch.scala 41:52:@29184.4]
  assign output_33_28 = io_outValid_28 & _T_68025; // @[Switch.scala 41:38:@29185.4]
  assign _T_68028 = select_29 == 6'h21; // @[Switch.scala 41:52:@29187.4]
  assign output_33_29 = io_outValid_29 & _T_68028; // @[Switch.scala 41:38:@29188.4]
  assign _T_68031 = select_30 == 6'h21; // @[Switch.scala 41:52:@29190.4]
  assign output_33_30 = io_outValid_30 & _T_68031; // @[Switch.scala 41:38:@29191.4]
  assign _T_68034 = select_31 == 6'h21; // @[Switch.scala 41:52:@29193.4]
  assign output_33_31 = io_outValid_31 & _T_68034; // @[Switch.scala 41:38:@29194.4]
  assign _T_68037 = select_32 == 6'h21; // @[Switch.scala 41:52:@29196.4]
  assign output_33_32 = io_outValid_32 & _T_68037; // @[Switch.scala 41:38:@29197.4]
  assign _T_68040 = select_33 == 6'h21; // @[Switch.scala 41:52:@29199.4]
  assign output_33_33 = io_outValid_33 & _T_68040; // @[Switch.scala 41:38:@29200.4]
  assign _T_68043 = select_34 == 6'h21; // @[Switch.scala 41:52:@29202.4]
  assign output_33_34 = io_outValid_34 & _T_68043; // @[Switch.scala 41:38:@29203.4]
  assign _T_68046 = select_35 == 6'h21; // @[Switch.scala 41:52:@29205.4]
  assign output_33_35 = io_outValid_35 & _T_68046; // @[Switch.scala 41:38:@29206.4]
  assign _T_68049 = select_36 == 6'h21; // @[Switch.scala 41:52:@29208.4]
  assign output_33_36 = io_outValid_36 & _T_68049; // @[Switch.scala 41:38:@29209.4]
  assign _T_68052 = select_37 == 6'h21; // @[Switch.scala 41:52:@29211.4]
  assign output_33_37 = io_outValid_37 & _T_68052; // @[Switch.scala 41:38:@29212.4]
  assign _T_68055 = select_38 == 6'h21; // @[Switch.scala 41:52:@29214.4]
  assign output_33_38 = io_outValid_38 & _T_68055; // @[Switch.scala 41:38:@29215.4]
  assign _T_68058 = select_39 == 6'h21; // @[Switch.scala 41:52:@29217.4]
  assign output_33_39 = io_outValid_39 & _T_68058; // @[Switch.scala 41:38:@29218.4]
  assign _T_68061 = select_40 == 6'h21; // @[Switch.scala 41:52:@29220.4]
  assign output_33_40 = io_outValid_40 & _T_68061; // @[Switch.scala 41:38:@29221.4]
  assign _T_68064 = select_41 == 6'h21; // @[Switch.scala 41:52:@29223.4]
  assign output_33_41 = io_outValid_41 & _T_68064; // @[Switch.scala 41:38:@29224.4]
  assign _T_68067 = select_42 == 6'h21; // @[Switch.scala 41:52:@29226.4]
  assign output_33_42 = io_outValid_42 & _T_68067; // @[Switch.scala 41:38:@29227.4]
  assign _T_68070 = select_43 == 6'h21; // @[Switch.scala 41:52:@29229.4]
  assign output_33_43 = io_outValid_43 & _T_68070; // @[Switch.scala 41:38:@29230.4]
  assign _T_68073 = select_44 == 6'h21; // @[Switch.scala 41:52:@29232.4]
  assign output_33_44 = io_outValid_44 & _T_68073; // @[Switch.scala 41:38:@29233.4]
  assign _T_68076 = select_45 == 6'h21; // @[Switch.scala 41:52:@29235.4]
  assign output_33_45 = io_outValid_45 & _T_68076; // @[Switch.scala 41:38:@29236.4]
  assign _T_68079 = select_46 == 6'h21; // @[Switch.scala 41:52:@29238.4]
  assign output_33_46 = io_outValid_46 & _T_68079; // @[Switch.scala 41:38:@29239.4]
  assign _T_68082 = select_47 == 6'h21; // @[Switch.scala 41:52:@29241.4]
  assign output_33_47 = io_outValid_47 & _T_68082; // @[Switch.scala 41:38:@29242.4]
  assign _T_68085 = select_48 == 6'h21; // @[Switch.scala 41:52:@29244.4]
  assign output_33_48 = io_outValid_48 & _T_68085; // @[Switch.scala 41:38:@29245.4]
  assign _T_68088 = select_49 == 6'h21; // @[Switch.scala 41:52:@29247.4]
  assign output_33_49 = io_outValid_49 & _T_68088; // @[Switch.scala 41:38:@29248.4]
  assign _T_68091 = select_50 == 6'h21; // @[Switch.scala 41:52:@29250.4]
  assign output_33_50 = io_outValid_50 & _T_68091; // @[Switch.scala 41:38:@29251.4]
  assign _T_68094 = select_51 == 6'h21; // @[Switch.scala 41:52:@29253.4]
  assign output_33_51 = io_outValid_51 & _T_68094; // @[Switch.scala 41:38:@29254.4]
  assign _T_68097 = select_52 == 6'h21; // @[Switch.scala 41:52:@29256.4]
  assign output_33_52 = io_outValid_52 & _T_68097; // @[Switch.scala 41:38:@29257.4]
  assign _T_68100 = select_53 == 6'h21; // @[Switch.scala 41:52:@29259.4]
  assign output_33_53 = io_outValid_53 & _T_68100; // @[Switch.scala 41:38:@29260.4]
  assign _T_68103 = select_54 == 6'h21; // @[Switch.scala 41:52:@29262.4]
  assign output_33_54 = io_outValid_54 & _T_68103; // @[Switch.scala 41:38:@29263.4]
  assign _T_68106 = select_55 == 6'h21; // @[Switch.scala 41:52:@29265.4]
  assign output_33_55 = io_outValid_55 & _T_68106; // @[Switch.scala 41:38:@29266.4]
  assign _T_68109 = select_56 == 6'h21; // @[Switch.scala 41:52:@29268.4]
  assign output_33_56 = io_outValid_56 & _T_68109; // @[Switch.scala 41:38:@29269.4]
  assign _T_68112 = select_57 == 6'h21; // @[Switch.scala 41:52:@29271.4]
  assign output_33_57 = io_outValid_57 & _T_68112; // @[Switch.scala 41:38:@29272.4]
  assign _T_68115 = select_58 == 6'h21; // @[Switch.scala 41:52:@29274.4]
  assign output_33_58 = io_outValid_58 & _T_68115; // @[Switch.scala 41:38:@29275.4]
  assign _T_68118 = select_59 == 6'h21; // @[Switch.scala 41:52:@29277.4]
  assign output_33_59 = io_outValid_59 & _T_68118; // @[Switch.scala 41:38:@29278.4]
  assign _T_68121 = select_60 == 6'h21; // @[Switch.scala 41:52:@29280.4]
  assign output_33_60 = io_outValid_60 & _T_68121; // @[Switch.scala 41:38:@29281.4]
  assign _T_68124 = select_61 == 6'h21; // @[Switch.scala 41:52:@29283.4]
  assign output_33_61 = io_outValid_61 & _T_68124; // @[Switch.scala 41:38:@29284.4]
  assign _T_68127 = select_62 == 6'h21; // @[Switch.scala 41:52:@29286.4]
  assign output_33_62 = io_outValid_62 & _T_68127; // @[Switch.scala 41:38:@29287.4]
  assign _T_68130 = select_63 == 6'h21; // @[Switch.scala 41:52:@29289.4]
  assign output_33_63 = io_outValid_63 & _T_68130; // @[Switch.scala 41:38:@29290.4]
  assign _T_68138 = {output_33_7,output_33_6,output_33_5,output_33_4,output_33_3,output_33_2,output_33_1,output_33_0}; // @[Switch.scala 43:31:@29298.4]
  assign _T_68146 = {output_33_15,output_33_14,output_33_13,output_33_12,output_33_11,output_33_10,output_33_9,output_33_8,_T_68138}; // @[Switch.scala 43:31:@29306.4]
  assign _T_68153 = {output_33_23,output_33_22,output_33_21,output_33_20,output_33_19,output_33_18,output_33_17,output_33_16}; // @[Switch.scala 43:31:@29313.4]
  assign _T_68162 = {output_33_31,output_33_30,output_33_29,output_33_28,output_33_27,output_33_26,output_33_25,output_33_24,_T_68153,_T_68146}; // @[Switch.scala 43:31:@29322.4]
  assign _T_68169 = {output_33_39,output_33_38,output_33_37,output_33_36,output_33_35,output_33_34,output_33_33,output_33_32}; // @[Switch.scala 43:31:@29329.4]
  assign _T_68177 = {output_33_47,output_33_46,output_33_45,output_33_44,output_33_43,output_33_42,output_33_41,output_33_40,_T_68169}; // @[Switch.scala 43:31:@29337.4]
  assign _T_68184 = {output_33_55,output_33_54,output_33_53,output_33_52,output_33_51,output_33_50,output_33_49,output_33_48}; // @[Switch.scala 43:31:@29344.4]
  assign _T_68193 = {output_33_63,output_33_62,output_33_61,output_33_60,output_33_59,output_33_58,output_33_57,output_33_56,_T_68184,_T_68177}; // @[Switch.scala 43:31:@29353.4]
  assign _T_68194 = {_T_68193,_T_68162}; // @[Switch.scala 43:31:@29354.4]
  assign _T_68198 = select_0 == 6'h22; // @[Switch.scala 41:52:@29357.4]
  assign output_34_0 = io_outValid_0 & _T_68198; // @[Switch.scala 41:38:@29358.4]
  assign _T_68201 = select_1 == 6'h22; // @[Switch.scala 41:52:@29360.4]
  assign output_34_1 = io_outValid_1 & _T_68201; // @[Switch.scala 41:38:@29361.4]
  assign _T_68204 = select_2 == 6'h22; // @[Switch.scala 41:52:@29363.4]
  assign output_34_2 = io_outValid_2 & _T_68204; // @[Switch.scala 41:38:@29364.4]
  assign _T_68207 = select_3 == 6'h22; // @[Switch.scala 41:52:@29366.4]
  assign output_34_3 = io_outValid_3 & _T_68207; // @[Switch.scala 41:38:@29367.4]
  assign _T_68210 = select_4 == 6'h22; // @[Switch.scala 41:52:@29369.4]
  assign output_34_4 = io_outValid_4 & _T_68210; // @[Switch.scala 41:38:@29370.4]
  assign _T_68213 = select_5 == 6'h22; // @[Switch.scala 41:52:@29372.4]
  assign output_34_5 = io_outValid_5 & _T_68213; // @[Switch.scala 41:38:@29373.4]
  assign _T_68216 = select_6 == 6'h22; // @[Switch.scala 41:52:@29375.4]
  assign output_34_6 = io_outValid_6 & _T_68216; // @[Switch.scala 41:38:@29376.4]
  assign _T_68219 = select_7 == 6'h22; // @[Switch.scala 41:52:@29378.4]
  assign output_34_7 = io_outValid_7 & _T_68219; // @[Switch.scala 41:38:@29379.4]
  assign _T_68222 = select_8 == 6'h22; // @[Switch.scala 41:52:@29381.4]
  assign output_34_8 = io_outValid_8 & _T_68222; // @[Switch.scala 41:38:@29382.4]
  assign _T_68225 = select_9 == 6'h22; // @[Switch.scala 41:52:@29384.4]
  assign output_34_9 = io_outValid_9 & _T_68225; // @[Switch.scala 41:38:@29385.4]
  assign _T_68228 = select_10 == 6'h22; // @[Switch.scala 41:52:@29387.4]
  assign output_34_10 = io_outValid_10 & _T_68228; // @[Switch.scala 41:38:@29388.4]
  assign _T_68231 = select_11 == 6'h22; // @[Switch.scala 41:52:@29390.4]
  assign output_34_11 = io_outValid_11 & _T_68231; // @[Switch.scala 41:38:@29391.4]
  assign _T_68234 = select_12 == 6'h22; // @[Switch.scala 41:52:@29393.4]
  assign output_34_12 = io_outValid_12 & _T_68234; // @[Switch.scala 41:38:@29394.4]
  assign _T_68237 = select_13 == 6'h22; // @[Switch.scala 41:52:@29396.4]
  assign output_34_13 = io_outValid_13 & _T_68237; // @[Switch.scala 41:38:@29397.4]
  assign _T_68240 = select_14 == 6'h22; // @[Switch.scala 41:52:@29399.4]
  assign output_34_14 = io_outValid_14 & _T_68240; // @[Switch.scala 41:38:@29400.4]
  assign _T_68243 = select_15 == 6'h22; // @[Switch.scala 41:52:@29402.4]
  assign output_34_15 = io_outValid_15 & _T_68243; // @[Switch.scala 41:38:@29403.4]
  assign _T_68246 = select_16 == 6'h22; // @[Switch.scala 41:52:@29405.4]
  assign output_34_16 = io_outValid_16 & _T_68246; // @[Switch.scala 41:38:@29406.4]
  assign _T_68249 = select_17 == 6'h22; // @[Switch.scala 41:52:@29408.4]
  assign output_34_17 = io_outValid_17 & _T_68249; // @[Switch.scala 41:38:@29409.4]
  assign _T_68252 = select_18 == 6'h22; // @[Switch.scala 41:52:@29411.4]
  assign output_34_18 = io_outValid_18 & _T_68252; // @[Switch.scala 41:38:@29412.4]
  assign _T_68255 = select_19 == 6'h22; // @[Switch.scala 41:52:@29414.4]
  assign output_34_19 = io_outValid_19 & _T_68255; // @[Switch.scala 41:38:@29415.4]
  assign _T_68258 = select_20 == 6'h22; // @[Switch.scala 41:52:@29417.4]
  assign output_34_20 = io_outValid_20 & _T_68258; // @[Switch.scala 41:38:@29418.4]
  assign _T_68261 = select_21 == 6'h22; // @[Switch.scala 41:52:@29420.4]
  assign output_34_21 = io_outValid_21 & _T_68261; // @[Switch.scala 41:38:@29421.4]
  assign _T_68264 = select_22 == 6'h22; // @[Switch.scala 41:52:@29423.4]
  assign output_34_22 = io_outValid_22 & _T_68264; // @[Switch.scala 41:38:@29424.4]
  assign _T_68267 = select_23 == 6'h22; // @[Switch.scala 41:52:@29426.4]
  assign output_34_23 = io_outValid_23 & _T_68267; // @[Switch.scala 41:38:@29427.4]
  assign _T_68270 = select_24 == 6'h22; // @[Switch.scala 41:52:@29429.4]
  assign output_34_24 = io_outValid_24 & _T_68270; // @[Switch.scala 41:38:@29430.4]
  assign _T_68273 = select_25 == 6'h22; // @[Switch.scala 41:52:@29432.4]
  assign output_34_25 = io_outValid_25 & _T_68273; // @[Switch.scala 41:38:@29433.4]
  assign _T_68276 = select_26 == 6'h22; // @[Switch.scala 41:52:@29435.4]
  assign output_34_26 = io_outValid_26 & _T_68276; // @[Switch.scala 41:38:@29436.4]
  assign _T_68279 = select_27 == 6'h22; // @[Switch.scala 41:52:@29438.4]
  assign output_34_27 = io_outValid_27 & _T_68279; // @[Switch.scala 41:38:@29439.4]
  assign _T_68282 = select_28 == 6'h22; // @[Switch.scala 41:52:@29441.4]
  assign output_34_28 = io_outValid_28 & _T_68282; // @[Switch.scala 41:38:@29442.4]
  assign _T_68285 = select_29 == 6'h22; // @[Switch.scala 41:52:@29444.4]
  assign output_34_29 = io_outValid_29 & _T_68285; // @[Switch.scala 41:38:@29445.4]
  assign _T_68288 = select_30 == 6'h22; // @[Switch.scala 41:52:@29447.4]
  assign output_34_30 = io_outValid_30 & _T_68288; // @[Switch.scala 41:38:@29448.4]
  assign _T_68291 = select_31 == 6'h22; // @[Switch.scala 41:52:@29450.4]
  assign output_34_31 = io_outValid_31 & _T_68291; // @[Switch.scala 41:38:@29451.4]
  assign _T_68294 = select_32 == 6'h22; // @[Switch.scala 41:52:@29453.4]
  assign output_34_32 = io_outValid_32 & _T_68294; // @[Switch.scala 41:38:@29454.4]
  assign _T_68297 = select_33 == 6'h22; // @[Switch.scala 41:52:@29456.4]
  assign output_34_33 = io_outValid_33 & _T_68297; // @[Switch.scala 41:38:@29457.4]
  assign _T_68300 = select_34 == 6'h22; // @[Switch.scala 41:52:@29459.4]
  assign output_34_34 = io_outValid_34 & _T_68300; // @[Switch.scala 41:38:@29460.4]
  assign _T_68303 = select_35 == 6'h22; // @[Switch.scala 41:52:@29462.4]
  assign output_34_35 = io_outValid_35 & _T_68303; // @[Switch.scala 41:38:@29463.4]
  assign _T_68306 = select_36 == 6'h22; // @[Switch.scala 41:52:@29465.4]
  assign output_34_36 = io_outValid_36 & _T_68306; // @[Switch.scala 41:38:@29466.4]
  assign _T_68309 = select_37 == 6'h22; // @[Switch.scala 41:52:@29468.4]
  assign output_34_37 = io_outValid_37 & _T_68309; // @[Switch.scala 41:38:@29469.4]
  assign _T_68312 = select_38 == 6'h22; // @[Switch.scala 41:52:@29471.4]
  assign output_34_38 = io_outValid_38 & _T_68312; // @[Switch.scala 41:38:@29472.4]
  assign _T_68315 = select_39 == 6'h22; // @[Switch.scala 41:52:@29474.4]
  assign output_34_39 = io_outValid_39 & _T_68315; // @[Switch.scala 41:38:@29475.4]
  assign _T_68318 = select_40 == 6'h22; // @[Switch.scala 41:52:@29477.4]
  assign output_34_40 = io_outValid_40 & _T_68318; // @[Switch.scala 41:38:@29478.4]
  assign _T_68321 = select_41 == 6'h22; // @[Switch.scala 41:52:@29480.4]
  assign output_34_41 = io_outValid_41 & _T_68321; // @[Switch.scala 41:38:@29481.4]
  assign _T_68324 = select_42 == 6'h22; // @[Switch.scala 41:52:@29483.4]
  assign output_34_42 = io_outValid_42 & _T_68324; // @[Switch.scala 41:38:@29484.4]
  assign _T_68327 = select_43 == 6'h22; // @[Switch.scala 41:52:@29486.4]
  assign output_34_43 = io_outValid_43 & _T_68327; // @[Switch.scala 41:38:@29487.4]
  assign _T_68330 = select_44 == 6'h22; // @[Switch.scala 41:52:@29489.4]
  assign output_34_44 = io_outValid_44 & _T_68330; // @[Switch.scala 41:38:@29490.4]
  assign _T_68333 = select_45 == 6'h22; // @[Switch.scala 41:52:@29492.4]
  assign output_34_45 = io_outValid_45 & _T_68333; // @[Switch.scala 41:38:@29493.4]
  assign _T_68336 = select_46 == 6'h22; // @[Switch.scala 41:52:@29495.4]
  assign output_34_46 = io_outValid_46 & _T_68336; // @[Switch.scala 41:38:@29496.4]
  assign _T_68339 = select_47 == 6'h22; // @[Switch.scala 41:52:@29498.4]
  assign output_34_47 = io_outValid_47 & _T_68339; // @[Switch.scala 41:38:@29499.4]
  assign _T_68342 = select_48 == 6'h22; // @[Switch.scala 41:52:@29501.4]
  assign output_34_48 = io_outValid_48 & _T_68342; // @[Switch.scala 41:38:@29502.4]
  assign _T_68345 = select_49 == 6'h22; // @[Switch.scala 41:52:@29504.4]
  assign output_34_49 = io_outValid_49 & _T_68345; // @[Switch.scala 41:38:@29505.4]
  assign _T_68348 = select_50 == 6'h22; // @[Switch.scala 41:52:@29507.4]
  assign output_34_50 = io_outValid_50 & _T_68348; // @[Switch.scala 41:38:@29508.4]
  assign _T_68351 = select_51 == 6'h22; // @[Switch.scala 41:52:@29510.4]
  assign output_34_51 = io_outValid_51 & _T_68351; // @[Switch.scala 41:38:@29511.4]
  assign _T_68354 = select_52 == 6'h22; // @[Switch.scala 41:52:@29513.4]
  assign output_34_52 = io_outValid_52 & _T_68354; // @[Switch.scala 41:38:@29514.4]
  assign _T_68357 = select_53 == 6'h22; // @[Switch.scala 41:52:@29516.4]
  assign output_34_53 = io_outValid_53 & _T_68357; // @[Switch.scala 41:38:@29517.4]
  assign _T_68360 = select_54 == 6'h22; // @[Switch.scala 41:52:@29519.4]
  assign output_34_54 = io_outValid_54 & _T_68360; // @[Switch.scala 41:38:@29520.4]
  assign _T_68363 = select_55 == 6'h22; // @[Switch.scala 41:52:@29522.4]
  assign output_34_55 = io_outValid_55 & _T_68363; // @[Switch.scala 41:38:@29523.4]
  assign _T_68366 = select_56 == 6'h22; // @[Switch.scala 41:52:@29525.4]
  assign output_34_56 = io_outValid_56 & _T_68366; // @[Switch.scala 41:38:@29526.4]
  assign _T_68369 = select_57 == 6'h22; // @[Switch.scala 41:52:@29528.4]
  assign output_34_57 = io_outValid_57 & _T_68369; // @[Switch.scala 41:38:@29529.4]
  assign _T_68372 = select_58 == 6'h22; // @[Switch.scala 41:52:@29531.4]
  assign output_34_58 = io_outValid_58 & _T_68372; // @[Switch.scala 41:38:@29532.4]
  assign _T_68375 = select_59 == 6'h22; // @[Switch.scala 41:52:@29534.4]
  assign output_34_59 = io_outValid_59 & _T_68375; // @[Switch.scala 41:38:@29535.4]
  assign _T_68378 = select_60 == 6'h22; // @[Switch.scala 41:52:@29537.4]
  assign output_34_60 = io_outValid_60 & _T_68378; // @[Switch.scala 41:38:@29538.4]
  assign _T_68381 = select_61 == 6'h22; // @[Switch.scala 41:52:@29540.4]
  assign output_34_61 = io_outValid_61 & _T_68381; // @[Switch.scala 41:38:@29541.4]
  assign _T_68384 = select_62 == 6'h22; // @[Switch.scala 41:52:@29543.4]
  assign output_34_62 = io_outValid_62 & _T_68384; // @[Switch.scala 41:38:@29544.4]
  assign _T_68387 = select_63 == 6'h22; // @[Switch.scala 41:52:@29546.4]
  assign output_34_63 = io_outValid_63 & _T_68387; // @[Switch.scala 41:38:@29547.4]
  assign _T_68395 = {output_34_7,output_34_6,output_34_5,output_34_4,output_34_3,output_34_2,output_34_1,output_34_0}; // @[Switch.scala 43:31:@29555.4]
  assign _T_68403 = {output_34_15,output_34_14,output_34_13,output_34_12,output_34_11,output_34_10,output_34_9,output_34_8,_T_68395}; // @[Switch.scala 43:31:@29563.4]
  assign _T_68410 = {output_34_23,output_34_22,output_34_21,output_34_20,output_34_19,output_34_18,output_34_17,output_34_16}; // @[Switch.scala 43:31:@29570.4]
  assign _T_68419 = {output_34_31,output_34_30,output_34_29,output_34_28,output_34_27,output_34_26,output_34_25,output_34_24,_T_68410,_T_68403}; // @[Switch.scala 43:31:@29579.4]
  assign _T_68426 = {output_34_39,output_34_38,output_34_37,output_34_36,output_34_35,output_34_34,output_34_33,output_34_32}; // @[Switch.scala 43:31:@29586.4]
  assign _T_68434 = {output_34_47,output_34_46,output_34_45,output_34_44,output_34_43,output_34_42,output_34_41,output_34_40,_T_68426}; // @[Switch.scala 43:31:@29594.4]
  assign _T_68441 = {output_34_55,output_34_54,output_34_53,output_34_52,output_34_51,output_34_50,output_34_49,output_34_48}; // @[Switch.scala 43:31:@29601.4]
  assign _T_68450 = {output_34_63,output_34_62,output_34_61,output_34_60,output_34_59,output_34_58,output_34_57,output_34_56,_T_68441,_T_68434}; // @[Switch.scala 43:31:@29610.4]
  assign _T_68451 = {_T_68450,_T_68419}; // @[Switch.scala 43:31:@29611.4]
  assign _T_68455 = select_0 == 6'h23; // @[Switch.scala 41:52:@29614.4]
  assign output_35_0 = io_outValid_0 & _T_68455; // @[Switch.scala 41:38:@29615.4]
  assign _T_68458 = select_1 == 6'h23; // @[Switch.scala 41:52:@29617.4]
  assign output_35_1 = io_outValid_1 & _T_68458; // @[Switch.scala 41:38:@29618.4]
  assign _T_68461 = select_2 == 6'h23; // @[Switch.scala 41:52:@29620.4]
  assign output_35_2 = io_outValid_2 & _T_68461; // @[Switch.scala 41:38:@29621.4]
  assign _T_68464 = select_3 == 6'h23; // @[Switch.scala 41:52:@29623.4]
  assign output_35_3 = io_outValid_3 & _T_68464; // @[Switch.scala 41:38:@29624.4]
  assign _T_68467 = select_4 == 6'h23; // @[Switch.scala 41:52:@29626.4]
  assign output_35_4 = io_outValid_4 & _T_68467; // @[Switch.scala 41:38:@29627.4]
  assign _T_68470 = select_5 == 6'h23; // @[Switch.scala 41:52:@29629.4]
  assign output_35_5 = io_outValid_5 & _T_68470; // @[Switch.scala 41:38:@29630.4]
  assign _T_68473 = select_6 == 6'h23; // @[Switch.scala 41:52:@29632.4]
  assign output_35_6 = io_outValid_6 & _T_68473; // @[Switch.scala 41:38:@29633.4]
  assign _T_68476 = select_7 == 6'h23; // @[Switch.scala 41:52:@29635.4]
  assign output_35_7 = io_outValid_7 & _T_68476; // @[Switch.scala 41:38:@29636.4]
  assign _T_68479 = select_8 == 6'h23; // @[Switch.scala 41:52:@29638.4]
  assign output_35_8 = io_outValid_8 & _T_68479; // @[Switch.scala 41:38:@29639.4]
  assign _T_68482 = select_9 == 6'h23; // @[Switch.scala 41:52:@29641.4]
  assign output_35_9 = io_outValid_9 & _T_68482; // @[Switch.scala 41:38:@29642.4]
  assign _T_68485 = select_10 == 6'h23; // @[Switch.scala 41:52:@29644.4]
  assign output_35_10 = io_outValid_10 & _T_68485; // @[Switch.scala 41:38:@29645.4]
  assign _T_68488 = select_11 == 6'h23; // @[Switch.scala 41:52:@29647.4]
  assign output_35_11 = io_outValid_11 & _T_68488; // @[Switch.scala 41:38:@29648.4]
  assign _T_68491 = select_12 == 6'h23; // @[Switch.scala 41:52:@29650.4]
  assign output_35_12 = io_outValid_12 & _T_68491; // @[Switch.scala 41:38:@29651.4]
  assign _T_68494 = select_13 == 6'h23; // @[Switch.scala 41:52:@29653.4]
  assign output_35_13 = io_outValid_13 & _T_68494; // @[Switch.scala 41:38:@29654.4]
  assign _T_68497 = select_14 == 6'h23; // @[Switch.scala 41:52:@29656.4]
  assign output_35_14 = io_outValid_14 & _T_68497; // @[Switch.scala 41:38:@29657.4]
  assign _T_68500 = select_15 == 6'h23; // @[Switch.scala 41:52:@29659.4]
  assign output_35_15 = io_outValid_15 & _T_68500; // @[Switch.scala 41:38:@29660.4]
  assign _T_68503 = select_16 == 6'h23; // @[Switch.scala 41:52:@29662.4]
  assign output_35_16 = io_outValid_16 & _T_68503; // @[Switch.scala 41:38:@29663.4]
  assign _T_68506 = select_17 == 6'h23; // @[Switch.scala 41:52:@29665.4]
  assign output_35_17 = io_outValid_17 & _T_68506; // @[Switch.scala 41:38:@29666.4]
  assign _T_68509 = select_18 == 6'h23; // @[Switch.scala 41:52:@29668.4]
  assign output_35_18 = io_outValid_18 & _T_68509; // @[Switch.scala 41:38:@29669.4]
  assign _T_68512 = select_19 == 6'h23; // @[Switch.scala 41:52:@29671.4]
  assign output_35_19 = io_outValid_19 & _T_68512; // @[Switch.scala 41:38:@29672.4]
  assign _T_68515 = select_20 == 6'h23; // @[Switch.scala 41:52:@29674.4]
  assign output_35_20 = io_outValid_20 & _T_68515; // @[Switch.scala 41:38:@29675.4]
  assign _T_68518 = select_21 == 6'h23; // @[Switch.scala 41:52:@29677.4]
  assign output_35_21 = io_outValid_21 & _T_68518; // @[Switch.scala 41:38:@29678.4]
  assign _T_68521 = select_22 == 6'h23; // @[Switch.scala 41:52:@29680.4]
  assign output_35_22 = io_outValid_22 & _T_68521; // @[Switch.scala 41:38:@29681.4]
  assign _T_68524 = select_23 == 6'h23; // @[Switch.scala 41:52:@29683.4]
  assign output_35_23 = io_outValid_23 & _T_68524; // @[Switch.scala 41:38:@29684.4]
  assign _T_68527 = select_24 == 6'h23; // @[Switch.scala 41:52:@29686.4]
  assign output_35_24 = io_outValid_24 & _T_68527; // @[Switch.scala 41:38:@29687.4]
  assign _T_68530 = select_25 == 6'h23; // @[Switch.scala 41:52:@29689.4]
  assign output_35_25 = io_outValid_25 & _T_68530; // @[Switch.scala 41:38:@29690.4]
  assign _T_68533 = select_26 == 6'h23; // @[Switch.scala 41:52:@29692.4]
  assign output_35_26 = io_outValid_26 & _T_68533; // @[Switch.scala 41:38:@29693.4]
  assign _T_68536 = select_27 == 6'h23; // @[Switch.scala 41:52:@29695.4]
  assign output_35_27 = io_outValid_27 & _T_68536; // @[Switch.scala 41:38:@29696.4]
  assign _T_68539 = select_28 == 6'h23; // @[Switch.scala 41:52:@29698.4]
  assign output_35_28 = io_outValid_28 & _T_68539; // @[Switch.scala 41:38:@29699.4]
  assign _T_68542 = select_29 == 6'h23; // @[Switch.scala 41:52:@29701.4]
  assign output_35_29 = io_outValid_29 & _T_68542; // @[Switch.scala 41:38:@29702.4]
  assign _T_68545 = select_30 == 6'h23; // @[Switch.scala 41:52:@29704.4]
  assign output_35_30 = io_outValid_30 & _T_68545; // @[Switch.scala 41:38:@29705.4]
  assign _T_68548 = select_31 == 6'h23; // @[Switch.scala 41:52:@29707.4]
  assign output_35_31 = io_outValid_31 & _T_68548; // @[Switch.scala 41:38:@29708.4]
  assign _T_68551 = select_32 == 6'h23; // @[Switch.scala 41:52:@29710.4]
  assign output_35_32 = io_outValid_32 & _T_68551; // @[Switch.scala 41:38:@29711.4]
  assign _T_68554 = select_33 == 6'h23; // @[Switch.scala 41:52:@29713.4]
  assign output_35_33 = io_outValid_33 & _T_68554; // @[Switch.scala 41:38:@29714.4]
  assign _T_68557 = select_34 == 6'h23; // @[Switch.scala 41:52:@29716.4]
  assign output_35_34 = io_outValid_34 & _T_68557; // @[Switch.scala 41:38:@29717.4]
  assign _T_68560 = select_35 == 6'h23; // @[Switch.scala 41:52:@29719.4]
  assign output_35_35 = io_outValid_35 & _T_68560; // @[Switch.scala 41:38:@29720.4]
  assign _T_68563 = select_36 == 6'h23; // @[Switch.scala 41:52:@29722.4]
  assign output_35_36 = io_outValid_36 & _T_68563; // @[Switch.scala 41:38:@29723.4]
  assign _T_68566 = select_37 == 6'h23; // @[Switch.scala 41:52:@29725.4]
  assign output_35_37 = io_outValid_37 & _T_68566; // @[Switch.scala 41:38:@29726.4]
  assign _T_68569 = select_38 == 6'h23; // @[Switch.scala 41:52:@29728.4]
  assign output_35_38 = io_outValid_38 & _T_68569; // @[Switch.scala 41:38:@29729.4]
  assign _T_68572 = select_39 == 6'h23; // @[Switch.scala 41:52:@29731.4]
  assign output_35_39 = io_outValid_39 & _T_68572; // @[Switch.scala 41:38:@29732.4]
  assign _T_68575 = select_40 == 6'h23; // @[Switch.scala 41:52:@29734.4]
  assign output_35_40 = io_outValid_40 & _T_68575; // @[Switch.scala 41:38:@29735.4]
  assign _T_68578 = select_41 == 6'h23; // @[Switch.scala 41:52:@29737.4]
  assign output_35_41 = io_outValid_41 & _T_68578; // @[Switch.scala 41:38:@29738.4]
  assign _T_68581 = select_42 == 6'h23; // @[Switch.scala 41:52:@29740.4]
  assign output_35_42 = io_outValid_42 & _T_68581; // @[Switch.scala 41:38:@29741.4]
  assign _T_68584 = select_43 == 6'h23; // @[Switch.scala 41:52:@29743.4]
  assign output_35_43 = io_outValid_43 & _T_68584; // @[Switch.scala 41:38:@29744.4]
  assign _T_68587 = select_44 == 6'h23; // @[Switch.scala 41:52:@29746.4]
  assign output_35_44 = io_outValid_44 & _T_68587; // @[Switch.scala 41:38:@29747.4]
  assign _T_68590 = select_45 == 6'h23; // @[Switch.scala 41:52:@29749.4]
  assign output_35_45 = io_outValid_45 & _T_68590; // @[Switch.scala 41:38:@29750.4]
  assign _T_68593 = select_46 == 6'h23; // @[Switch.scala 41:52:@29752.4]
  assign output_35_46 = io_outValid_46 & _T_68593; // @[Switch.scala 41:38:@29753.4]
  assign _T_68596 = select_47 == 6'h23; // @[Switch.scala 41:52:@29755.4]
  assign output_35_47 = io_outValid_47 & _T_68596; // @[Switch.scala 41:38:@29756.4]
  assign _T_68599 = select_48 == 6'h23; // @[Switch.scala 41:52:@29758.4]
  assign output_35_48 = io_outValid_48 & _T_68599; // @[Switch.scala 41:38:@29759.4]
  assign _T_68602 = select_49 == 6'h23; // @[Switch.scala 41:52:@29761.4]
  assign output_35_49 = io_outValid_49 & _T_68602; // @[Switch.scala 41:38:@29762.4]
  assign _T_68605 = select_50 == 6'h23; // @[Switch.scala 41:52:@29764.4]
  assign output_35_50 = io_outValid_50 & _T_68605; // @[Switch.scala 41:38:@29765.4]
  assign _T_68608 = select_51 == 6'h23; // @[Switch.scala 41:52:@29767.4]
  assign output_35_51 = io_outValid_51 & _T_68608; // @[Switch.scala 41:38:@29768.4]
  assign _T_68611 = select_52 == 6'h23; // @[Switch.scala 41:52:@29770.4]
  assign output_35_52 = io_outValid_52 & _T_68611; // @[Switch.scala 41:38:@29771.4]
  assign _T_68614 = select_53 == 6'h23; // @[Switch.scala 41:52:@29773.4]
  assign output_35_53 = io_outValid_53 & _T_68614; // @[Switch.scala 41:38:@29774.4]
  assign _T_68617 = select_54 == 6'h23; // @[Switch.scala 41:52:@29776.4]
  assign output_35_54 = io_outValid_54 & _T_68617; // @[Switch.scala 41:38:@29777.4]
  assign _T_68620 = select_55 == 6'h23; // @[Switch.scala 41:52:@29779.4]
  assign output_35_55 = io_outValid_55 & _T_68620; // @[Switch.scala 41:38:@29780.4]
  assign _T_68623 = select_56 == 6'h23; // @[Switch.scala 41:52:@29782.4]
  assign output_35_56 = io_outValid_56 & _T_68623; // @[Switch.scala 41:38:@29783.4]
  assign _T_68626 = select_57 == 6'h23; // @[Switch.scala 41:52:@29785.4]
  assign output_35_57 = io_outValid_57 & _T_68626; // @[Switch.scala 41:38:@29786.4]
  assign _T_68629 = select_58 == 6'h23; // @[Switch.scala 41:52:@29788.4]
  assign output_35_58 = io_outValid_58 & _T_68629; // @[Switch.scala 41:38:@29789.4]
  assign _T_68632 = select_59 == 6'h23; // @[Switch.scala 41:52:@29791.4]
  assign output_35_59 = io_outValid_59 & _T_68632; // @[Switch.scala 41:38:@29792.4]
  assign _T_68635 = select_60 == 6'h23; // @[Switch.scala 41:52:@29794.4]
  assign output_35_60 = io_outValid_60 & _T_68635; // @[Switch.scala 41:38:@29795.4]
  assign _T_68638 = select_61 == 6'h23; // @[Switch.scala 41:52:@29797.4]
  assign output_35_61 = io_outValid_61 & _T_68638; // @[Switch.scala 41:38:@29798.4]
  assign _T_68641 = select_62 == 6'h23; // @[Switch.scala 41:52:@29800.4]
  assign output_35_62 = io_outValid_62 & _T_68641; // @[Switch.scala 41:38:@29801.4]
  assign _T_68644 = select_63 == 6'h23; // @[Switch.scala 41:52:@29803.4]
  assign output_35_63 = io_outValid_63 & _T_68644; // @[Switch.scala 41:38:@29804.4]
  assign _T_68652 = {output_35_7,output_35_6,output_35_5,output_35_4,output_35_3,output_35_2,output_35_1,output_35_0}; // @[Switch.scala 43:31:@29812.4]
  assign _T_68660 = {output_35_15,output_35_14,output_35_13,output_35_12,output_35_11,output_35_10,output_35_9,output_35_8,_T_68652}; // @[Switch.scala 43:31:@29820.4]
  assign _T_68667 = {output_35_23,output_35_22,output_35_21,output_35_20,output_35_19,output_35_18,output_35_17,output_35_16}; // @[Switch.scala 43:31:@29827.4]
  assign _T_68676 = {output_35_31,output_35_30,output_35_29,output_35_28,output_35_27,output_35_26,output_35_25,output_35_24,_T_68667,_T_68660}; // @[Switch.scala 43:31:@29836.4]
  assign _T_68683 = {output_35_39,output_35_38,output_35_37,output_35_36,output_35_35,output_35_34,output_35_33,output_35_32}; // @[Switch.scala 43:31:@29843.4]
  assign _T_68691 = {output_35_47,output_35_46,output_35_45,output_35_44,output_35_43,output_35_42,output_35_41,output_35_40,_T_68683}; // @[Switch.scala 43:31:@29851.4]
  assign _T_68698 = {output_35_55,output_35_54,output_35_53,output_35_52,output_35_51,output_35_50,output_35_49,output_35_48}; // @[Switch.scala 43:31:@29858.4]
  assign _T_68707 = {output_35_63,output_35_62,output_35_61,output_35_60,output_35_59,output_35_58,output_35_57,output_35_56,_T_68698,_T_68691}; // @[Switch.scala 43:31:@29867.4]
  assign _T_68708 = {_T_68707,_T_68676}; // @[Switch.scala 43:31:@29868.4]
  assign _T_68712 = select_0 == 6'h24; // @[Switch.scala 41:52:@29871.4]
  assign output_36_0 = io_outValid_0 & _T_68712; // @[Switch.scala 41:38:@29872.4]
  assign _T_68715 = select_1 == 6'h24; // @[Switch.scala 41:52:@29874.4]
  assign output_36_1 = io_outValid_1 & _T_68715; // @[Switch.scala 41:38:@29875.4]
  assign _T_68718 = select_2 == 6'h24; // @[Switch.scala 41:52:@29877.4]
  assign output_36_2 = io_outValid_2 & _T_68718; // @[Switch.scala 41:38:@29878.4]
  assign _T_68721 = select_3 == 6'h24; // @[Switch.scala 41:52:@29880.4]
  assign output_36_3 = io_outValid_3 & _T_68721; // @[Switch.scala 41:38:@29881.4]
  assign _T_68724 = select_4 == 6'h24; // @[Switch.scala 41:52:@29883.4]
  assign output_36_4 = io_outValid_4 & _T_68724; // @[Switch.scala 41:38:@29884.4]
  assign _T_68727 = select_5 == 6'h24; // @[Switch.scala 41:52:@29886.4]
  assign output_36_5 = io_outValid_5 & _T_68727; // @[Switch.scala 41:38:@29887.4]
  assign _T_68730 = select_6 == 6'h24; // @[Switch.scala 41:52:@29889.4]
  assign output_36_6 = io_outValid_6 & _T_68730; // @[Switch.scala 41:38:@29890.4]
  assign _T_68733 = select_7 == 6'h24; // @[Switch.scala 41:52:@29892.4]
  assign output_36_7 = io_outValid_7 & _T_68733; // @[Switch.scala 41:38:@29893.4]
  assign _T_68736 = select_8 == 6'h24; // @[Switch.scala 41:52:@29895.4]
  assign output_36_8 = io_outValid_8 & _T_68736; // @[Switch.scala 41:38:@29896.4]
  assign _T_68739 = select_9 == 6'h24; // @[Switch.scala 41:52:@29898.4]
  assign output_36_9 = io_outValid_9 & _T_68739; // @[Switch.scala 41:38:@29899.4]
  assign _T_68742 = select_10 == 6'h24; // @[Switch.scala 41:52:@29901.4]
  assign output_36_10 = io_outValid_10 & _T_68742; // @[Switch.scala 41:38:@29902.4]
  assign _T_68745 = select_11 == 6'h24; // @[Switch.scala 41:52:@29904.4]
  assign output_36_11 = io_outValid_11 & _T_68745; // @[Switch.scala 41:38:@29905.4]
  assign _T_68748 = select_12 == 6'h24; // @[Switch.scala 41:52:@29907.4]
  assign output_36_12 = io_outValid_12 & _T_68748; // @[Switch.scala 41:38:@29908.4]
  assign _T_68751 = select_13 == 6'h24; // @[Switch.scala 41:52:@29910.4]
  assign output_36_13 = io_outValid_13 & _T_68751; // @[Switch.scala 41:38:@29911.4]
  assign _T_68754 = select_14 == 6'h24; // @[Switch.scala 41:52:@29913.4]
  assign output_36_14 = io_outValid_14 & _T_68754; // @[Switch.scala 41:38:@29914.4]
  assign _T_68757 = select_15 == 6'h24; // @[Switch.scala 41:52:@29916.4]
  assign output_36_15 = io_outValid_15 & _T_68757; // @[Switch.scala 41:38:@29917.4]
  assign _T_68760 = select_16 == 6'h24; // @[Switch.scala 41:52:@29919.4]
  assign output_36_16 = io_outValid_16 & _T_68760; // @[Switch.scala 41:38:@29920.4]
  assign _T_68763 = select_17 == 6'h24; // @[Switch.scala 41:52:@29922.4]
  assign output_36_17 = io_outValid_17 & _T_68763; // @[Switch.scala 41:38:@29923.4]
  assign _T_68766 = select_18 == 6'h24; // @[Switch.scala 41:52:@29925.4]
  assign output_36_18 = io_outValid_18 & _T_68766; // @[Switch.scala 41:38:@29926.4]
  assign _T_68769 = select_19 == 6'h24; // @[Switch.scala 41:52:@29928.4]
  assign output_36_19 = io_outValid_19 & _T_68769; // @[Switch.scala 41:38:@29929.4]
  assign _T_68772 = select_20 == 6'h24; // @[Switch.scala 41:52:@29931.4]
  assign output_36_20 = io_outValid_20 & _T_68772; // @[Switch.scala 41:38:@29932.4]
  assign _T_68775 = select_21 == 6'h24; // @[Switch.scala 41:52:@29934.4]
  assign output_36_21 = io_outValid_21 & _T_68775; // @[Switch.scala 41:38:@29935.4]
  assign _T_68778 = select_22 == 6'h24; // @[Switch.scala 41:52:@29937.4]
  assign output_36_22 = io_outValid_22 & _T_68778; // @[Switch.scala 41:38:@29938.4]
  assign _T_68781 = select_23 == 6'h24; // @[Switch.scala 41:52:@29940.4]
  assign output_36_23 = io_outValid_23 & _T_68781; // @[Switch.scala 41:38:@29941.4]
  assign _T_68784 = select_24 == 6'h24; // @[Switch.scala 41:52:@29943.4]
  assign output_36_24 = io_outValid_24 & _T_68784; // @[Switch.scala 41:38:@29944.4]
  assign _T_68787 = select_25 == 6'h24; // @[Switch.scala 41:52:@29946.4]
  assign output_36_25 = io_outValid_25 & _T_68787; // @[Switch.scala 41:38:@29947.4]
  assign _T_68790 = select_26 == 6'h24; // @[Switch.scala 41:52:@29949.4]
  assign output_36_26 = io_outValid_26 & _T_68790; // @[Switch.scala 41:38:@29950.4]
  assign _T_68793 = select_27 == 6'h24; // @[Switch.scala 41:52:@29952.4]
  assign output_36_27 = io_outValid_27 & _T_68793; // @[Switch.scala 41:38:@29953.4]
  assign _T_68796 = select_28 == 6'h24; // @[Switch.scala 41:52:@29955.4]
  assign output_36_28 = io_outValid_28 & _T_68796; // @[Switch.scala 41:38:@29956.4]
  assign _T_68799 = select_29 == 6'h24; // @[Switch.scala 41:52:@29958.4]
  assign output_36_29 = io_outValid_29 & _T_68799; // @[Switch.scala 41:38:@29959.4]
  assign _T_68802 = select_30 == 6'h24; // @[Switch.scala 41:52:@29961.4]
  assign output_36_30 = io_outValid_30 & _T_68802; // @[Switch.scala 41:38:@29962.4]
  assign _T_68805 = select_31 == 6'h24; // @[Switch.scala 41:52:@29964.4]
  assign output_36_31 = io_outValid_31 & _T_68805; // @[Switch.scala 41:38:@29965.4]
  assign _T_68808 = select_32 == 6'h24; // @[Switch.scala 41:52:@29967.4]
  assign output_36_32 = io_outValid_32 & _T_68808; // @[Switch.scala 41:38:@29968.4]
  assign _T_68811 = select_33 == 6'h24; // @[Switch.scala 41:52:@29970.4]
  assign output_36_33 = io_outValid_33 & _T_68811; // @[Switch.scala 41:38:@29971.4]
  assign _T_68814 = select_34 == 6'h24; // @[Switch.scala 41:52:@29973.4]
  assign output_36_34 = io_outValid_34 & _T_68814; // @[Switch.scala 41:38:@29974.4]
  assign _T_68817 = select_35 == 6'h24; // @[Switch.scala 41:52:@29976.4]
  assign output_36_35 = io_outValid_35 & _T_68817; // @[Switch.scala 41:38:@29977.4]
  assign _T_68820 = select_36 == 6'h24; // @[Switch.scala 41:52:@29979.4]
  assign output_36_36 = io_outValid_36 & _T_68820; // @[Switch.scala 41:38:@29980.4]
  assign _T_68823 = select_37 == 6'h24; // @[Switch.scala 41:52:@29982.4]
  assign output_36_37 = io_outValid_37 & _T_68823; // @[Switch.scala 41:38:@29983.4]
  assign _T_68826 = select_38 == 6'h24; // @[Switch.scala 41:52:@29985.4]
  assign output_36_38 = io_outValid_38 & _T_68826; // @[Switch.scala 41:38:@29986.4]
  assign _T_68829 = select_39 == 6'h24; // @[Switch.scala 41:52:@29988.4]
  assign output_36_39 = io_outValid_39 & _T_68829; // @[Switch.scala 41:38:@29989.4]
  assign _T_68832 = select_40 == 6'h24; // @[Switch.scala 41:52:@29991.4]
  assign output_36_40 = io_outValid_40 & _T_68832; // @[Switch.scala 41:38:@29992.4]
  assign _T_68835 = select_41 == 6'h24; // @[Switch.scala 41:52:@29994.4]
  assign output_36_41 = io_outValid_41 & _T_68835; // @[Switch.scala 41:38:@29995.4]
  assign _T_68838 = select_42 == 6'h24; // @[Switch.scala 41:52:@29997.4]
  assign output_36_42 = io_outValid_42 & _T_68838; // @[Switch.scala 41:38:@29998.4]
  assign _T_68841 = select_43 == 6'h24; // @[Switch.scala 41:52:@30000.4]
  assign output_36_43 = io_outValid_43 & _T_68841; // @[Switch.scala 41:38:@30001.4]
  assign _T_68844 = select_44 == 6'h24; // @[Switch.scala 41:52:@30003.4]
  assign output_36_44 = io_outValid_44 & _T_68844; // @[Switch.scala 41:38:@30004.4]
  assign _T_68847 = select_45 == 6'h24; // @[Switch.scala 41:52:@30006.4]
  assign output_36_45 = io_outValid_45 & _T_68847; // @[Switch.scala 41:38:@30007.4]
  assign _T_68850 = select_46 == 6'h24; // @[Switch.scala 41:52:@30009.4]
  assign output_36_46 = io_outValid_46 & _T_68850; // @[Switch.scala 41:38:@30010.4]
  assign _T_68853 = select_47 == 6'h24; // @[Switch.scala 41:52:@30012.4]
  assign output_36_47 = io_outValid_47 & _T_68853; // @[Switch.scala 41:38:@30013.4]
  assign _T_68856 = select_48 == 6'h24; // @[Switch.scala 41:52:@30015.4]
  assign output_36_48 = io_outValid_48 & _T_68856; // @[Switch.scala 41:38:@30016.4]
  assign _T_68859 = select_49 == 6'h24; // @[Switch.scala 41:52:@30018.4]
  assign output_36_49 = io_outValid_49 & _T_68859; // @[Switch.scala 41:38:@30019.4]
  assign _T_68862 = select_50 == 6'h24; // @[Switch.scala 41:52:@30021.4]
  assign output_36_50 = io_outValid_50 & _T_68862; // @[Switch.scala 41:38:@30022.4]
  assign _T_68865 = select_51 == 6'h24; // @[Switch.scala 41:52:@30024.4]
  assign output_36_51 = io_outValid_51 & _T_68865; // @[Switch.scala 41:38:@30025.4]
  assign _T_68868 = select_52 == 6'h24; // @[Switch.scala 41:52:@30027.4]
  assign output_36_52 = io_outValid_52 & _T_68868; // @[Switch.scala 41:38:@30028.4]
  assign _T_68871 = select_53 == 6'h24; // @[Switch.scala 41:52:@30030.4]
  assign output_36_53 = io_outValid_53 & _T_68871; // @[Switch.scala 41:38:@30031.4]
  assign _T_68874 = select_54 == 6'h24; // @[Switch.scala 41:52:@30033.4]
  assign output_36_54 = io_outValid_54 & _T_68874; // @[Switch.scala 41:38:@30034.4]
  assign _T_68877 = select_55 == 6'h24; // @[Switch.scala 41:52:@30036.4]
  assign output_36_55 = io_outValid_55 & _T_68877; // @[Switch.scala 41:38:@30037.4]
  assign _T_68880 = select_56 == 6'h24; // @[Switch.scala 41:52:@30039.4]
  assign output_36_56 = io_outValid_56 & _T_68880; // @[Switch.scala 41:38:@30040.4]
  assign _T_68883 = select_57 == 6'h24; // @[Switch.scala 41:52:@30042.4]
  assign output_36_57 = io_outValid_57 & _T_68883; // @[Switch.scala 41:38:@30043.4]
  assign _T_68886 = select_58 == 6'h24; // @[Switch.scala 41:52:@30045.4]
  assign output_36_58 = io_outValid_58 & _T_68886; // @[Switch.scala 41:38:@30046.4]
  assign _T_68889 = select_59 == 6'h24; // @[Switch.scala 41:52:@30048.4]
  assign output_36_59 = io_outValid_59 & _T_68889; // @[Switch.scala 41:38:@30049.4]
  assign _T_68892 = select_60 == 6'h24; // @[Switch.scala 41:52:@30051.4]
  assign output_36_60 = io_outValid_60 & _T_68892; // @[Switch.scala 41:38:@30052.4]
  assign _T_68895 = select_61 == 6'h24; // @[Switch.scala 41:52:@30054.4]
  assign output_36_61 = io_outValid_61 & _T_68895; // @[Switch.scala 41:38:@30055.4]
  assign _T_68898 = select_62 == 6'h24; // @[Switch.scala 41:52:@30057.4]
  assign output_36_62 = io_outValid_62 & _T_68898; // @[Switch.scala 41:38:@30058.4]
  assign _T_68901 = select_63 == 6'h24; // @[Switch.scala 41:52:@30060.4]
  assign output_36_63 = io_outValid_63 & _T_68901; // @[Switch.scala 41:38:@30061.4]
  assign _T_68909 = {output_36_7,output_36_6,output_36_5,output_36_4,output_36_3,output_36_2,output_36_1,output_36_0}; // @[Switch.scala 43:31:@30069.4]
  assign _T_68917 = {output_36_15,output_36_14,output_36_13,output_36_12,output_36_11,output_36_10,output_36_9,output_36_8,_T_68909}; // @[Switch.scala 43:31:@30077.4]
  assign _T_68924 = {output_36_23,output_36_22,output_36_21,output_36_20,output_36_19,output_36_18,output_36_17,output_36_16}; // @[Switch.scala 43:31:@30084.4]
  assign _T_68933 = {output_36_31,output_36_30,output_36_29,output_36_28,output_36_27,output_36_26,output_36_25,output_36_24,_T_68924,_T_68917}; // @[Switch.scala 43:31:@30093.4]
  assign _T_68940 = {output_36_39,output_36_38,output_36_37,output_36_36,output_36_35,output_36_34,output_36_33,output_36_32}; // @[Switch.scala 43:31:@30100.4]
  assign _T_68948 = {output_36_47,output_36_46,output_36_45,output_36_44,output_36_43,output_36_42,output_36_41,output_36_40,_T_68940}; // @[Switch.scala 43:31:@30108.4]
  assign _T_68955 = {output_36_55,output_36_54,output_36_53,output_36_52,output_36_51,output_36_50,output_36_49,output_36_48}; // @[Switch.scala 43:31:@30115.4]
  assign _T_68964 = {output_36_63,output_36_62,output_36_61,output_36_60,output_36_59,output_36_58,output_36_57,output_36_56,_T_68955,_T_68948}; // @[Switch.scala 43:31:@30124.4]
  assign _T_68965 = {_T_68964,_T_68933}; // @[Switch.scala 43:31:@30125.4]
  assign _T_68969 = select_0 == 6'h25; // @[Switch.scala 41:52:@30128.4]
  assign output_37_0 = io_outValid_0 & _T_68969; // @[Switch.scala 41:38:@30129.4]
  assign _T_68972 = select_1 == 6'h25; // @[Switch.scala 41:52:@30131.4]
  assign output_37_1 = io_outValid_1 & _T_68972; // @[Switch.scala 41:38:@30132.4]
  assign _T_68975 = select_2 == 6'h25; // @[Switch.scala 41:52:@30134.4]
  assign output_37_2 = io_outValid_2 & _T_68975; // @[Switch.scala 41:38:@30135.4]
  assign _T_68978 = select_3 == 6'h25; // @[Switch.scala 41:52:@30137.4]
  assign output_37_3 = io_outValid_3 & _T_68978; // @[Switch.scala 41:38:@30138.4]
  assign _T_68981 = select_4 == 6'h25; // @[Switch.scala 41:52:@30140.4]
  assign output_37_4 = io_outValid_4 & _T_68981; // @[Switch.scala 41:38:@30141.4]
  assign _T_68984 = select_5 == 6'h25; // @[Switch.scala 41:52:@30143.4]
  assign output_37_5 = io_outValid_5 & _T_68984; // @[Switch.scala 41:38:@30144.4]
  assign _T_68987 = select_6 == 6'h25; // @[Switch.scala 41:52:@30146.4]
  assign output_37_6 = io_outValid_6 & _T_68987; // @[Switch.scala 41:38:@30147.4]
  assign _T_68990 = select_7 == 6'h25; // @[Switch.scala 41:52:@30149.4]
  assign output_37_7 = io_outValid_7 & _T_68990; // @[Switch.scala 41:38:@30150.4]
  assign _T_68993 = select_8 == 6'h25; // @[Switch.scala 41:52:@30152.4]
  assign output_37_8 = io_outValid_8 & _T_68993; // @[Switch.scala 41:38:@30153.4]
  assign _T_68996 = select_9 == 6'h25; // @[Switch.scala 41:52:@30155.4]
  assign output_37_9 = io_outValid_9 & _T_68996; // @[Switch.scala 41:38:@30156.4]
  assign _T_68999 = select_10 == 6'h25; // @[Switch.scala 41:52:@30158.4]
  assign output_37_10 = io_outValid_10 & _T_68999; // @[Switch.scala 41:38:@30159.4]
  assign _T_69002 = select_11 == 6'h25; // @[Switch.scala 41:52:@30161.4]
  assign output_37_11 = io_outValid_11 & _T_69002; // @[Switch.scala 41:38:@30162.4]
  assign _T_69005 = select_12 == 6'h25; // @[Switch.scala 41:52:@30164.4]
  assign output_37_12 = io_outValid_12 & _T_69005; // @[Switch.scala 41:38:@30165.4]
  assign _T_69008 = select_13 == 6'h25; // @[Switch.scala 41:52:@30167.4]
  assign output_37_13 = io_outValid_13 & _T_69008; // @[Switch.scala 41:38:@30168.4]
  assign _T_69011 = select_14 == 6'h25; // @[Switch.scala 41:52:@30170.4]
  assign output_37_14 = io_outValid_14 & _T_69011; // @[Switch.scala 41:38:@30171.4]
  assign _T_69014 = select_15 == 6'h25; // @[Switch.scala 41:52:@30173.4]
  assign output_37_15 = io_outValid_15 & _T_69014; // @[Switch.scala 41:38:@30174.4]
  assign _T_69017 = select_16 == 6'h25; // @[Switch.scala 41:52:@30176.4]
  assign output_37_16 = io_outValid_16 & _T_69017; // @[Switch.scala 41:38:@30177.4]
  assign _T_69020 = select_17 == 6'h25; // @[Switch.scala 41:52:@30179.4]
  assign output_37_17 = io_outValid_17 & _T_69020; // @[Switch.scala 41:38:@30180.4]
  assign _T_69023 = select_18 == 6'h25; // @[Switch.scala 41:52:@30182.4]
  assign output_37_18 = io_outValid_18 & _T_69023; // @[Switch.scala 41:38:@30183.4]
  assign _T_69026 = select_19 == 6'h25; // @[Switch.scala 41:52:@30185.4]
  assign output_37_19 = io_outValid_19 & _T_69026; // @[Switch.scala 41:38:@30186.4]
  assign _T_69029 = select_20 == 6'h25; // @[Switch.scala 41:52:@30188.4]
  assign output_37_20 = io_outValid_20 & _T_69029; // @[Switch.scala 41:38:@30189.4]
  assign _T_69032 = select_21 == 6'h25; // @[Switch.scala 41:52:@30191.4]
  assign output_37_21 = io_outValid_21 & _T_69032; // @[Switch.scala 41:38:@30192.4]
  assign _T_69035 = select_22 == 6'h25; // @[Switch.scala 41:52:@30194.4]
  assign output_37_22 = io_outValid_22 & _T_69035; // @[Switch.scala 41:38:@30195.4]
  assign _T_69038 = select_23 == 6'h25; // @[Switch.scala 41:52:@30197.4]
  assign output_37_23 = io_outValid_23 & _T_69038; // @[Switch.scala 41:38:@30198.4]
  assign _T_69041 = select_24 == 6'h25; // @[Switch.scala 41:52:@30200.4]
  assign output_37_24 = io_outValid_24 & _T_69041; // @[Switch.scala 41:38:@30201.4]
  assign _T_69044 = select_25 == 6'h25; // @[Switch.scala 41:52:@30203.4]
  assign output_37_25 = io_outValid_25 & _T_69044; // @[Switch.scala 41:38:@30204.4]
  assign _T_69047 = select_26 == 6'h25; // @[Switch.scala 41:52:@30206.4]
  assign output_37_26 = io_outValid_26 & _T_69047; // @[Switch.scala 41:38:@30207.4]
  assign _T_69050 = select_27 == 6'h25; // @[Switch.scala 41:52:@30209.4]
  assign output_37_27 = io_outValid_27 & _T_69050; // @[Switch.scala 41:38:@30210.4]
  assign _T_69053 = select_28 == 6'h25; // @[Switch.scala 41:52:@30212.4]
  assign output_37_28 = io_outValid_28 & _T_69053; // @[Switch.scala 41:38:@30213.4]
  assign _T_69056 = select_29 == 6'h25; // @[Switch.scala 41:52:@30215.4]
  assign output_37_29 = io_outValid_29 & _T_69056; // @[Switch.scala 41:38:@30216.4]
  assign _T_69059 = select_30 == 6'h25; // @[Switch.scala 41:52:@30218.4]
  assign output_37_30 = io_outValid_30 & _T_69059; // @[Switch.scala 41:38:@30219.4]
  assign _T_69062 = select_31 == 6'h25; // @[Switch.scala 41:52:@30221.4]
  assign output_37_31 = io_outValid_31 & _T_69062; // @[Switch.scala 41:38:@30222.4]
  assign _T_69065 = select_32 == 6'h25; // @[Switch.scala 41:52:@30224.4]
  assign output_37_32 = io_outValid_32 & _T_69065; // @[Switch.scala 41:38:@30225.4]
  assign _T_69068 = select_33 == 6'h25; // @[Switch.scala 41:52:@30227.4]
  assign output_37_33 = io_outValid_33 & _T_69068; // @[Switch.scala 41:38:@30228.4]
  assign _T_69071 = select_34 == 6'h25; // @[Switch.scala 41:52:@30230.4]
  assign output_37_34 = io_outValid_34 & _T_69071; // @[Switch.scala 41:38:@30231.4]
  assign _T_69074 = select_35 == 6'h25; // @[Switch.scala 41:52:@30233.4]
  assign output_37_35 = io_outValid_35 & _T_69074; // @[Switch.scala 41:38:@30234.4]
  assign _T_69077 = select_36 == 6'h25; // @[Switch.scala 41:52:@30236.4]
  assign output_37_36 = io_outValid_36 & _T_69077; // @[Switch.scala 41:38:@30237.4]
  assign _T_69080 = select_37 == 6'h25; // @[Switch.scala 41:52:@30239.4]
  assign output_37_37 = io_outValid_37 & _T_69080; // @[Switch.scala 41:38:@30240.4]
  assign _T_69083 = select_38 == 6'h25; // @[Switch.scala 41:52:@30242.4]
  assign output_37_38 = io_outValid_38 & _T_69083; // @[Switch.scala 41:38:@30243.4]
  assign _T_69086 = select_39 == 6'h25; // @[Switch.scala 41:52:@30245.4]
  assign output_37_39 = io_outValid_39 & _T_69086; // @[Switch.scala 41:38:@30246.4]
  assign _T_69089 = select_40 == 6'h25; // @[Switch.scala 41:52:@30248.4]
  assign output_37_40 = io_outValid_40 & _T_69089; // @[Switch.scala 41:38:@30249.4]
  assign _T_69092 = select_41 == 6'h25; // @[Switch.scala 41:52:@30251.4]
  assign output_37_41 = io_outValid_41 & _T_69092; // @[Switch.scala 41:38:@30252.4]
  assign _T_69095 = select_42 == 6'h25; // @[Switch.scala 41:52:@30254.4]
  assign output_37_42 = io_outValid_42 & _T_69095; // @[Switch.scala 41:38:@30255.4]
  assign _T_69098 = select_43 == 6'h25; // @[Switch.scala 41:52:@30257.4]
  assign output_37_43 = io_outValid_43 & _T_69098; // @[Switch.scala 41:38:@30258.4]
  assign _T_69101 = select_44 == 6'h25; // @[Switch.scala 41:52:@30260.4]
  assign output_37_44 = io_outValid_44 & _T_69101; // @[Switch.scala 41:38:@30261.4]
  assign _T_69104 = select_45 == 6'h25; // @[Switch.scala 41:52:@30263.4]
  assign output_37_45 = io_outValid_45 & _T_69104; // @[Switch.scala 41:38:@30264.4]
  assign _T_69107 = select_46 == 6'h25; // @[Switch.scala 41:52:@30266.4]
  assign output_37_46 = io_outValid_46 & _T_69107; // @[Switch.scala 41:38:@30267.4]
  assign _T_69110 = select_47 == 6'h25; // @[Switch.scala 41:52:@30269.4]
  assign output_37_47 = io_outValid_47 & _T_69110; // @[Switch.scala 41:38:@30270.4]
  assign _T_69113 = select_48 == 6'h25; // @[Switch.scala 41:52:@30272.4]
  assign output_37_48 = io_outValid_48 & _T_69113; // @[Switch.scala 41:38:@30273.4]
  assign _T_69116 = select_49 == 6'h25; // @[Switch.scala 41:52:@30275.4]
  assign output_37_49 = io_outValid_49 & _T_69116; // @[Switch.scala 41:38:@30276.4]
  assign _T_69119 = select_50 == 6'h25; // @[Switch.scala 41:52:@30278.4]
  assign output_37_50 = io_outValid_50 & _T_69119; // @[Switch.scala 41:38:@30279.4]
  assign _T_69122 = select_51 == 6'h25; // @[Switch.scala 41:52:@30281.4]
  assign output_37_51 = io_outValid_51 & _T_69122; // @[Switch.scala 41:38:@30282.4]
  assign _T_69125 = select_52 == 6'h25; // @[Switch.scala 41:52:@30284.4]
  assign output_37_52 = io_outValid_52 & _T_69125; // @[Switch.scala 41:38:@30285.4]
  assign _T_69128 = select_53 == 6'h25; // @[Switch.scala 41:52:@30287.4]
  assign output_37_53 = io_outValid_53 & _T_69128; // @[Switch.scala 41:38:@30288.4]
  assign _T_69131 = select_54 == 6'h25; // @[Switch.scala 41:52:@30290.4]
  assign output_37_54 = io_outValid_54 & _T_69131; // @[Switch.scala 41:38:@30291.4]
  assign _T_69134 = select_55 == 6'h25; // @[Switch.scala 41:52:@30293.4]
  assign output_37_55 = io_outValid_55 & _T_69134; // @[Switch.scala 41:38:@30294.4]
  assign _T_69137 = select_56 == 6'h25; // @[Switch.scala 41:52:@30296.4]
  assign output_37_56 = io_outValid_56 & _T_69137; // @[Switch.scala 41:38:@30297.4]
  assign _T_69140 = select_57 == 6'h25; // @[Switch.scala 41:52:@30299.4]
  assign output_37_57 = io_outValid_57 & _T_69140; // @[Switch.scala 41:38:@30300.4]
  assign _T_69143 = select_58 == 6'h25; // @[Switch.scala 41:52:@30302.4]
  assign output_37_58 = io_outValid_58 & _T_69143; // @[Switch.scala 41:38:@30303.4]
  assign _T_69146 = select_59 == 6'h25; // @[Switch.scala 41:52:@30305.4]
  assign output_37_59 = io_outValid_59 & _T_69146; // @[Switch.scala 41:38:@30306.4]
  assign _T_69149 = select_60 == 6'h25; // @[Switch.scala 41:52:@30308.4]
  assign output_37_60 = io_outValid_60 & _T_69149; // @[Switch.scala 41:38:@30309.4]
  assign _T_69152 = select_61 == 6'h25; // @[Switch.scala 41:52:@30311.4]
  assign output_37_61 = io_outValid_61 & _T_69152; // @[Switch.scala 41:38:@30312.4]
  assign _T_69155 = select_62 == 6'h25; // @[Switch.scala 41:52:@30314.4]
  assign output_37_62 = io_outValid_62 & _T_69155; // @[Switch.scala 41:38:@30315.4]
  assign _T_69158 = select_63 == 6'h25; // @[Switch.scala 41:52:@30317.4]
  assign output_37_63 = io_outValid_63 & _T_69158; // @[Switch.scala 41:38:@30318.4]
  assign _T_69166 = {output_37_7,output_37_6,output_37_5,output_37_4,output_37_3,output_37_2,output_37_1,output_37_0}; // @[Switch.scala 43:31:@30326.4]
  assign _T_69174 = {output_37_15,output_37_14,output_37_13,output_37_12,output_37_11,output_37_10,output_37_9,output_37_8,_T_69166}; // @[Switch.scala 43:31:@30334.4]
  assign _T_69181 = {output_37_23,output_37_22,output_37_21,output_37_20,output_37_19,output_37_18,output_37_17,output_37_16}; // @[Switch.scala 43:31:@30341.4]
  assign _T_69190 = {output_37_31,output_37_30,output_37_29,output_37_28,output_37_27,output_37_26,output_37_25,output_37_24,_T_69181,_T_69174}; // @[Switch.scala 43:31:@30350.4]
  assign _T_69197 = {output_37_39,output_37_38,output_37_37,output_37_36,output_37_35,output_37_34,output_37_33,output_37_32}; // @[Switch.scala 43:31:@30357.4]
  assign _T_69205 = {output_37_47,output_37_46,output_37_45,output_37_44,output_37_43,output_37_42,output_37_41,output_37_40,_T_69197}; // @[Switch.scala 43:31:@30365.4]
  assign _T_69212 = {output_37_55,output_37_54,output_37_53,output_37_52,output_37_51,output_37_50,output_37_49,output_37_48}; // @[Switch.scala 43:31:@30372.4]
  assign _T_69221 = {output_37_63,output_37_62,output_37_61,output_37_60,output_37_59,output_37_58,output_37_57,output_37_56,_T_69212,_T_69205}; // @[Switch.scala 43:31:@30381.4]
  assign _T_69222 = {_T_69221,_T_69190}; // @[Switch.scala 43:31:@30382.4]
  assign _T_69226 = select_0 == 6'h26; // @[Switch.scala 41:52:@30385.4]
  assign output_38_0 = io_outValid_0 & _T_69226; // @[Switch.scala 41:38:@30386.4]
  assign _T_69229 = select_1 == 6'h26; // @[Switch.scala 41:52:@30388.4]
  assign output_38_1 = io_outValid_1 & _T_69229; // @[Switch.scala 41:38:@30389.4]
  assign _T_69232 = select_2 == 6'h26; // @[Switch.scala 41:52:@30391.4]
  assign output_38_2 = io_outValid_2 & _T_69232; // @[Switch.scala 41:38:@30392.4]
  assign _T_69235 = select_3 == 6'h26; // @[Switch.scala 41:52:@30394.4]
  assign output_38_3 = io_outValid_3 & _T_69235; // @[Switch.scala 41:38:@30395.4]
  assign _T_69238 = select_4 == 6'h26; // @[Switch.scala 41:52:@30397.4]
  assign output_38_4 = io_outValid_4 & _T_69238; // @[Switch.scala 41:38:@30398.4]
  assign _T_69241 = select_5 == 6'h26; // @[Switch.scala 41:52:@30400.4]
  assign output_38_5 = io_outValid_5 & _T_69241; // @[Switch.scala 41:38:@30401.4]
  assign _T_69244 = select_6 == 6'h26; // @[Switch.scala 41:52:@30403.4]
  assign output_38_6 = io_outValid_6 & _T_69244; // @[Switch.scala 41:38:@30404.4]
  assign _T_69247 = select_7 == 6'h26; // @[Switch.scala 41:52:@30406.4]
  assign output_38_7 = io_outValid_7 & _T_69247; // @[Switch.scala 41:38:@30407.4]
  assign _T_69250 = select_8 == 6'h26; // @[Switch.scala 41:52:@30409.4]
  assign output_38_8 = io_outValid_8 & _T_69250; // @[Switch.scala 41:38:@30410.4]
  assign _T_69253 = select_9 == 6'h26; // @[Switch.scala 41:52:@30412.4]
  assign output_38_9 = io_outValid_9 & _T_69253; // @[Switch.scala 41:38:@30413.4]
  assign _T_69256 = select_10 == 6'h26; // @[Switch.scala 41:52:@30415.4]
  assign output_38_10 = io_outValid_10 & _T_69256; // @[Switch.scala 41:38:@30416.4]
  assign _T_69259 = select_11 == 6'h26; // @[Switch.scala 41:52:@30418.4]
  assign output_38_11 = io_outValid_11 & _T_69259; // @[Switch.scala 41:38:@30419.4]
  assign _T_69262 = select_12 == 6'h26; // @[Switch.scala 41:52:@30421.4]
  assign output_38_12 = io_outValid_12 & _T_69262; // @[Switch.scala 41:38:@30422.4]
  assign _T_69265 = select_13 == 6'h26; // @[Switch.scala 41:52:@30424.4]
  assign output_38_13 = io_outValid_13 & _T_69265; // @[Switch.scala 41:38:@30425.4]
  assign _T_69268 = select_14 == 6'h26; // @[Switch.scala 41:52:@30427.4]
  assign output_38_14 = io_outValid_14 & _T_69268; // @[Switch.scala 41:38:@30428.4]
  assign _T_69271 = select_15 == 6'h26; // @[Switch.scala 41:52:@30430.4]
  assign output_38_15 = io_outValid_15 & _T_69271; // @[Switch.scala 41:38:@30431.4]
  assign _T_69274 = select_16 == 6'h26; // @[Switch.scala 41:52:@30433.4]
  assign output_38_16 = io_outValid_16 & _T_69274; // @[Switch.scala 41:38:@30434.4]
  assign _T_69277 = select_17 == 6'h26; // @[Switch.scala 41:52:@30436.4]
  assign output_38_17 = io_outValid_17 & _T_69277; // @[Switch.scala 41:38:@30437.4]
  assign _T_69280 = select_18 == 6'h26; // @[Switch.scala 41:52:@30439.4]
  assign output_38_18 = io_outValid_18 & _T_69280; // @[Switch.scala 41:38:@30440.4]
  assign _T_69283 = select_19 == 6'h26; // @[Switch.scala 41:52:@30442.4]
  assign output_38_19 = io_outValid_19 & _T_69283; // @[Switch.scala 41:38:@30443.4]
  assign _T_69286 = select_20 == 6'h26; // @[Switch.scala 41:52:@30445.4]
  assign output_38_20 = io_outValid_20 & _T_69286; // @[Switch.scala 41:38:@30446.4]
  assign _T_69289 = select_21 == 6'h26; // @[Switch.scala 41:52:@30448.4]
  assign output_38_21 = io_outValid_21 & _T_69289; // @[Switch.scala 41:38:@30449.4]
  assign _T_69292 = select_22 == 6'h26; // @[Switch.scala 41:52:@30451.4]
  assign output_38_22 = io_outValid_22 & _T_69292; // @[Switch.scala 41:38:@30452.4]
  assign _T_69295 = select_23 == 6'h26; // @[Switch.scala 41:52:@30454.4]
  assign output_38_23 = io_outValid_23 & _T_69295; // @[Switch.scala 41:38:@30455.4]
  assign _T_69298 = select_24 == 6'h26; // @[Switch.scala 41:52:@30457.4]
  assign output_38_24 = io_outValid_24 & _T_69298; // @[Switch.scala 41:38:@30458.4]
  assign _T_69301 = select_25 == 6'h26; // @[Switch.scala 41:52:@30460.4]
  assign output_38_25 = io_outValid_25 & _T_69301; // @[Switch.scala 41:38:@30461.4]
  assign _T_69304 = select_26 == 6'h26; // @[Switch.scala 41:52:@30463.4]
  assign output_38_26 = io_outValid_26 & _T_69304; // @[Switch.scala 41:38:@30464.4]
  assign _T_69307 = select_27 == 6'h26; // @[Switch.scala 41:52:@30466.4]
  assign output_38_27 = io_outValid_27 & _T_69307; // @[Switch.scala 41:38:@30467.4]
  assign _T_69310 = select_28 == 6'h26; // @[Switch.scala 41:52:@30469.4]
  assign output_38_28 = io_outValid_28 & _T_69310; // @[Switch.scala 41:38:@30470.4]
  assign _T_69313 = select_29 == 6'h26; // @[Switch.scala 41:52:@30472.4]
  assign output_38_29 = io_outValid_29 & _T_69313; // @[Switch.scala 41:38:@30473.4]
  assign _T_69316 = select_30 == 6'h26; // @[Switch.scala 41:52:@30475.4]
  assign output_38_30 = io_outValid_30 & _T_69316; // @[Switch.scala 41:38:@30476.4]
  assign _T_69319 = select_31 == 6'h26; // @[Switch.scala 41:52:@30478.4]
  assign output_38_31 = io_outValid_31 & _T_69319; // @[Switch.scala 41:38:@30479.4]
  assign _T_69322 = select_32 == 6'h26; // @[Switch.scala 41:52:@30481.4]
  assign output_38_32 = io_outValid_32 & _T_69322; // @[Switch.scala 41:38:@30482.4]
  assign _T_69325 = select_33 == 6'h26; // @[Switch.scala 41:52:@30484.4]
  assign output_38_33 = io_outValid_33 & _T_69325; // @[Switch.scala 41:38:@30485.4]
  assign _T_69328 = select_34 == 6'h26; // @[Switch.scala 41:52:@30487.4]
  assign output_38_34 = io_outValid_34 & _T_69328; // @[Switch.scala 41:38:@30488.4]
  assign _T_69331 = select_35 == 6'h26; // @[Switch.scala 41:52:@30490.4]
  assign output_38_35 = io_outValid_35 & _T_69331; // @[Switch.scala 41:38:@30491.4]
  assign _T_69334 = select_36 == 6'h26; // @[Switch.scala 41:52:@30493.4]
  assign output_38_36 = io_outValid_36 & _T_69334; // @[Switch.scala 41:38:@30494.4]
  assign _T_69337 = select_37 == 6'h26; // @[Switch.scala 41:52:@30496.4]
  assign output_38_37 = io_outValid_37 & _T_69337; // @[Switch.scala 41:38:@30497.4]
  assign _T_69340 = select_38 == 6'h26; // @[Switch.scala 41:52:@30499.4]
  assign output_38_38 = io_outValid_38 & _T_69340; // @[Switch.scala 41:38:@30500.4]
  assign _T_69343 = select_39 == 6'h26; // @[Switch.scala 41:52:@30502.4]
  assign output_38_39 = io_outValid_39 & _T_69343; // @[Switch.scala 41:38:@30503.4]
  assign _T_69346 = select_40 == 6'h26; // @[Switch.scala 41:52:@30505.4]
  assign output_38_40 = io_outValid_40 & _T_69346; // @[Switch.scala 41:38:@30506.4]
  assign _T_69349 = select_41 == 6'h26; // @[Switch.scala 41:52:@30508.4]
  assign output_38_41 = io_outValid_41 & _T_69349; // @[Switch.scala 41:38:@30509.4]
  assign _T_69352 = select_42 == 6'h26; // @[Switch.scala 41:52:@30511.4]
  assign output_38_42 = io_outValid_42 & _T_69352; // @[Switch.scala 41:38:@30512.4]
  assign _T_69355 = select_43 == 6'h26; // @[Switch.scala 41:52:@30514.4]
  assign output_38_43 = io_outValid_43 & _T_69355; // @[Switch.scala 41:38:@30515.4]
  assign _T_69358 = select_44 == 6'h26; // @[Switch.scala 41:52:@30517.4]
  assign output_38_44 = io_outValid_44 & _T_69358; // @[Switch.scala 41:38:@30518.4]
  assign _T_69361 = select_45 == 6'h26; // @[Switch.scala 41:52:@30520.4]
  assign output_38_45 = io_outValid_45 & _T_69361; // @[Switch.scala 41:38:@30521.4]
  assign _T_69364 = select_46 == 6'h26; // @[Switch.scala 41:52:@30523.4]
  assign output_38_46 = io_outValid_46 & _T_69364; // @[Switch.scala 41:38:@30524.4]
  assign _T_69367 = select_47 == 6'h26; // @[Switch.scala 41:52:@30526.4]
  assign output_38_47 = io_outValid_47 & _T_69367; // @[Switch.scala 41:38:@30527.4]
  assign _T_69370 = select_48 == 6'h26; // @[Switch.scala 41:52:@30529.4]
  assign output_38_48 = io_outValid_48 & _T_69370; // @[Switch.scala 41:38:@30530.4]
  assign _T_69373 = select_49 == 6'h26; // @[Switch.scala 41:52:@30532.4]
  assign output_38_49 = io_outValid_49 & _T_69373; // @[Switch.scala 41:38:@30533.4]
  assign _T_69376 = select_50 == 6'h26; // @[Switch.scala 41:52:@30535.4]
  assign output_38_50 = io_outValid_50 & _T_69376; // @[Switch.scala 41:38:@30536.4]
  assign _T_69379 = select_51 == 6'h26; // @[Switch.scala 41:52:@30538.4]
  assign output_38_51 = io_outValid_51 & _T_69379; // @[Switch.scala 41:38:@30539.4]
  assign _T_69382 = select_52 == 6'h26; // @[Switch.scala 41:52:@30541.4]
  assign output_38_52 = io_outValid_52 & _T_69382; // @[Switch.scala 41:38:@30542.4]
  assign _T_69385 = select_53 == 6'h26; // @[Switch.scala 41:52:@30544.4]
  assign output_38_53 = io_outValid_53 & _T_69385; // @[Switch.scala 41:38:@30545.4]
  assign _T_69388 = select_54 == 6'h26; // @[Switch.scala 41:52:@30547.4]
  assign output_38_54 = io_outValid_54 & _T_69388; // @[Switch.scala 41:38:@30548.4]
  assign _T_69391 = select_55 == 6'h26; // @[Switch.scala 41:52:@30550.4]
  assign output_38_55 = io_outValid_55 & _T_69391; // @[Switch.scala 41:38:@30551.4]
  assign _T_69394 = select_56 == 6'h26; // @[Switch.scala 41:52:@30553.4]
  assign output_38_56 = io_outValid_56 & _T_69394; // @[Switch.scala 41:38:@30554.4]
  assign _T_69397 = select_57 == 6'h26; // @[Switch.scala 41:52:@30556.4]
  assign output_38_57 = io_outValid_57 & _T_69397; // @[Switch.scala 41:38:@30557.4]
  assign _T_69400 = select_58 == 6'h26; // @[Switch.scala 41:52:@30559.4]
  assign output_38_58 = io_outValid_58 & _T_69400; // @[Switch.scala 41:38:@30560.4]
  assign _T_69403 = select_59 == 6'h26; // @[Switch.scala 41:52:@30562.4]
  assign output_38_59 = io_outValid_59 & _T_69403; // @[Switch.scala 41:38:@30563.4]
  assign _T_69406 = select_60 == 6'h26; // @[Switch.scala 41:52:@30565.4]
  assign output_38_60 = io_outValid_60 & _T_69406; // @[Switch.scala 41:38:@30566.4]
  assign _T_69409 = select_61 == 6'h26; // @[Switch.scala 41:52:@30568.4]
  assign output_38_61 = io_outValid_61 & _T_69409; // @[Switch.scala 41:38:@30569.4]
  assign _T_69412 = select_62 == 6'h26; // @[Switch.scala 41:52:@30571.4]
  assign output_38_62 = io_outValid_62 & _T_69412; // @[Switch.scala 41:38:@30572.4]
  assign _T_69415 = select_63 == 6'h26; // @[Switch.scala 41:52:@30574.4]
  assign output_38_63 = io_outValid_63 & _T_69415; // @[Switch.scala 41:38:@30575.4]
  assign _T_69423 = {output_38_7,output_38_6,output_38_5,output_38_4,output_38_3,output_38_2,output_38_1,output_38_0}; // @[Switch.scala 43:31:@30583.4]
  assign _T_69431 = {output_38_15,output_38_14,output_38_13,output_38_12,output_38_11,output_38_10,output_38_9,output_38_8,_T_69423}; // @[Switch.scala 43:31:@30591.4]
  assign _T_69438 = {output_38_23,output_38_22,output_38_21,output_38_20,output_38_19,output_38_18,output_38_17,output_38_16}; // @[Switch.scala 43:31:@30598.4]
  assign _T_69447 = {output_38_31,output_38_30,output_38_29,output_38_28,output_38_27,output_38_26,output_38_25,output_38_24,_T_69438,_T_69431}; // @[Switch.scala 43:31:@30607.4]
  assign _T_69454 = {output_38_39,output_38_38,output_38_37,output_38_36,output_38_35,output_38_34,output_38_33,output_38_32}; // @[Switch.scala 43:31:@30614.4]
  assign _T_69462 = {output_38_47,output_38_46,output_38_45,output_38_44,output_38_43,output_38_42,output_38_41,output_38_40,_T_69454}; // @[Switch.scala 43:31:@30622.4]
  assign _T_69469 = {output_38_55,output_38_54,output_38_53,output_38_52,output_38_51,output_38_50,output_38_49,output_38_48}; // @[Switch.scala 43:31:@30629.4]
  assign _T_69478 = {output_38_63,output_38_62,output_38_61,output_38_60,output_38_59,output_38_58,output_38_57,output_38_56,_T_69469,_T_69462}; // @[Switch.scala 43:31:@30638.4]
  assign _T_69479 = {_T_69478,_T_69447}; // @[Switch.scala 43:31:@30639.4]
  assign _T_69483 = select_0 == 6'h27; // @[Switch.scala 41:52:@30642.4]
  assign output_39_0 = io_outValid_0 & _T_69483; // @[Switch.scala 41:38:@30643.4]
  assign _T_69486 = select_1 == 6'h27; // @[Switch.scala 41:52:@30645.4]
  assign output_39_1 = io_outValid_1 & _T_69486; // @[Switch.scala 41:38:@30646.4]
  assign _T_69489 = select_2 == 6'h27; // @[Switch.scala 41:52:@30648.4]
  assign output_39_2 = io_outValid_2 & _T_69489; // @[Switch.scala 41:38:@30649.4]
  assign _T_69492 = select_3 == 6'h27; // @[Switch.scala 41:52:@30651.4]
  assign output_39_3 = io_outValid_3 & _T_69492; // @[Switch.scala 41:38:@30652.4]
  assign _T_69495 = select_4 == 6'h27; // @[Switch.scala 41:52:@30654.4]
  assign output_39_4 = io_outValid_4 & _T_69495; // @[Switch.scala 41:38:@30655.4]
  assign _T_69498 = select_5 == 6'h27; // @[Switch.scala 41:52:@30657.4]
  assign output_39_5 = io_outValid_5 & _T_69498; // @[Switch.scala 41:38:@30658.4]
  assign _T_69501 = select_6 == 6'h27; // @[Switch.scala 41:52:@30660.4]
  assign output_39_6 = io_outValid_6 & _T_69501; // @[Switch.scala 41:38:@30661.4]
  assign _T_69504 = select_7 == 6'h27; // @[Switch.scala 41:52:@30663.4]
  assign output_39_7 = io_outValid_7 & _T_69504; // @[Switch.scala 41:38:@30664.4]
  assign _T_69507 = select_8 == 6'h27; // @[Switch.scala 41:52:@30666.4]
  assign output_39_8 = io_outValid_8 & _T_69507; // @[Switch.scala 41:38:@30667.4]
  assign _T_69510 = select_9 == 6'h27; // @[Switch.scala 41:52:@30669.4]
  assign output_39_9 = io_outValid_9 & _T_69510; // @[Switch.scala 41:38:@30670.4]
  assign _T_69513 = select_10 == 6'h27; // @[Switch.scala 41:52:@30672.4]
  assign output_39_10 = io_outValid_10 & _T_69513; // @[Switch.scala 41:38:@30673.4]
  assign _T_69516 = select_11 == 6'h27; // @[Switch.scala 41:52:@30675.4]
  assign output_39_11 = io_outValid_11 & _T_69516; // @[Switch.scala 41:38:@30676.4]
  assign _T_69519 = select_12 == 6'h27; // @[Switch.scala 41:52:@30678.4]
  assign output_39_12 = io_outValid_12 & _T_69519; // @[Switch.scala 41:38:@30679.4]
  assign _T_69522 = select_13 == 6'h27; // @[Switch.scala 41:52:@30681.4]
  assign output_39_13 = io_outValid_13 & _T_69522; // @[Switch.scala 41:38:@30682.4]
  assign _T_69525 = select_14 == 6'h27; // @[Switch.scala 41:52:@30684.4]
  assign output_39_14 = io_outValid_14 & _T_69525; // @[Switch.scala 41:38:@30685.4]
  assign _T_69528 = select_15 == 6'h27; // @[Switch.scala 41:52:@30687.4]
  assign output_39_15 = io_outValid_15 & _T_69528; // @[Switch.scala 41:38:@30688.4]
  assign _T_69531 = select_16 == 6'h27; // @[Switch.scala 41:52:@30690.4]
  assign output_39_16 = io_outValid_16 & _T_69531; // @[Switch.scala 41:38:@30691.4]
  assign _T_69534 = select_17 == 6'h27; // @[Switch.scala 41:52:@30693.4]
  assign output_39_17 = io_outValid_17 & _T_69534; // @[Switch.scala 41:38:@30694.4]
  assign _T_69537 = select_18 == 6'h27; // @[Switch.scala 41:52:@30696.4]
  assign output_39_18 = io_outValid_18 & _T_69537; // @[Switch.scala 41:38:@30697.4]
  assign _T_69540 = select_19 == 6'h27; // @[Switch.scala 41:52:@30699.4]
  assign output_39_19 = io_outValid_19 & _T_69540; // @[Switch.scala 41:38:@30700.4]
  assign _T_69543 = select_20 == 6'h27; // @[Switch.scala 41:52:@30702.4]
  assign output_39_20 = io_outValid_20 & _T_69543; // @[Switch.scala 41:38:@30703.4]
  assign _T_69546 = select_21 == 6'h27; // @[Switch.scala 41:52:@30705.4]
  assign output_39_21 = io_outValid_21 & _T_69546; // @[Switch.scala 41:38:@30706.4]
  assign _T_69549 = select_22 == 6'h27; // @[Switch.scala 41:52:@30708.4]
  assign output_39_22 = io_outValid_22 & _T_69549; // @[Switch.scala 41:38:@30709.4]
  assign _T_69552 = select_23 == 6'h27; // @[Switch.scala 41:52:@30711.4]
  assign output_39_23 = io_outValid_23 & _T_69552; // @[Switch.scala 41:38:@30712.4]
  assign _T_69555 = select_24 == 6'h27; // @[Switch.scala 41:52:@30714.4]
  assign output_39_24 = io_outValid_24 & _T_69555; // @[Switch.scala 41:38:@30715.4]
  assign _T_69558 = select_25 == 6'h27; // @[Switch.scala 41:52:@30717.4]
  assign output_39_25 = io_outValid_25 & _T_69558; // @[Switch.scala 41:38:@30718.4]
  assign _T_69561 = select_26 == 6'h27; // @[Switch.scala 41:52:@30720.4]
  assign output_39_26 = io_outValid_26 & _T_69561; // @[Switch.scala 41:38:@30721.4]
  assign _T_69564 = select_27 == 6'h27; // @[Switch.scala 41:52:@30723.4]
  assign output_39_27 = io_outValid_27 & _T_69564; // @[Switch.scala 41:38:@30724.4]
  assign _T_69567 = select_28 == 6'h27; // @[Switch.scala 41:52:@30726.4]
  assign output_39_28 = io_outValid_28 & _T_69567; // @[Switch.scala 41:38:@30727.4]
  assign _T_69570 = select_29 == 6'h27; // @[Switch.scala 41:52:@30729.4]
  assign output_39_29 = io_outValid_29 & _T_69570; // @[Switch.scala 41:38:@30730.4]
  assign _T_69573 = select_30 == 6'h27; // @[Switch.scala 41:52:@30732.4]
  assign output_39_30 = io_outValid_30 & _T_69573; // @[Switch.scala 41:38:@30733.4]
  assign _T_69576 = select_31 == 6'h27; // @[Switch.scala 41:52:@30735.4]
  assign output_39_31 = io_outValid_31 & _T_69576; // @[Switch.scala 41:38:@30736.4]
  assign _T_69579 = select_32 == 6'h27; // @[Switch.scala 41:52:@30738.4]
  assign output_39_32 = io_outValid_32 & _T_69579; // @[Switch.scala 41:38:@30739.4]
  assign _T_69582 = select_33 == 6'h27; // @[Switch.scala 41:52:@30741.4]
  assign output_39_33 = io_outValid_33 & _T_69582; // @[Switch.scala 41:38:@30742.4]
  assign _T_69585 = select_34 == 6'h27; // @[Switch.scala 41:52:@30744.4]
  assign output_39_34 = io_outValid_34 & _T_69585; // @[Switch.scala 41:38:@30745.4]
  assign _T_69588 = select_35 == 6'h27; // @[Switch.scala 41:52:@30747.4]
  assign output_39_35 = io_outValid_35 & _T_69588; // @[Switch.scala 41:38:@30748.4]
  assign _T_69591 = select_36 == 6'h27; // @[Switch.scala 41:52:@30750.4]
  assign output_39_36 = io_outValid_36 & _T_69591; // @[Switch.scala 41:38:@30751.4]
  assign _T_69594 = select_37 == 6'h27; // @[Switch.scala 41:52:@30753.4]
  assign output_39_37 = io_outValid_37 & _T_69594; // @[Switch.scala 41:38:@30754.4]
  assign _T_69597 = select_38 == 6'h27; // @[Switch.scala 41:52:@30756.4]
  assign output_39_38 = io_outValid_38 & _T_69597; // @[Switch.scala 41:38:@30757.4]
  assign _T_69600 = select_39 == 6'h27; // @[Switch.scala 41:52:@30759.4]
  assign output_39_39 = io_outValid_39 & _T_69600; // @[Switch.scala 41:38:@30760.4]
  assign _T_69603 = select_40 == 6'h27; // @[Switch.scala 41:52:@30762.4]
  assign output_39_40 = io_outValid_40 & _T_69603; // @[Switch.scala 41:38:@30763.4]
  assign _T_69606 = select_41 == 6'h27; // @[Switch.scala 41:52:@30765.4]
  assign output_39_41 = io_outValid_41 & _T_69606; // @[Switch.scala 41:38:@30766.4]
  assign _T_69609 = select_42 == 6'h27; // @[Switch.scala 41:52:@30768.4]
  assign output_39_42 = io_outValid_42 & _T_69609; // @[Switch.scala 41:38:@30769.4]
  assign _T_69612 = select_43 == 6'h27; // @[Switch.scala 41:52:@30771.4]
  assign output_39_43 = io_outValid_43 & _T_69612; // @[Switch.scala 41:38:@30772.4]
  assign _T_69615 = select_44 == 6'h27; // @[Switch.scala 41:52:@30774.4]
  assign output_39_44 = io_outValid_44 & _T_69615; // @[Switch.scala 41:38:@30775.4]
  assign _T_69618 = select_45 == 6'h27; // @[Switch.scala 41:52:@30777.4]
  assign output_39_45 = io_outValid_45 & _T_69618; // @[Switch.scala 41:38:@30778.4]
  assign _T_69621 = select_46 == 6'h27; // @[Switch.scala 41:52:@30780.4]
  assign output_39_46 = io_outValid_46 & _T_69621; // @[Switch.scala 41:38:@30781.4]
  assign _T_69624 = select_47 == 6'h27; // @[Switch.scala 41:52:@30783.4]
  assign output_39_47 = io_outValid_47 & _T_69624; // @[Switch.scala 41:38:@30784.4]
  assign _T_69627 = select_48 == 6'h27; // @[Switch.scala 41:52:@30786.4]
  assign output_39_48 = io_outValid_48 & _T_69627; // @[Switch.scala 41:38:@30787.4]
  assign _T_69630 = select_49 == 6'h27; // @[Switch.scala 41:52:@30789.4]
  assign output_39_49 = io_outValid_49 & _T_69630; // @[Switch.scala 41:38:@30790.4]
  assign _T_69633 = select_50 == 6'h27; // @[Switch.scala 41:52:@30792.4]
  assign output_39_50 = io_outValid_50 & _T_69633; // @[Switch.scala 41:38:@30793.4]
  assign _T_69636 = select_51 == 6'h27; // @[Switch.scala 41:52:@30795.4]
  assign output_39_51 = io_outValid_51 & _T_69636; // @[Switch.scala 41:38:@30796.4]
  assign _T_69639 = select_52 == 6'h27; // @[Switch.scala 41:52:@30798.4]
  assign output_39_52 = io_outValid_52 & _T_69639; // @[Switch.scala 41:38:@30799.4]
  assign _T_69642 = select_53 == 6'h27; // @[Switch.scala 41:52:@30801.4]
  assign output_39_53 = io_outValid_53 & _T_69642; // @[Switch.scala 41:38:@30802.4]
  assign _T_69645 = select_54 == 6'h27; // @[Switch.scala 41:52:@30804.4]
  assign output_39_54 = io_outValid_54 & _T_69645; // @[Switch.scala 41:38:@30805.4]
  assign _T_69648 = select_55 == 6'h27; // @[Switch.scala 41:52:@30807.4]
  assign output_39_55 = io_outValid_55 & _T_69648; // @[Switch.scala 41:38:@30808.4]
  assign _T_69651 = select_56 == 6'h27; // @[Switch.scala 41:52:@30810.4]
  assign output_39_56 = io_outValid_56 & _T_69651; // @[Switch.scala 41:38:@30811.4]
  assign _T_69654 = select_57 == 6'h27; // @[Switch.scala 41:52:@30813.4]
  assign output_39_57 = io_outValid_57 & _T_69654; // @[Switch.scala 41:38:@30814.4]
  assign _T_69657 = select_58 == 6'h27; // @[Switch.scala 41:52:@30816.4]
  assign output_39_58 = io_outValid_58 & _T_69657; // @[Switch.scala 41:38:@30817.4]
  assign _T_69660 = select_59 == 6'h27; // @[Switch.scala 41:52:@30819.4]
  assign output_39_59 = io_outValid_59 & _T_69660; // @[Switch.scala 41:38:@30820.4]
  assign _T_69663 = select_60 == 6'h27; // @[Switch.scala 41:52:@30822.4]
  assign output_39_60 = io_outValid_60 & _T_69663; // @[Switch.scala 41:38:@30823.4]
  assign _T_69666 = select_61 == 6'h27; // @[Switch.scala 41:52:@30825.4]
  assign output_39_61 = io_outValid_61 & _T_69666; // @[Switch.scala 41:38:@30826.4]
  assign _T_69669 = select_62 == 6'h27; // @[Switch.scala 41:52:@30828.4]
  assign output_39_62 = io_outValid_62 & _T_69669; // @[Switch.scala 41:38:@30829.4]
  assign _T_69672 = select_63 == 6'h27; // @[Switch.scala 41:52:@30831.4]
  assign output_39_63 = io_outValid_63 & _T_69672; // @[Switch.scala 41:38:@30832.4]
  assign _T_69680 = {output_39_7,output_39_6,output_39_5,output_39_4,output_39_3,output_39_2,output_39_1,output_39_0}; // @[Switch.scala 43:31:@30840.4]
  assign _T_69688 = {output_39_15,output_39_14,output_39_13,output_39_12,output_39_11,output_39_10,output_39_9,output_39_8,_T_69680}; // @[Switch.scala 43:31:@30848.4]
  assign _T_69695 = {output_39_23,output_39_22,output_39_21,output_39_20,output_39_19,output_39_18,output_39_17,output_39_16}; // @[Switch.scala 43:31:@30855.4]
  assign _T_69704 = {output_39_31,output_39_30,output_39_29,output_39_28,output_39_27,output_39_26,output_39_25,output_39_24,_T_69695,_T_69688}; // @[Switch.scala 43:31:@30864.4]
  assign _T_69711 = {output_39_39,output_39_38,output_39_37,output_39_36,output_39_35,output_39_34,output_39_33,output_39_32}; // @[Switch.scala 43:31:@30871.4]
  assign _T_69719 = {output_39_47,output_39_46,output_39_45,output_39_44,output_39_43,output_39_42,output_39_41,output_39_40,_T_69711}; // @[Switch.scala 43:31:@30879.4]
  assign _T_69726 = {output_39_55,output_39_54,output_39_53,output_39_52,output_39_51,output_39_50,output_39_49,output_39_48}; // @[Switch.scala 43:31:@30886.4]
  assign _T_69735 = {output_39_63,output_39_62,output_39_61,output_39_60,output_39_59,output_39_58,output_39_57,output_39_56,_T_69726,_T_69719}; // @[Switch.scala 43:31:@30895.4]
  assign _T_69736 = {_T_69735,_T_69704}; // @[Switch.scala 43:31:@30896.4]
  assign _T_69740 = select_0 == 6'h28; // @[Switch.scala 41:52:@30899.4]
  assign output_40_0 = io_outValid_0 & _T_69740; // @[Switch.scala 41:38:@30900.4]
  assign _T_69743 = select_1 == 6'h28; // @[Switch.scala 41:52:@30902.4]
  assign output_40_1 = io_outValid_1 & _T_69743; // @[Switch.scala 41:38:@30903.4]
  assign _T_69746 = select_2 == 6'h28; // @[Switch.scala 41:52:@30905.4]
  assign output_40_2 = io_outValid_2 & _T_69746; // @[Switch.scala 41:38:@30906.4]
  assign _T_69749 = select_3 == 6'h28; // @[Switch.scala 41:52:@30908.4]
  assign output_40_3 = io_outValid_3 & _T_69749; // @[Switch.scala 41:38:@30909.4]
  assign _T_69752 = select_4 == 6'h28; // @[Switch.scala 41:52:@30911.4]
  assign output_40_4 = io_outValid_4 & _T_69752; // @[Switch.scala 41:38:@30912.4]
  assign _T_69755 = select_5 == 6'h28; // @[Switch.scala 41:52:@30914.4]
  assign output_40_5 = io_outValid_5 & _T_69755; // @[Switch.scala 41:38:@30915.4]
  assign _T_69758 = select_6 == 6'h28; // @[Switch.scala 41:52:@30917.4]
  assign output_40_6 = io_outValid_6 & _T_69758; // @[Switch.scala 41:38:@30918.4]
  assign _T_69761 = select_7 == 6'h28; // @[Switch.scala 41:52:@30920.4]
  assign output_40_7 = io_outValid_7 & _T_69761; // @[Switch.scala 41:38:@30921.4]
  assign _T_69764 = select_8 == 6'h28; // @[Switch.scala 41:52:@30923.4]
  assign output_40_8 = io_outValid_8 & _T_69764; // @[Switch.scala 41:38:@30924.4]
  assign _T_69767 = select_9 == 6'h28; // @[Switch.scala 41:52:@30926.4]
  assign output_40_9 = io_outValid_9 & _T_69767; // @[Switch.scala 41:38:@30927.4]
  assign _T_69770 = select_10 == 6'h28; // @[Switch.scala 41:52:@30929.4]
  assign output_40_10 = io_outValid_10 & _T_69770; // @[Switch.scala 41:38:@30930.4]
  assign _T_69773 = select_11 == 6'h28; // @[Switch.scala 41:52:@30932.4]
  assign output_40_11 = io_outValid_11 & _T_69773; // @[Switch.scala 41:38:@30933.4]
  assign _T_69776 = select_12 == 6'h28; // @[Switch.scala 41:52:@30935.4]
  assign output_40_12 = io_outValid_12 & _T_69776; // @[Switch.scala 41:38:@30936.4]
  assign _T_69779 = select_13 == 6'h28; // @[Switch.scala 41:52:@30938.4]
  assign output_40_13 = io_outValid_13 & _T_69779; // @[Switch.scala 41:38:@30939.4]
  assign _T_69782 = select_14 == 6'h28; // @[Switch.scala 41:52:@30941.4]
  assign output_40_14 = io_outValid_14 & _T_69782; // @[Switch.scala 41:38:@30942.4]
  assign _T_69785 = select_15 == 6'h28; // @[Switch.scala 41:52:@30944.4]
  assign output_40_15 = io_outValid_15 & _T_69785; // @[Switch.scala 41:38:@30945.4]
  assign _T_69788 = select_16 == 6'h28; // @[Switch.scala 41:52:@30947.4]
  assign output_40_16 = io_outValid_16 & _T_69788; // @[Switch.scala 41:38:@30948.4]
  assign _T_69791 = select_17 == 6'h28; // @[Switch.scala 41:52:@30950.4]
  assign output_40_17 = io_outValid_17 & _T_69791; // @[Switch.scala 41:38:@30951.4]
  assign _T_69794 = select_18 == 6'h28; // @[Switch.scala 41:52:@30953.4]
  assign output_40_18 = io_outValid_18 & _T_69794; // @[Switch.scala 41:38:@30954.4]
  assign _T_69797 = select_19 == 6'h28; // @[Switch.scala 41:52:@30956.4]
  assign output_40_19 = io_outValid_19 & _T_69797; // @[Switch.scala 41:38:@30957.4]
  assign _T_69800 = select_20 == 6'h28; // @[Switch.scala 41:52:@30959.4]
  assign output_40_20 = io_outValid_20 & _T_69800; // @[Switch.scala 41:38:@30960.4]
  assign _T_69803 = select_21 == 6'h28; // @[Switch.scala 41:52:@30962.4]
  assign output_40_21 = io_outValid_21 & _T_69803; // @[Switch.scala 41:38:@30963.4]
  assign _T_69806 = select_22 == 6'h28; // @[Switch.scala 41:52:@30965.4]
  assign output_40_22 = io_outValid_22 & _T_69806; // @[Switch.scala 41:38:@30966.4]
  assign _T_69809 = select_23 == 6'h28; // @[Switch.scala 41:52:@30968.4]
  assign output_40_23 = io_outValid_23 & _T_69809; // @[Switch.scala 41:38:@30969.4]
  assign _T_69812 = select_24 == 6'h28; // @[Switch.scala 41:52:@30971.4]
  assign output_40_24 = io_outValid_24 & _T_69812; // @[Switch.scala 41:38:@30972.4]
  assign _T_69815 = select_25 == 6'h28; // @[Switch.scala 41:52:@30974.4]
  assign output_40_25 = io_outValid_25 & _T_69815; // @[Switch.scala 41:38:@30975.4]
  assign _T_69818 = select_26 == 6'h28; // @[Switch.scala 41:52:@30977.4]
  assign output_40_26 = io_outValid_26 & _T_69818; // @[Switch.scala 41:38:@30978.4]
  assign _T_69821 = select_27 == 6'h28; // @[Switch.scala 41:52:@30980.4]
  assign output_40_27 = io_outValid_27 & _T_69821; // @[Switch.scala 41:38:@30981.4]
  assign _T_69824 = select_28 == 6'h28; // @[Switch.scala 41:52:@30983.4]
  assign output_40_28 = io_outValid_28 & _T_69824; // @[Switch.scala 41:38:@30984.4]
  assign _T_69827 = select_29 == 6'h28; // @[Switch.scala 41:52:@30986.4]
  assign output_40_29 = io_outValid_29 & _T_69827; // @[Switch.scala 41:38:@30987.4]
  assign _T_69830 = select_30 == 6'h28; // @[Switch.scala 41:52:@30989.4]
  assign output_40_30 = io_outValid_30 & _T_69830; // @[Switch.scala 41:38:@30990.4]
  assign _T_69833 = select_31 == 6'h28; // @[Switch.scala 41:52:@30992.4]
  assign output_40_31 = io_outValid_31 & _T_69833; // @[Switch.scala 41:38:@30993.4]
  assign _T_69836 = select_32 == 6'h28; // @[Switch.scala 41:52:@30995.4]
  assign output_40_32 = io_outValid_32 & _T_69836; // @[Switch.scala 41:38:@30996.4]
  assign _T_69839 = select_33 == 6'h28; // @[Switch.scala 41:52:@30998.4]
  assign output_40_33 = io_outValid_33 & _T_69839; // @[Switch.scala 41:38:@30999.4]
  assign _T_69842 = select_34 == 6'h28; // @[Switch.scala 41:52:@31001.4]
  assign output_40_34 = io_outValid_34 & _T_69842; // @[Switch.scala 41:38:@31002.4]
  assign _T_69845 = select_35 == 6'h28; // @[Switch.scala 41:52:@31004.4]
  assign output_40_35 = io_outValid_35 & _T_69845; // @[Switch.scala 41:38:@31005.4]
  assign _T_69848 = select_36 == 6'h28; // @[Switch.scala 41:52:@31007.4]
  assign output_40_36 = io_outValid_36 & _T_69848; // @[Switch.scala 41:38:@31008.4]
  assign _T_69851 = select_37 == 6'h28; // @[Switch.scala 41:52:@31010.4]
  assign output_40_37 = io_outValid_37 & _T_69851; // @[Switch.scala 41:38:@31011.4]
  assign _T_69854 = select_38 == 6'h28; // @[Switch.scala 41:52:@31013.4]
  assign output_40_38 = io_outValid_38 & _T_69854; // @[Switch.scala 41:38:@31014.4]
  assign _T_69857 = select_39 == 6'h28; // @[Switch.scala 41:52:@31016.4]
  assign output_40_39 = io_outValid_39 & _T_69857; // @[Switch.scala 41:38:@31017.4]
  assign _T_69860 = select_40 == 6'h28; // @[Switch.scala 41:52:@31019.4]
  assign output_40_40 = io_outValid_40 & _T_69860; // @[Switch.scala 41:38:@31020.4]
  assign _T_69863 = select_41 == 6'h28; // @[Switch.scala 41:52:@31022.4]
  assign output_40_41 = io_outValid_41 & _T_69863; // @[Switch.scala 41:38:@31023.4]
  assign _T_69866 = select_42 == 6'h28; // @[Switch.scala 41:52:@31025.4]
  assign output_40_42 = io_outValid_42 & _T_69866; // @[Switch.scala 41:38:@31026.4]
  assign _T_69869 = select_43 == 6'h28; // @[Switch.scala 41:52:@31028.4]
  assign output_40_43 = io_outValid_43 & _T_69869; // @[Switch.scala 41:38:@31029.4]
  assign _T_69872 = select_44 == 6'h28; // @[Switch.scala 41:52:@31031.4]
  assign output_40_44 = io_outValid_44 & _T_69872; // @[Switch.scala 41:38:@31032.4]
  assign _T_69875 = select_45 == 6'h28; // @[Switch.scala 41:52:@31034.4]
  assign output_40_45 = io_outValid_45 & _T_69875; // @[Switch.scala 41:38:@31035.4]
  assign _T_69878 = select_46 == 6'h28; // @[Switch.scala 41:52:@31037.4]
  assign output_40_46 = io_outValid_46 & _T_69878; // @[Switch.scala 41:38:@31038.4]
  assign _T_69881 = select_47 == 6'h28; // @[Switch.scala 41:52:@31040.4]
  assign output_40_47 = io_outValid_47 & _T_69881; // @[Switch.scala 41:38:@31041.4]
  assign _T_69884 = select_48 == 6'h28; // @[Switch.scala 41:52:@31043.4]
  assign output_40_48 = io_outValid_48 & _T_69884; // @[Switch.scala 41:38:@31044.4]
  assign _T_69887 = select_49 == 6'h28; // @[Switch.scala 41:52:@31046.4]
  assign output_40_49 = io_outValid_49 & _T_69887; // @[Switch.scala 41:38:@31047.4]
  assign _T_69890 = select_50 == 6'h28; // @[Switch.scala 41:52:@31049.4]
  assign output_40_50 = io_outValid_50 & _T_69890; // @[Switch.scala 41:38:@31050.4]
  assign _T_69893 = select_51 == 6'h28; // @[Switch.scala 41:52:@31052.4]
  assign output_40_51 = io_outValid_51 & _T_69893; // @[Switch.scala 41:38:@31053.4]
  assign _T_69896 = select_52 == 6'h28; // @[Switch.scala 41:52:@31055.4]
  assign output_40_52 = io_outValid_52 & _T_69896; // @[Switch.scala 41:38:@31056.4]
  assign _T_69899 = select_53 == 6'h28; // @[Switch.scala 41:52:@31058.4]
  assign output_40_53 = io_outValid_53 & _T_69899; // @[Switch.scala 41:38:@31059.4]
  assign _T_69902 = select_54 == 6'h28; // @[Switch.scala 41:52:@31061.4]
  assign output_40_54 = io_outValid_54 & _T_69902; // @[Switch.scala 41:38:@31062.4]
  assign _T_69905 = select_55 == 6'h28; // @[Switch.scala 41:52:@31064.4]
  assign output_40_55 = io_outValid_55 & _T_69905; // @[Switch.scala 41:38:@31065.4]
  assign _T_69908 = select_56 == 6'h28; // @[Switch.scala 41:52:@31067.4]
  assign output_40_56 = io_outValid_56 & _T_69908; // @[Switch.scala 41:38:@31068.4]
  assign _T_69911 = select_57 == 6'h28; // @[Switch.scala 41:52:@31070.4]
  assign output_40_57 = io_outValid_57 & _T_69911; // @[Switch.scala 41:38:@31071.4]
  assign _T_69914 = select_58 == 6'h28; // @[Switch.scala 41:52:@31073.4]
  assign output_40_58 = io_outValid_58 & _T_69914; // @[Switch.scala 41:38:@31074.4]
  assign _T_69917 = select_59 == 6'h28; // @[Switch.scala 41:52:@31076.4]
  assign output_40_59 = io_outValid_59 & _T_69917; // @[Switch.scala 41:38:@31077.4]
  assign _T_69920 = select_60 == 6'h28; // @[Switch.scala 41:52:@31079.4]
  assign output_40_60 = io_outValid_60 & _T_69920; // @[Switch.scala 41:38:@31080.4]
  assign _T_69923 = select_61 == 6'h28; // @[Switch.scala 41:52:@31082.4]
  assign output_40_61 = io_outValid_61 & _T_69923; // @[Switch.scala 41:38:@31083.4]
  assign _T_69926 = select_62 == 6'h28; // @[Switch.scala 41:52:@31085.4]
  assign output_40_62 = io_outValid_62 & _T_69926; // @[Switch.scala 41:38:@31086.4]
  assign _T_69929 = select_63 == 6'h28; // @[Switch.scala 41:52:@31088.4]
  assign output_40_63 = io_outValid_63 & _T_69929; // @[Switch.scala 41:38:@31089.4]
  assign _T_69937 = {output_40_7,output_40_6,output_40_5,output_40_4,output_40_3,output_40_2,output_40_1,output_40_0}; // @[Switch.scala 43:31:@31097.4]
  assign _T_69945 = {output_40_15,output_40_14,output_40_13,output_40_12,output_40_11,output_40_10,output_40_9,output_40_8,_T_69937}; // @[Switch.scala 43:31:@31105.4]
  assign _T_69952 = {output_40_23,output_40_22,output_40_21,output_40_20,output_40_19,output_40_18,output_40_17,output_40_16}; // @[Switch.scala 43:31:@31112.4]
  assign _T_69961 = {output_40_31,output_40_30,output_40_29,output_40_28,output_40_27,output_40_26,output_40_25,output_40_24,_T_69952,_T_69945}; // @[Switch.scala 43:31:@31121.4]
  assign _T_69968 = {output_40_39,output_40_38,output_40_37,output_40_36,output_40_35,output_40_34,output_40_33,output_40_32}; // @[Switch.scala 43:31:@31128.4]
  assign _T_69976 = {output_40_47,output_40_46,output_40_45,output_40_44,output_40_43,output_40_42,output_40_41,output_40_40,_T_69968}; // @[Switch.scala 43:31:@31136.4]
  assign _T_69983 = {output_40_55,output_40_54,output_40_53,output_40_52,output_40_51,output_40_50,output_40_49,output_40_48}; // @[Switch.scala 43:31:@31143.4]
  assign _T_69992 = {output_40_63,output_40_62,output_40_61,output_40_60,output_40_59,output_40_58,output_40_57,output_40_56,_T_69983,_T_69976}; // @[Switch.scala 43:31:@31152.4]
  assign _T_69993 = {_T_69992,_T_69961}; // @[Switch.scala 43:31:@31153.4]
  assign _T_69997 = select_0 == 6'h29; // @[Switch.scala 41:52:@31156.4]
  assign output_41_0 = io_outValid_0 & _T_69997; // @[Switch.scala 41:38:@31157.4]
  assign _T_70000 = select_1 == 6'h29; // @[Switch.scala 41:52:@31159.4]
  assign output_41_1 = io_outValid_1 & _T_70000; // @[Switch.scala 41:38:@31160.4]
  assign _T_70003 = select_2 == 6'h29; // @[Switch.scala 41:52:@31162.4]
  assign output_41_2 = io_outValid_2 & _T_70003; // @[Switch.scala 41:38:@31163.4]
  assign _T_70006 = select_3 == 6'h29; // @[Switch.scala 41:52:@31165.4]
  assign output_41_3 = io_outValid_3 & _T_70006; // @[Switch.scala 41:38:@31166.4]
  assign _T_70009 = select_4 == 6'h29; // @[Switch.scala 41:52:@31168.4]
  assign output_41_4 = io_outValid_4 & _T_70009; // @[Switch.scala 41:38:@31169.4]
  assign _T_70012 = select_5 == 6'h29; // @[Switch.scala 41:52:@31171.4]
  assign output_41_5 = io_outValid_5 & _T_70012; // @[Switch.scala 41:38:@31172.4]
  assign _T_70015 = select_6 == 6'h29; // @[Switch.scala 41:52:@31174.4]
  assign output_41_6 = io_outValid_6 & _T_70015; // @[Switch.scala 41:38:@31175.4]
  assign _T_70018 = select_7 == 6'h29; // @[Switch.scala 41:52:@31177.4]
  assign output_41_7 = io_outValid_7 & _T_70018; // @[Switch.scala 41:38:@31178.4]
  assign _T_70021 = select_8 == 6'h29; // @[Switch.scala 41:52:@31180.4]
  assign output_41_8 = io_outValid_8 & _T_70021; // @[Switch.scala 41:38:@31181.4]
  assign _T_70024 = select_9 == 6'h29; // @[Switch.scala 41:52:@31183.4]
  assign output_41_9 = io_outValid_9 & _T_70024; // @[Switch.scala 41:38:@31184.4]
  assign _T_70027 = select_10 == 6'h29; // @[Switch.scala 41:52:@31186.4]
  assign output_41_10 = io_outValid_10 & _T_70027; // @[Switch.scala 41:38:@31187.4]
  assign _T_70030 = select_11 == 6'h29; // @[Switch.scala 41:52:@31189.4]
  assign output_41_11 = io_outValid_11 & _T_70030; // @[Switch.scala 41:38:@31190.4]
  assign _T_70033 = select_12 == 6'h29; // @[Switch.scala 41:52:@31192.4]
  assign output_41_12 = io_outValid_12 & _T_70033; // @[Switch.scala 41:38:@31193.4]
  assign _T_70036 = select_13 == 6'h29; // @[Switch.scala 41:52:@31195.4]
  assign output_41_13 = io_outValid_13 & _T_70036; // @[Switch.scala 41:38:@31196.4]
  assign _T_70039 = select_14 == 6'h29; // @[Switch.scala 41:52:@31198.4]
  assign output_41_14 = io_outValid_14 & _T_70039; // @[Switch.scala 41:38:@31199.4]
  assign _T_70042 = select_15 == 6'h29; // @[Switch.scala 41:52:@31201.4]
  assign output_41_15 = io_outValid_15 & _T_70042; // @[Switch.scala 41:38:@31202.4]
  assign _T_70045 = select_16 == 6'h29; // @[Switch.scala 41:52:@31204.4]
  assign output_41_16 = io_outValid_16 & _T_70045; // @[Switch.scala 41:38:@31205.4]
  assign _T_70048 = select_17 == 6'h29; // @[Switch.scala 41:52:@31207.4]
  assign output_41_17 = io_outValid_17 & _T_70048; // @[Switch.scala 41:38:@31208.4]
  assign _T_70051 = select_18 == 6'h29; // @[Switch.scala 41:52:@31210.4]
  assign output_41_18 = io_outValid_18 & _T_70051; // @[Switch.scala 41:38:@31211.4]
  assign _T_70054 = select_19 == 6'h29; // @[Switch.scala 41:52:@31213.4]
  assign output_41_19 = io_outValid_19 & _T_70054; // @[Switch.scala 41:38:@31214.4]
  assign _T_70057 = select_20 == 6'h29; // @[Switch.scala 41:52:@31216.4]
  assign output_41_20 = io_outValid_20 & _T_70057; // @[Switch.scala 41:38:@31217.4]
  assign _T_70060 = select_21 == 6'h29; // @[Switch.scala 41:52:@31219.4]
  assign output_41_21 = io_outValid_21 & _T_70060; // @[Switch.scala 41:38:@31220.4]
  assign _T_70063 = select_22 == 6'h29; // @[Switch.scala 41:52:@31222.4]
  assign output_41_22 = io_outValid_22 & _T_70063; // @[Switch.scala 41:38:@31223.4]
  assign _T_70066 = select_23 == 6'h29; // @[Switch.scala 41:52:@31225.4]
  assign output_41_23 = io_outValid_23 & _T_70066; // @[Switch.scala 41:38:@31226.4]
  assign _T_70069 = select_24 == 6'h29; // @[Switch.scala 41:52:@31228.4]
  assign output_41_24 = io_outValid_24 & _T_70069; // @[Switch.scala 41:38:@31229.4]
  assign _T_70072 = select_25 == 6'h29; // @[Switch.scala 41:52:@31231.4]
  assign output_41_25 = io_outValid_25 & _T_70072; // @[Switch.scala 41:38:@31232.4]
  assign _T_70075 = select_26 == 6'h29; // @[Switch.scala 41:52:@31234.4]
  assign output_41_26 = io_outValid_26 & _T_70075; // @[Switch.scala 41:38:@31235.4]
  assign _T_70078 = select_27 == 6'h29; // @[Switch.scala 41:52:@31237.4]
  assign output_41_27 = io_outValid_27 & _T_70078; // @[Switch.scala 41:38:@31238.4]
  assign _T_70081 = select_28 == 6'h29; // @[Switch.scala 41:52:@31240.4]
  assign output_41_28 = io_outValid_28 & _T_70081; // @[Switch.scala 41:38:@31241.4]
  assign _T_70084 = select_29 == 6'h29; // @[Switch.scala 41:52:@31243.4]
  assign output_41_29 = io_outValid_29 & _T_70084; // @[Switch.scala 41:38:@31244.4]
  assign _T_70087 = select_30 == 6'h29; // @[Switch.scala 41:52:@31246.4]
  assign output_41_30 = io_outValid_30 & _T_70087; // @[Switch.scala 41:38:@31247.4]
  assign _T_70090 = select_31 == 6'h29; // @[Switch.scala 41:52:@31249.4]
  assign output_41_31 = io_outValid_31 & _T_70090; // @[Switch.scala 41:38:@31250.4]
  assign _T_70093 = select_32 == 6'h29; // @[Switch.scala 41:52:@31252.4]
  assign output_41_32 = io_outValid_32 & _T_70093; // @[Switch.scala 41:38:@31253.4]
  assign _T_70096 = select_33 == 6'h29; // @[Switch.scala 41:52:@31255.4]
  assign output_41_33 = io_outValid_33 & _T_70096; // @[Switch.scala 41:38:@31256.4]
  assign _T_70099 = select_34 == 6'h29; // @[Switch.scala 41:52:@31258.4]
  assign output_41_34 = io_outValid_34 & _T_70099; // @[Switch.scala 41:38:@31259.4]
  assign _T_70102 = select_35 == 6'h29; // @[Switch.scala 41:52:@31261.4]
  assign output_41_35 = io_outValid_35 & _T_70102; // @[Switch.scala 41:38:@31262.4]
  assign _T_70105 = select_36 == 6'h29; // @[Switch.scala 41:52:@31264.4]
  assign output_41_36 = io_outValid_36 & _T_70105; // @[Switch.scala 41:38:@31265.4]
  assign _T_70108 = select_37 == 6'h29; // @[Switch.scala 41:52:@31267.4]
  assign output_41_37 = io_outValid_37 & _T_70108; // @[Switch.scala 41:38:@31268.4]
  assign _T_70111 = select_38 == 6'h29; // @[Switch.scala 41:52:@31270.4]
  assign output_41_38 = io_outValid_38 & _T_70111; // @[Switch.scala 41:38:@31271.4]
  assign _T_70114 = select_39 == 6'h29; // @[Switch.scala 41:52:@31273.4]
  assign output_41_39 = io_outValid_39 & _T_70114; // @[Switch.scala 41:38:@31274.4]
  assign _T_70117 = select_40 == 6'h29; // @[Switch.scala 41:52:@31276.4]
  assign output_41_40 = io_outValid_40 & _T_70117; // @[Switch.scala 41:38:@31277.4]
  assign _T_70120 = select_41 == 6'h29; // @[Switch.scala 41:52:@31279.4]
  assign output_41_41 = io_outValid_41 & _T_70120; // @[Switch.scala 41:38:@31280.4]
  assign _T_70123 = select_42 == 6'h29; // @[Switch.scala 41:52:@31282.4]
  assign output_41_42 = io_outValid_42 & _T_70123; // @[Switch.scala 41:38:@31283.4]
  assign _T_70126 = select_43 == 6'h29; // @[Switch.scala 41:52:@31285.4]
  assign output_41_43 = io_outValid_43 & _T_70126; // @[Switch.scala 41:38:@31286.4]
  assign _T_70129 = select_44 == 6'h29; // @[Switch.scala 41:52:@31288.4]
  assign output_41_44 = io_outValid_44 & _T_70129; // @[Switch.scala 41:38:@31289.4]
  assign _T_70132 = select_45 == 6'h29; // @[Switch.scala 41:52:@31291.4]
  assign output_41_45 = io_outValid_45 & _T_70132; // @[Switch.scala 41:38:@31292.4]
  assign _T_70135 = select_46 == 6'h29; // @[Switch.scala 41:52:@31294.4]
  assign output_41_46 = io_outValid_46 & _T_70135; // @[Switch.scala 41:38:@31295.4]
  assign _T_70138 = select_47 == 6'h29; // @[Switch.scala 41:52:@31297.4]
  assign output_41_47 = io_outValid_47 & _T_70138; // @[Switch.scala 41:38:@31298.4]
  assign _T_70141 = select_48 == 6'h29; // @[Switch.scala 41:52:@31300.4]
  assign output_41_48 = io_outValid_48 & _T_70141; // @[Switch.scala 41:38:@31301.4]
  assign _T_70144 = select_49 == 6'h29; // @[Switch.scala 41:52:@31303.4]
  assign output_41_49 = io_outValid_49 & _T_70144; // @[Switch.scala 41:38:@31304.4]
  assign _T_70147 = select_50 == 6'h29; // @[Switch.scala 41:52:@31306.4]
  assign output_41_50 = io_outValid_50 & _T_70147; // @[Switch.scala 41:38:@31307.4]
  assign _T_70150 = select_51 == 6'h29; // @[Switch.scala 41:52:@31309.4]
  assign output_41_51 = io_outValid_51 & _T_70150; // @[Switch.scala 41:38:@31310.4]
  assign _T_70153 = select_52 == 6'h29; // @[Switch.scala 41:52:@31312.4]
  assign output_41_52 = io_outValid_52 & _T_70153; // @[Switch.scala 41:38:@31313.4]
  assign _T_70156 = select_53 == 6'h29; // @[Switch.scala 41:52:@31315.4]
  assign output_41_53 = io_outValid_53 & _T_70156; // @[Switch.scala 41:38:@31316.4]
  assign _T_70159 = select_54 == 6'h29; // @[Switch.scala 41:52:@31318.4]
  assign output_41_54 = io_outValid_54 & _T_70159; // @[Switch.scala 41:38:@31319.4]
  assign _T_70162 = select_55 == 6'h29; // @[Switch.scala 41:52:@31321.4]
  assign output_41_55 = io_outValid_55 & _T_70162; // @[Switch.scala 41:38:@31322.4]
  assign _T_70165 = select_56 == 6'h29; // @[Switch.scala 41:52:@31324.4]
  assign output_41_56 = io_outValid_56 & _T_70165; // @[Switch.scala 41:38:@31325.4]
  assign _T_70168 = select_57 == 6'h29; // @[Switch.scala 41:52:@31327.4]
  assign output_41_57 = io_outValid_57 & _T_70168; // @[Switch.scala 41:38:@31328.4]
  assign _T_70171 = select_58 == 6'h29; // @[Switch.scala 41:52:@31330.4]
  assign output_41_58 = io_outValid_58 & _T_70171; // @[Switch.scala 41:38:@31331.4]
  assign _T_70174 = select_59 == 6'h29; // @[Switch.scala 41:52:@31333.4]
  assign output_41_59 = io_outValid_59 & _T_70174; // @[Switch.scala 41:38:@31334.4]
  assign _T_70177 = select_60 == 6'h29; // @[Switch.scala 41:52:@31336.4]
  assign output_41_60 = io_outValid_60 & _T_70177; // @[Switch.scala 41:38:@31337.4]
  assign _T_70180 = select_61 == 6'h29; // @[Switch.scala 41:52:@31339.4]
  assign output_41_61 = io_outValid_61 & _T_70180; // @[Switch.scala 41:38:@31340.4]
  assign _T_70183 = select_62 == 6'h29; // @[Switch.scala 41:52:@31342.4]
  assign output_41_62 = io_outValid_62 & _T_70183; // @[Switch.scala 41:38:@31343.4]
  assign _T_70186 = select_63 == 6'h29; // @[Switch.scala 41:52:@31345.4]
  assign output_41_63 = io_outValid_63 & _T_70186; // @[Switch.scala 41:38:@31346.4]
  assign _T_70194 = {output_41_7,output_41_6,output_41_5,output_41_4,output_41_3,output_41_2,output_41_1,output_41_0}; // @[Switch.scala 43:31:@31354.4]
  assign _T_70202 = {output_41_15,output_41_14,output_41_13,output_41_12,output_41_11,output_41_10,output_41_9,output_41_8,_T_70194}; // @[Switch.scala 43:31:@31362.4]
  assign _T_70209 = {output_41_23,output_41_22,output_41_21,output_41_20,output_41_19,output_41_18,output_41_17,output_41_16}; // @[Switch.scala 43:31:@31369.4]
  assign _T_70218 = {output_41_31,output_41_30,output_41_29,output_41_28,output_41_27,output_41_26,output_41_25,output_41_24,_T_70209,_T_70202}; // @[Switch.scala 43:31:@31378.4]
  assign _T_70225 = {output_41_39,output_41_38,output_41_37,output_41_36,output_41_35,output_41_34,output_41_33,output_41_32}; // @[Switch.scala 43:31:@31385.4]
  assign _T_70233 = {output_41_47,output_41_46,output_41_45,output_41_44,output_41_43,output_41_42,output_41_41,output_41_40,_T_70225}; // @[Switch.scala 43:31:@31393.4]
  assign _T_70240 = {output_41_55,output_41_54,output_41_53,output_41_52,output_41_51,output_41_50,output_41_49,output_41_48}; // @[Switch.scala 43:31:@31400.4]
  assign _T_70249 = {output_41_63,output_41_62,output_41_61,output_41_60,output_41_59,output_41_58,output_41_57,output_41_56,_T_70240,_T_70233}; // @[Switch.scala 43:31:@31409.4]
  assign _T_70250 = {_T_70249,_T_70218}; // @[Switch.scala 43:31:@31410.4]
  assign _T_70254 = select_0 == 6'h2a; // @[Switch.scala 41:52:@31413.4]
  assign output_42_0 = io_outValid_0 & _T_70254; // @[Switch.scala 41:38:@31414.4]
  assign _T_70257 = select_1 == 6'h2a; // @[Switch.scala 41:52:@31416.4]
  assign output_42_1 = io_outValid_1 & _T_70257; // @[Switch.scala 41:38:@31417.4]
  assign _T_70260 = select_2 == 6'h2a; // @[Switch.scala 41:52:@31419.4]
  assign output_42_2 = io_outValid_2 & _T_70260; // @[Switch.scala 41:38:@31420.4]
  assign _T_70263 = select_3 == 6'h2a; // @[Switch.scala 41:52:@31422.4]
  assign output_42_3 = io_outValid_3 & _T_70263; // @[Switch.scala 41:38:@31423.4]
  assign _T_70266 = select_4 == 6'h2a; // @[Switch.scala 41:52:@31425.4]
  assign output_42_4 = io_outValid_4 & _T_70266; // @[Switch.scala 41:38:@31426.4]
  assign _T_70269 = select_5 == 6'h2a; // @[Switch.scala 41:52:@31428.4]
  assign output_42_5 = io_outValid_5 & _T_70269; // @[Switch.scala 41:38:@31429.4]
  assign _T_70272 = select_6 == 6'h2a; // @[Switch.scala 41:52:@31431.4]
  assign output_42_6 = io_outValid_6 & _T_70272; // @[Switch.scala 41:38:@31432.4]
  assign _T_70275 = select_7 == 6'h2a; // @[Switch.scala 41:52:@31434.4]
  assign output_42_7 = io_outValid_7 & _T_70275; // @[Switch.scala 41:38:@31435.4]
  assign _T_70278 = select_8 == 6'h2a; // @[Switch.scala 41:52:@31437.4]
  assign output_42_8 = io_outValid_8 & _T_70278; // @[Switch.scala 41:38:@31438.4]
  assign _T_70281 = select_9 == 6'h2a; // @[Switch.scala 41:52:@31440.4]
  assign output_42_9 = io_outValid_9 & _T_70281; // @[Switch.scala 41:38:@31441.4]
  assign _T_70284 = select_10 == 6'h2a; // @[Switch.scala 41:52:@31443.4]
  assign output_42_10 = io_outValid_10 & _T_70284; // @[Switch.scala 41:38:@31444.4]
  assign _T_70287 = select_11 == 6'h2a; // @[Switch.scala 41:52:@31446.4]
  assign output_42_11 = io_outValid_11 & _T_70287; // @[Switch.scala 41:38:@31447.4]
  assign _T_70290 = select_12 == 6'h2a; // @[Switch.scala 41:52:@31449.4]
  assign output_42_12 = io_outValid_12 & _T_70290; // @[Switch.scala 41:38:@31450.4]
  assign _T_70293 = select_13 == 6'h2a; // @[Switch.scala 41:52:@31452.4]
  assign output_42_13 = io_outValid_13 & _T_70293; // @[Switch.scala 41:38:@31453.4]
  assign _T_70296 = select_14 == 6'h2a; // @[Switch.scala 41:52:@31455.4]
  assign output_42_14 = io_outValid_14 & _T_70296; // @[Switch.scala 41:38:@31456.4]
  assign _T_70299 = select_15 == 6'h2a; // @[Switch.scala 41:52:@31458.4]
  assign output_42_15 = io_outValid_15 & _T_70299; // @[Switch.scala 41:38:@31459.4]
  assign _T_70302 = select_16 == 6'h2a; // @[Switch.scala 41:52:@31461.4]
  assign output_42_16 = io_outValid_16 & _T_70302; // @[Switch.scala 41:38:@31462.4]
  assign _T_70305 = select_17 == 6'h2a; // @[Switch.scala 41:52:@31464.4]
  assign output_42_17 = io_outValid_17 & _T_70305; // @[Switch.scala 41:38:@31465.4]
  assign _T_70308 = select_18 == 6'h2a; // @[Switch.scala 41:52:@31467.4]
  assign output_42_18 = io_outValid_18 & _T_70308; // @[Switch.scala 41:38:@31468.4]
  assign _T_70311 = select_19 == 6'h2a; // @[Switch.scala 41:52:@31470.4]
  assign output_42_19 = io_outValid_19 & _T_70311; // @[Switch.scala 41:38:@31471.4]
  assign _T_70314 = select_20 == 6'h2a; // @[Switch.scala 41:52:@31473.4]
  assign output_42_20 = io_outValid_20 & _T_70314; // @[Switch.scala 41:38:@31474.4]
  assign _T_70317 = select_21 == 6'h2a; // @[Switch.scala 41:52:@31476.4]
  assign output_42_21 = io_outValid_21 & _T_70317; // @[Switch.scala 41:38:@31477.4]
  assign _T_70320 = select_22 == 6'h2a; // @[Switch.scala 41:52:@31479.4]
  assign output_42_22 = io_outValid_22 & _T_70320; // @[Switch.scala 41:38:@31480.4]
  assign _T_70323 = select_23 == 6'h2a; // @[Switch.scala 41:52:@31482.4]
  assign output_42_23 = io_outValid_23 & _T_70323; // @[Switch.scala 41:38:@31483.4]
  assign _T_70326 = select_24 == 6'h2a; // @[Switch.scala 41:52:@31485.4]
  assign output_42_24 = io_outValid_24 & _T_70326; // @[Switch.scala 41:38:@31486.4]
  assign _T_70329 = select_25 == 6'h2a; // @[Switch.scala 41:52:@31488.4]
  assign output_42_25 = io_outValid_25 & _T_70329; // @[Switch.scala 41:38:@31489.4]
  assign _T_70332 = select_26 == 6'h2a; // @[Switch.scala 41:52:@31491.4]
  assign output_42_26 = io_outValid_26 & _T_70332; // @[Switch.scala 41:38:@31492.4]
  assign _T_70335 = select_27 == 6'h2a; // @[Switch.scala 41:52:@31494.4]
  assign output_42_27 = io_outValid_27 & _T_70335; // @[Switch.scala 41:38:@31495.4]
  assign _T_70338 = select_28 == 6'h2a; // @[Switch.scala 41:52:@31497.4]
  assign output_42_28 = io_outValid_28 & _T_70338; // @[Switch.scala 41:38:@31498.4]
  assign _T_70341 = select_29 == 6'h2a; // @[Switch.scala 41:52:@31500.4]
  assign output_42_29 = io_outValid_29 & _T_70341; // @[Switch.scala 41:38:@31501.4]
  assign _T_70344 = select_30 == 6'h2a; // @[Switch.scala 41:52:@31503.4]
  assign output_42_30 = io_outValid_30 & _T_70344; // @[Switch.scala 41:38:@31504.4]
  assign _T_70347 = select_31 == 6'h2a; // @[Switch.scala 41:52:@31506.4]
  assign output_42_31 = io_outValid_31 & _T_70347; // @[Switch.scala 41:38:@31507.4]
  assign _T_70350 = select_32 == 6'h2a; // @[Switch.scala 41:52:@31509.4]
  assign output_42_32 = io_outValid_32 & _T_70350; // @[Switch.scala 41:38:@31510.4]
  assign _T_70353 = select_33 == 6'h2a; // @[Switch.scala 41:52:@31512.4]
  assign output_42_33 = io_outValid_33 & _T_70353; // @[Switch.scala 41:38:@31513.4]
  assign _T_70356 = select_34 == 6'h2a; // @[Switch.scala 41:52:@31515.4]
  assign output_42_34 = io_outValid_34 & _T_70356; // @[Switch.scala 41:38:@31516.4]
  assign _T_70359 = select_35 == 6'h2a; // @[Switch.scala 41:52:@31518.4]
  assign output_42_35 = io_outValid_35 & _T_70359; // @[Switch.scala 41:38:@31519.4]
  assign _T_70362 = select_36 == 6'h2a; // @[Switch.scala 41:52:@31521.4]
  assign output_42_36 = io_outValid_36 & _T_70362; // @[Switch.scala 41:38:@31522.4]
  assign _T_70365 = select_37 == 6'h2a; // @[Switch.scala 41:52:@31524.4]
  assign output_42_37 = io_outValid_37 & _T_70365; // @[Switch.scala 41:38:@31525.4]
  assign _T_70368 = select_38 == 6'h2a; // @[Switch.scala 41:52:@31527.4]
  assign output_42_38 = io_outValid_38 & _T_70368; // @[Switch.scala 41:38:@31528.4]
  assign _T_70371 = select_39 == 6'h2a; // @[Switch.scala 41:52:@31530.4]
  assign output_42_39 = io_outValid_39 & _T_70371; // @[Switch.scala 41:38:@31531.4]
  assign _T_70374 = select_40 == 6'h2a; // @[Switch.scala 41:52:@31533.4]
  assign output_42_40 = io_outValid_40 & _T_70374; // @[Switch.scala 41:38:@31534.4]
  assign _T_70377 = select_41 == 6'h2a; // @[Switch.scala 41:52:@31536.4]
  assign output_42_41 = io_outValid_41 & _T_70377; // @[Switch.scala 41:38:@31537.4]
  assign _T_70380 = select_42 == 6'h2a; // @[Switch.scala 41:52:@31539.4]
  assign output_42_42 = io_outValid_42 & _T_70380; // @[Switch.scala 41:38:@31540.4]
  assign _T_70383 = select_43 == 6'h2a; // @[Switch.scala 41:52:@31542.4]
  assign output_42_43 = io_outValid_43 & _T_70383; // @[Switch.scala 41:38:@31543.4]
  assign _T_70386 = select_44 == 6'h2a; // @[Switch.scala 41:52:@31545.4]
  assign output_42_44 = io_outValid_44 & _T_70386; // @[Switch.scala 41:38:@31546.4]
  assign _T_70389 = select_45 == 6'h2a; // @[Switch.scala 41:52:@31548.4]
  assign output_42_45 = io_outValid_45 & _T_70389; // @[Switch.scala 41:38:@31549.4]
  assign _T_70392 = select_46 == 6'h2a; // @[Switch.scala 41:52:@31551.4]
  assign output_42_46 = io_outValid_46 & _T_70392; // @[Switch.scala 41:38:@31552.4]
  assign _T_70395 = select_47 == 6'h2a; // @[Switch.scala 41:52:@31554.4]
  assign output_42_47 = io_outValid_47 & _T_70395; // @[Switch.scala 41:38:@31555.4]
  assign _T_70398 = select_48 == 6'h2a; // @[Switch.scala 41:52:@31557.4]
  assign output_42_48 = io_outValid_48 & _T_70398; // @[Switch.scala 41:38:@31558.4]
  assign _T_70401 = select_49 == 6'h2a; // @[Switch.scala 41:52:@31560.4]
  assign output_42_49 = io_outValid_49 & _T_70401; // @[Switch.scala 41:38:@31561.4]
  assign _T_70404 = select_50 == 6'h2a; // @[Switch.scala 41:52:@31563.4]
  assign output_42_50 = io_outValid_50 & _T_70404; // @[Switch.scala 41:38:@31564.4]
  assign _T_70407 = select_51 == 6'h2a; // @[Switch.scala 41:52:@31566.4]
  assign output_42_51 = io_outValid_51 & _T_70407; // @[Switch.scala 41:38:@31567.4]
  assign _T_70410 = select_52 == 6'h2a; // @[Switch.scala 41:52:@31569.4]
  assign output_42_52 = io_outValid_52 & _T_70410; // @[Switch.scala 41:38:@31570.4]
  assign _T_70413 = select_53 == 6'h2a; // @[Switch.scala 41:52:@31572.4]
  assign output_42_53 = io_outValid_53 & _T_70413; // @[Switch.scala 41:38:@31573.4]
  assign _T_70416 = select_54 == 6'h2a; // @[Switch.scala 41:52:@31575.4]
  assign output_42_54 = io_outValid_54 & _T_70416; // @[Switch.scala 41:38:@31576.4]
  assign _T_70419 = select_55 == 6'h2a; // @[Switch.scala 41:52:@31578.4]
  assign output_42_55 = io_outValid_55 & _T_70419; // @[Switch.scala 41:38:@31579.4]
  assign _T_70422 = select_56 == 6'h2a; // @[Switch.scala 41:52:@31581.4]
  assign output_42_56 = io_outValid_56 & _T_70422; // @[Switch.scala 41:38:@31582.4]
  assign _T_70425 = select_57 == 6'h2a; // @[Switch.scala 41:52:@31584.4]
  assign output_42_57 = io_outValid_57 & _T_70425; // @[Switch.scala 41:38:@31585.4]
  assign _T_70428 = select_58 == 6'h2a; // @[Switch.scala 41:52:@31587.4]
  assign output_42_58 = io_outValid_58 & _T_70428; // @[Switch.scala 41:38:@31588.4]
  assign _T_70431 = select_59 == 6'h2a; // @[Switch.scala 41:52:@31590.4]
  assign output_42_59 = io_outValid_59 & _T_70431; // @[Switch.scala 41:38:@31591.4]
  assign _T_70434 = select_60 == 6'h2a; // @[Switch.scala 41:52:@31593.4]
  assign output_42_60 = io_outValid_60 & _T_70434; // @[Switch.scala 41:38:@31594.4]
  assign _T_70437 = select_61 == 6'h2a; // @[Switch.scala 41:52:@31596.4]
  assign output_42_61 = io_outValid_61 & _T_70437; // @[Switch.scala 41:38:@31597.4]
  assign _T_70440 = select_62 == 6'h2a; // @[Switch.scala 41:52:@31599.4]
  assign output_42_62 = io_outValid_62 & _T_70440; // @[Switch.scala 41:38:@31600.4]
  assign _T_70443 = select_63 == 6'h2a; // @[Switch.scala 41:52:@31602.4]
  assign output_42_63 = io_outValid_63 & _T_70443; // @[Switch.scala 41:38:@31603.4]
  assign _T_70451 = {output_42_7,output_42_6,output_42_5,output_42_4,output_42_3,output_42_2,output_42_1,output_42_0}; // @[Switch.scala 43:31:@31611.4]
  assign _T_70459 = {output_42_15,output_42_14,output_42_13,output_42_12,output_42_11,output_42_10,output_42_9,output_42_8,_T_70451}; // @[Switch.scala 43:31:@31619.4]
  assign _T_70466 = {output_42_23,output_42_22,output_42_21,output_42_20,output_42_19,output_42_18,output_42_17,output_42_16}; // @[Switch.scala 43:31:@31626.4]
  assign _T_70475 = {output_42_31,output_42_30,output_42_29,output_42_28,output_42_27,output_42_26,output_42_25,output_42_24,_T_70466,_T_70459}; // @[Switch.scala 43:31:@31635.4]
  assign _T_70482 = {output_42_39,output_42_38,output_42_37,output_42_36,output_42_35,output_42_34,output_42_33,output_42_32}; // @[Switch.scala 43:31:@31642.4]
  assign _T_70490 = {output_42_47,output_42_46,output_42_45,output_42_44,output_42_43,output_42_42,output_42_41,output_42_40,_T_70482}; // @[Switch.scala 43:31:@31650.4]
  assign _T_70497 = {output_42_55,output_42_54,output_42_53,output_42_52,output_42_51,output_42_50,output_42_49,output_42_48}; // @[Switch.scala 43:31:@31657.4]
  assign _T_70506 = {output_42_63,output_42_62,output_42_61,output_42_60,output_42_59,output_42_58,output_42_57,output_42_56,_T_70497,_T_70490}; // @[Switch.scala 43:31:@31666.4]
  assign _T_70507 = {_T_70506,_T_70475}; // @[Switch.scala 43:31:@31667.4]
  assign _T_70511 = select_0 == 6'h2b; // @[Switch.scala 41:52:@31670.4]
  assign output_43_0 = io_outValid_0 & _T_70511; // @[Switch.scala 41:38:@31671.4]
  assign _T_70514 = select_1 == 6'h2b; // @[Switch.scala 41:52:@31673.4]
  assign output_43_1 = io_outValid_1 & _T_70514; // @[Switch.scala 41:38:@31674.4]
  assign _T_70517 = select_2 == 6'h2b; // @[Switch.scala 41:52:@31676.4]
  assign output_43_2 = io_outValid_2 & _T_70517; // @[Switch.scala 41:38:@31677.4]
  assign _T_70520 = select_3 == 6'h2b; // @[Switch.scala 41:52:@31679.4]
  assign output_43_3 = io_outValid_3 & _T_70520; // @[Switch.scala 41:38:@31680.4]
  assign _T_70523 = select_4 == 6'h2b; // @[Switch.scala 41:52:@31682.4]
  assign output_43_4 = io_outValid_4 & _T_70523; // @[Switch.scala 41:38:@31683.4]
  assign _T_70526 = select_5 == 6'h2b; // @[Switch.scala 41:52:@31685.4]
  assign output_43_5 = io_outValid_5 & _T_70526; // @[Switch.scala 41:38:@31686.4]
  assign _T_70529 = select_6 == 6'h2b; // @[Switch.scala 41:52:@31688.4]
  assign output_43_6 = io_outValid_6 & _T_70529; // @[Switch.scala 41:38:@31689.4]
  assign _T_70532 = select_7 == 6'h2b; // @[Switch.scala 41:52:@31691.4]
  assign output_43_7 = io_outValid_7 & _T_70532; // @[Switch.scala 41:38:@31692.4]
  assign _T_70535 = select_8 == 6'h2b; // @[Switch.scala 41:52:@31694.4]
  assign output_43_8 = io_outValid_8 & _T_70535; // @[Switch.scala 41:38:@31695.4]
  assign _T_70538 = select_9 == 6'h2b; // @[Switch.scala 41:52:@31697.4]
  assign output_43_9 = io_outValid_9 & _T_70538; // @[Switch.scala 41:38:@31698.4]
  assign _T_70541 = select_10 == 6'h2b; // @[Switch.scala 41:52:@31700.4]
  assign output_43_10 = io_outValid_10 & _T_70541; // @[Switch.scala 41:38:@31701.4]
  assign _T_70544 = select_11 == 6'h2b; // @[Switch.scala 41:52:@31703.4]
  assign output_43_11 = io_outValid_11 & _T_70544; // @[Switch.scala 41:38:@31704.4]
  assign _T_70547 = select_12 == 6'h2b; // @[Switch.scala 41:52:@31706.4]
  assign output_43_12 = io_outValid_12 & _T_70547; // @[Switch.scala 41:38:@31707.4]
  assign _T_70550 = select_13 == 6'h2b; // @[Switch.scala 41:52:@31709.4]
  assign output_43_13 = io_outValid_13 & _T_70550; // @[Switch.scala 41:38:@31710.4]
  assign _T_70553 = select_14 == 6'h2b; // @[Switch.scala 41:52:@31712.4]
  assign output_43_14 = io_outValid_14 & _T_70553; // @[Switch.scala 41:38:@31713.4]
  assign _T_70556 = select_15 == 6'h2b; // @[Switch.scala 41:52:@31715.4]
  assign output_43_15 = io_outValid_15 & _T_70556; // @[Switch.scala 41:38:@31716.4]
  assign _T_70559 = select_16 == 6'h2b; // @[Switch.scala 41:52:@31718.4]
  assign output_43_16 = io_outValid_16 & _T_70559; // @[Switch.scala 41:38:@31719.4]
  assign _T_70562 = select_17 == 6'h2b; // @[Switch.scala 41:52:@31721.4]
  assign output_43_17 = io_outValid_17 & _T_70562; // @[Switch.scala 41:38:@31722.4]
  assign _T_70565 = select_18 == 6'h2b; // @[Switch.scala 41:52:@31724.4]
  assign output_43_18 = io_outValid_18 & _T_70565; // @[Switch.scala 41:38:@31725.4]
  assign _T_70568 = select_19 == 6'h2b; // @[Switch.scala 41:52:@31727.4]
  assign output_43_19 = io_outValid_19 & _T_70568; // @[Switch.scala 41:38:@31728.4]
  assign _T_70571 = select_20 == 6'h2b; // @[Switch.scala 41:52:@31730.4]
  assign output_43_20 = io_outValid_20 & _T_70571; // @[Switch.scala 41:38:@31731.4]
  assign _T_70574 = select_21 == 6'h2b; // @[Switch.scala 41:52:@31733.4]
  assign output_43_21 = io_outValid_21 & _T_70574; // @[Switch.scala 41:38:@31734.4]
  assign _T_70577 = select_22 == 6'h2b; // @[Switch.scala 41:52:@31736.4]
  assign output_43_22 = io_outValid_22 & _T_70577; // @[Switch.scala 41:38:@31737.4]
  assign _T_70580 = select_23 == 6'h2b; // @[Switch.scala 41:52:@31739.4]
  assign output_43_23 = io_outValid_23 & _T_70580; // @[Switch.scala 41:38:@31740.4]
  assign _T_70583 = select_24 == 6'h2b; // @[Switch.scala 41:52:@31742.4]
  assign output_43_24 = io_outValid_24 & _T_70583; // @[Switch.scala 41:38:@31743.4]
  assign _T_70586 = select_25 == 6'h2b; // @[Switch.scala 41:52:@31745.4]
  assign output_43_25 = io_outValid_25 & _T_70586; // @[Switch.scala 41:38:@31746.4]
  assign _T_70589 = select_26 == 6'h2b; // @[Switch.scala 41:52:@31748.4]
  assign output_43_26 = io_outValid_26 & _T_70589; // @[Switch.scala 41:38:@31749.4]
  assign _T_70592 = select_27 == 6'h2b; // @[Switch.scala 41:52:@31751.4]
  assign output_43_27 = io_outValid_27 & _T_70592; // @[Switch.scala 41:38:@31752.4]
  assign _T_70595 = select_28 == 6'h2b; // @[Switch.scala 41:52:@31754.4]
  assign output_43_28 = io_outValid_28 & _T_70595; // @[Switch.scala 41:38:@31755.4]
  assign _T_70598 = select_29 == 6'h2b; // @[Switch.scala 41:52:@31757.4]
  assign output_43_29 = io_outValid_29 & _T_70598; // @[Switch.scala 41:38:@31758.4]
  assign _T_70601 = select_30 == 6'h2b; // @[Switch.scala 41:52:@31760.4]
  assign output_43_30 = io_outValid_30 & _T_70601; // @[Switch.scala 41:38:@31761.4]
  assign _T_70604 = select_31 == 6'h2b; // @[Switch.scala 41:52:@31763.4]
  assign output_43_31 = io_outValid_31 & _T_70604; // @[Switch.scala 41:38:@31764.4]
  assign _T_70607 = select_32 == 6'h2b; // @[Switch.scala 41:52:@31766.4]
  assign output_43_32 = io_outValid_32 & _T_70607; // @[Switch.scala 41:38:@31767.4]
  assign _T_70610 = select_33 == 6'h2b; // @[Switch.scala 41:52:@31769.4]
  assign output_43_33 = io_outValid_33 & _T_70610; // @[Switch.scala 41:38:@31770.4]
  assign _T_70613 = select_34 == 6'h2b; // @[Switch.scala 41:52:@31772.4]
  assign output_43_34 = io_outValid_34 & _T_70613; // @[Switch.scala 41:38:@31773.4]
  assign _T_70616 = select_35 == 6'h2b; // @[Switch.scala 41:52:@31775.4]
  assign output_43_35 = io_outValid_35 & _T_70616; // @[Switch.scala 41:38:@31776.4]
  assign _T_70619 = select_36 == 6'h2b; // @[Switch.scala 41:52:@31778.4]
  assign output_43_36 = io_outValid_36 & _T_70619; // @[Switch.scala 41:38:@31779.4]
  assign _T_70622 = select_37 == 6'h2b; // @[Switch.scala 41:52:@31781.4]
  assign output_43_37 = io_outValid_37 & _T_70622; // @[Switch.scala 41:38:@31782.4]
  assign _T_70625 = select_38 == 6'h2b; // @[Switch.scala 41:52:@31784.4]
  assign output_43_38 = io_outValid_38 & _T_70625; // @[Switch.scala 41:38:@31785.4]
  assign _T_70628 = select_39 == 6'h2b; // @[Switch.scala 41:52:@31787.4]
  assign output_43_39 = io_outValid_39 & _T_70628; // @[Switch.scala 41:38:@31788.4]
  assign _T_70631 = select_40 == 6'h2b; // @[Switch.scala 41:52:@31790.4]
  assign output_43_40 = io_outValid_40 & _T_70631; // @[Switch.scala 41:38:@31791.4]
  assign _T_70634 = select_41 == 6'h2b; // @[Switch.scala 41:52:@31793.4]
  assign output_43_41 = io_outValid_41 & _T_70634; // @[Switch.scala 41:38:@31794.4]
  assign _T_70637 = select_42 == 6'h2b; // @[Switch.scala 41:52:@31796.4]
  assign output_43_42 = io_outValid_42 & _T_70637; // @[Switch.scala 41:38:@31797.4]
  assign _T_70640 = select_43 == 6'h2b; // @[Switch.scala 41:52:@31799.4]
  assign output_43_43 = io_outValid_43 & _T_70640; // @[Switch.scala 41:38:@31800.4]
  assign _T_70643 = select_44 == 6'h2b; // @[Switch.scala 41:52:@31802.4]
  assign output_43_44 = io_outValid_44 & _T_70643; // @[Switch.scala 41:38:@31803.4]
  assign _T_70646 = select_45 == 6'h2b; // @[Switch.scala 41:52:@31805.4]
  assign output_43_45 = io_outValid_45 & _T_70646; // @[Switch.scala 41:38:@31806.4]
  assign _T_70649 = select_46 == 6'h2b; // @[Switch.scala 41:52:@31808.4]
  assign output_43_46 = io_outValid_46 & _T_70649; // @[Switch.scala 41:38:@31809.4]
  assign _T_70652 = select_47 == 6'h2b; // @[Switch.scala 41:52:@31811.4]
  assign output_43_47 = io_outValid_47 & _T_70652; // @[Switch.scala 41:38:@31812.4]
  assign _T_70655 = select_48 == 6'h2b; // @[Switch.scala 41:52:@31814.4]
  assign output_43_48 = io_outValid_48 & _T_70655; // @[Switch.scala 41:38:@31815.4]
  assign _T_70658 = select_49 == 6'h2b; // @[Switch.scala 41:52:@31817.4]
  assign output_43_49 = io_outValid_49 & _T_70658; // @[Switch.scala 41:38:@31818.4]
  assign _T_70661 = select_50 == 6'h2b; // @[Switch.scala 41:52:@31820.4]
  assign output_43_50 = io_outValid_50 & _T_70661; // @[Switch.scala 41:38:@31821.4]
  assign _T_70664 = select_51 == 6'h2b; // @[Switch.scala 41:52:@31823.4]
  assign output_43_51 = io_outValid_51 & _T_70664; // @[Switch.scala 41:38:@31824.4]
  assign _T_70667 = select_52 == 6'h2b; // @[Switch.scala 41:52:@31826.4]
  assign output_43_52 = io_outValid_52 & _T_70667; // @[Switch.scala 41:38:@31827.4]
  assign _T_70670 = select_53 == 6'h2b; // @[Switch.scala 41:52:@31829.4]
  assign output_43_53 = io_outValid_53 & _T_70670; // @[Switch.scala 41:38:@31830.4]
  assign _T_70673 = select_54 == 6'h2b; // @[Switch.scala 41:52:@31832.4]
  assign output_43_54 = io_outValid_54 & _T_70673; // @[Switch.scala 41:38:@31833.4]
  assign _T_70676 = select_55 == 6'h2b; // @[Switch.scala 41:52:@31835.4]
  assign output_43_55 = io_outValid_55 & _T_70676; // @[Switch.scala 41:38:@31836.4]
  assign _T_70679 = select_56 == 6'h2b; // @[Switch.scala 41:52:@31838.4]
  assign output_43_56 = io_outValid_56 & _T_70679; // @[Switch.scala 41:38:@31839.4]
  assign _T_70682 = select_57 == 6'h2b; // @[Switch.scala 41:52:@31841.4]
  assign output_43_57 = io_outValid_57 & _T_70682; // @[Switch.scala 41:38:@31842.4]
  assign _T_70685 = select_58 == 6'h2b; // @[Switch.scala 41:52:@31844.4]
  assign output_43_58 = io_outValid_58 & _T_70685; // @[Switch.scala 41:38:@31845.4]
  assign _T_70688 = select_59 == 6'h2b; // @[Switch.scala 41:52:@31847.4]
  assign output_43_59 = io_outValid_59 & _T_70688; // @[Switch.scala 41:38:@31848.4]
  assign _T_70691 = select_60 == 6'h2b; // @[Switch.scala 41:52:@31850.4]
  assign output_43_60 = io_outValid_60 & _T_70691; // @[Switch.scala 41:38:@31851.4]
  assign _T_70694 = select_61 == 6'h2b; // @[Switch.scala 41:52:@31853.4]
  assign output_43_61 = io_outValid_61 & _T_70694; // @[Switch.scala 41:38:@31854.4]
  assign _T_70697 = select_62 == 6'h2b; // @[Switch.scala 41:52:@31856.4]
  assign output_43_62 = io_outValid_62 & _T_70697; // @[Switch.scala 41:38:@31857.4]
  assign _T_70700 = select_63 == 6'h2b; // @[Switch.scala 41:52:@31859.4]
  assign output_43_63 = io_outValid_63 & _T_70700; // @[Switch.scala 41:38:@31860.4]
  assign _T_70708 = {output_43_7,output_43_6,output_43_5,output_43_4,output_43_3,output_43_2,output_43_1,output_43_0}; // @[Switch.scala 43:31:@31868.4]
  assign _T_70716 = {output_43_15,output_43_14,output_43_13,output_43_12,output_43_11,output_43_10,output_43_9,output_43_8,_T_70708}; // @[Switch.scala 43:31:@31876.4]
  assign _T_70723 = {output_43_23,output_43_22,output_43_21,output_43_20,output_43_19,output_43_18,output_43_17,output_43_16}; // @[Switch.scala 43:31:@31883.4]
  assign _T_70732 = {output_43_31,output_43_30,output_43_29,output_43_28,output_43_27,output_43_26,output_43_25,output_43_24,_T_70723,_T_70716}; // @[Switch.scala 43:31:@31892.4]
  assign _T_70739 = {output_43_39,output_43_38,output_43_37,output_43_36,output_43_35,output_43_34,output_43_33,output_43_32}; // @[Switch.scala 43:31:@31899.4]
  assign _T_70747 = {output_43_47,output_43_46,output_43_45,output_43_44,output_43_43,output_43_42,output_43_41,output_43_40,_T_70739}; // @[Switch.scala 43:31:@31907.4]
  assign _T_70754 = {output_43_55,output_43_54,output_43_53,output_43_52,output_43_51,output_43_50,output_43_49,output_43_48}; // @[Switch.scala 43:31:@31914.4]
  assign _T_70763 = {output_43_63,output_43_62,output_43_61,output_43_60,output_43_59,output_43_58,output_43_57,output_43_56,_T_70754,_T_70747}; // @[Switch.scala 43:31:@31923.4]
  assign _T_70764 = {_T_70763,_T_70732}; // @[Switch.scala 43:31:@31924.4]
  assign _T_70768 = select_0 == 6'h2c; // @[Switch.scala 41:52:@31927.4]
  assign output_44_0 = io_outValid_0 & _T_70768; // @[Switch.scala 41:38:@31928.4]
  assign _T_70771 = select_1 == 6'h2c; // @[Switch.scala 41:52:@31930.4]
  assign output_44_1 = io_outValid_1 & _T_70771; // @[Switch.scala 41:38:@31931.4]
  assign _T_70774 = select_2 == 6'h2c; // @[Switch.scala 41:52:@31933.4]
  assign output_44_2 = io_outValid_2 & _T_70774; // @[Switch.scala 41:38:@31934.4]
  assign _T_70777 = select_3 == 6'h2c; // @[Switch.scala 41:52:@31936.4]
  assign output_44_3 = io_outValid_3 & _T_70777; // @[Switch.scala 41:38:@31937.4]
  assign _T_70780 = select_4 == 6'h2c; // @[Switch.scala 41:52:@31939.4]
  assign output_44_4 = io_outValid_4 & _T_70780; // @[Switch.scala 41:38:@31940.4]
  assign _T_70783 = select_5 == 6'h2c; // @[Switch.scala 41:52:@31942.4]
  assign output_44_5 = io_outValid_5 & _T_70783; // @[Switch.scala 41:38:@31943.4]
  assign _T_70786 = select_6 == 6'h2c; // @[Switch.scala 41:52:@31945.4]
  assign output_44_6 = io_outValid_6 & _T_70786; // @[Switch.scala 41:38:@31946.4]
  assign _T_70789 = select_7 == 6'h2c; // @[Switch.scala 41:52:@31948.4]
  assign output_44_7 = io_outValid_7 & _T_70789; // @[Switch.scala 41:38:@31949.4]
  assign _T_70792 = select_8 == 6'h2c; // @[Switch.scala 41:52:@31951.4]
  assign output_44_8 = io_outValid_8 & _T_70792; // @[Switch.scala 41:38:@31952.4]
  assign _T_70795 = select_9 == 6'h2c; // @[Switch.scala 41:52:@31954.4]
  assign output_44_9 = io_outValid_9 & _T_70795; // @[Switch.scala 41:38:@31955.4]
  assign _T_70798 = select_10 == 6'h2c; // @[Switch.scala 41:52:@31957.4]
  assign output_44_10 = io_outValid_10 & _T_70798; // @[Switch.scala 41:38:@31958.4]
  assign _T_70801 = select_11 == 6'h2c; // @[Switch.scala 41:52:@31960.4]
  assign output_44_11 = io_outValid_11 & _T_70801; // @[Switch.scala 41:38:@31961.4]
  assign _T_70804 = select_12 == 6'h2c; // @[Switch.scala 41:52:@31963.4]
  assign output_44_12 = io_outValid_12 & _T_70804; // @[Switch.scala 41:38:@31964.4]
  assign _T_70807 = select_13 == 6'h2c; // @[Switch.scala 41:52:@31966.4]
  assign output_44_13 = io_outValid_13 & _T_70807; // @[Switch.scala 41:38:@31967.4]
  assign _T_70810 = select_14 == 6'h2c; // @[Switch.scala 41:52:@31969.4]
  assign output_44_14 = io_outValid_14 & _T_70810; // @[Switch.scala 41:38:@31970.4]
  assign _T_70813 = select_15 == 6'h2c; // @[Switch.scala 41:52:@31972.4]
  assign output_44_15 = io_outValid_15 & _T_70813; // @[Switch.scala 41:38:@31973.4]
  assign _T_70816 = select_16 == 6'h2c; // @[Switch.scala 41:52:@31975.4]
  assign output_44_16 = io_outValid_16 & _T_70816; // @[Switch.scala 41:38:@31976.4]
  assign _T_70819 = select_17 == 6'h2c; // @[Switch.scala 41:52:@31978.4]
  assign output_44_17 = io_outValid_17 & _T_70819; // @[Switch.scala 41:38:@31979.4]
  assign _T_70822 = select_18 == 6'h2c; // @[Switch.scala 41:52:@31981.4]
  assign output_44_18 = io_outValid_18 & _T_70822; // @[Switch.scala 41:38:@31982.4]
  assign _T_70825 = select_19 == 6'h2c; // @[Switch.scala 41:52:@31984.4]
  assign output_44_19 = io_outValid_19 & _T_70825; // @[Switch.scala 41:38:@31985.4]
  assign _T_70828 = select_20 == 6'h2c; // @[Switch.scala 41:52:@31987.4]
  assign output_44_20 = io_outValid_20 & _T_70828; // @[Switch.scala 41:38:@31988.4]
  assign _T_70831 = select_21 == 6'h2c; // @[Switch.scala 41:52:@31990.4]
  assign output_44_21 = io_outValid_21 & _T_70831; // @[Switch.scala 41:38:@31991.4]
  assign _T_70834 = select_22 == 6'h2c; // @[Switch.scala 41:52:@31993.4]
  assign output_44_22 = io_outValid_22 & _T_70834; // @[Switch.scala 41:38:@31994.4]
  assign _T_70837 = select_23 == 6'h2c; // @[Switch.scala 41:52:@31996.4]
  assign output_44_23 = io_outValid_23 & _T_70837; // @[Switch.scala 41:38:@31997.4]
  assign _T_70840 = select_24 == 6'h2c; // @[Switch.scala 41:52:@31999.4]
  assign output_44_24 = io_outValid_24 & _T_70840; // @[Switch.scala 41:38:@32000.4]
  assign _T_70843 = select_25 == 6'h2c; // @[Switch.scala 41:52:@32002.4]
  assign output_44_25 = io_outValid_25 & _T_70843; // @[Switch.scala 41:38:@32003.4]
  assign _T_70846 = select_26 == 6'h2c; // @[Switch.scala 41:52:@32005.4]
  assign output_44_26 = io_outValid_26 & _T_70846; // @[Switch.scala 41:38:@32006.4]
  assign _T_70849 = select_27 == 6'h2c; // @[Switch.scala 41:52:@32008.4]
  assign output_44_27 = io_outValid_27 & _T_70849; // @[Switch.scala 41:38:@32009.4]
  assign _T_70852 = select_28 == 6'h2c; // @[Switch.scala 41:52:@32011.4]
  assign output_44_28 = io_outValid_28 & _T_70852; // @[Switch.scala 41:38:@32012.4]
  assign _T_70855 = select_29 == 6'h2c; // @[Switch.scala 41:52:@32014.4]
  assign output_44_29 = io_outValid_29 & _T_70855; // @[Switch.scala 41:38:@32015.4]
  assign _T_70858 = select_30 == 6'h2c; // @[Switch.scala 41:52:@32017.4]
  assign output_44_30 = io_outValid_30 & _T_70858; // @[Switch.scala 41:38:@32018.4]
  assign _T_70861 = select_31 == 6'h2c; // @[Switch.scala 41:52:@32020.4]
  assign output_44_31 = io_outValid_31 & _T_70861; // @[Switch.scala 41:38:@32021.4]
  assign _T_70864 = select_32 == 6'h2c; // @[Switch.scala 41:52:@32023.4]
  assign output_44_32 = io_outValid_32 & _T_70864; // @[Switch.scala 41:38:@32024.4]
  assign _T_70867 = select_33 == 6'h2c; // @[Switch.scala 41:52:@32026.4]
  assign output_44_33 = io_outValid_33 & _T_70867; // @[Switch.scala 41:38:@32027.4]
  assign _T_70870 = select_34 == 6'h2c; // @[Switch.scala 41:52:@32029.4]
  assign output_44_34 = io_outValid_34 & _T_70870; // @[Switch.scala 41:38:@32030.4]
  assign _T_70873 = select_35 == 6'h2c; // @[Switch.scala 41:52:@32032.4]
  assign output_44_35 = io_outValid_35 & _T_70873; // @[Switch.scala 41:38:@32033.4]
  assign _T_70876 = select_36 == 6'h2c; // @[Switch.scala 41:52:@32035.4]
  assign output_44_36 = io_outValid_36 & _T_70876; // @[Switch.scala 41:38:@32036.4]
  assign _T_70879 = select_37 == 6'h2c; // @[Switch.scala 41:52:@32038.4]
  assign output_44_37 = io_outValid_37 & _T_70879; // @[Switch.scala 41:38:@32039.4]
  assign _T_70882 = select_38 == 6'h2c; // @[Switch.scala 41:52:@32041.4]
  assign output_44_38 = io_outValid_38 & _T_70882; // @[Switch.scala 41:38:@32042.4]
  assign _T_70885 = select_39 == 6'h2c; // @[Switch.scala 41:52:@32044.4]
  assign output_44_39 = io_outValid_39 & _T_70885; // @[Switch.scala 41:38:@32045.4]
  assign _T_70888 = select_40 == 6'h2c; // @[Switch.scala 41:52:@32047.4]
  assign output_44_40 = io_outValid_40 & _T_70888; // @[Switch.scala 41:38:@32048.4]
  assign _T_70891 = select_41 == 6'h2c; // @[Switch.scala 41:52:@32050.4]
  assign output_44_41 = io_outValid_41 & _T_70891; // @[Switch.scala 41:38:@32051.4]
  assign _T_70894 = select_42 == 6'h2c; // @[Switch.scala 41:52:@32053.4]
  assign output_44_42 = io_outValid_42 & _T_70894; // @[Switch.scala 41:38:@32054.4]
  assign _T_70897 = select_43 == 6'h2c; // @[Switch.scala 41:52:@32056.4]
  assign output_44_43 = io_outValid_43 & _T_70897; // @[Switch.scala 41:38:@32057.4]
  assign _T_70900 = select_44 == 6'h2c; // @[Switch.scala 41:52:@32059.4]
  assign output_44_44 = io_outValid_44 & _T_70900; // @[Switch.scala 41:38:@32060.4]
  assign _T_70903 = select_45 == 6'h2c; // @[Switch.scala 41:52:@32062.4]
  assign output_44_45 = io_outValid_45 & _T_70903; // @[Switch.scala 41:38:@32063.4]
  assign _T_70906 = select_46 == 6'h2c; // @[Switch.scala 41:52:@32065.4]
  assign output_44_46 = io_outValid_46 & _T_70906; // @[Switch.scala 41:38:@32066.4]
  assign _T_70909 = select_47 == 6'h2c; // @[Switch.scala 41:52:@32068.4]
  assign output_44_47 = io_outValid_47 & _T_70909; // @[Switch.scala 41:38:@32069.4]
  assign _T_70912 = select_48 == 6'h2c; // @[Switch.scala 41:52:@32071.4]
  assign output_44_48 = io_outValid_48 & _T_70912; // @[Switch.scala 41:38:@32072.4]
  assign _T_70915 = select_49 == 6'h2c; // @[Switch.scala 41:52:@32074.4]
  assign output_44_49 = io_outValid_49 & _T_70915; // @[Switch.scala 41:38:@32075.4]
  assign _T_70918 = select_50 == 6'h2c; // @[Switch.scala 41:52:@32077.4]
  assign output_44_50 = io_outValid_50 & _T_70918; // @[Switch.scala 41:38:@32078.4]
  assign _T_70921 = select_51 == 6'h2c; // @[Switch.scala 41:52:@32080.4]
  assign output_44_51 = io_outValid_51 & _T_70921; // @[Switch.scala 41:38:@32081.4]
  assign _T_70924 = select_52 == 6'h2c; // @[Switch.scala 41:52:@32083.4]
  assign output_44_52 = io_outValid_52 & _T_70924; // @[Switch.scala 41:38:@32084.4]
  assign _T_70927 = select_53 == 6'h2c; // @[Switch.scala 41:52:@32086.4]
  assign output_44_53 = io_outValid_53 & _T_70927; // @[Switch.scala 41:38:@32087.4]
  assign _T_70930 = select_54 == 6'h2c; // @[Switch.scala 41:52:@32089.4]
  assign output_44_54 = io_outValid_54 & _T_70930; // @[Switch.scala 41:38:@32090.4]
  assign _T_70933 = select_55 == 6'h2c; // @[Switch.scala 41:52:@32092.4]
  assign output_44_55 = io_outValid_55 & _T_70933; // @[Switch.scala 41:38:@32093.4]
  assign _T_70936 = select_56 == 6'h2c; // @[Switch.scala 41:52:@32095.4]
  assign output_44_56 = io_outValid_56 & _T_70936; // @[Switch.scala 41:38:@32096.4]
  assign _T_70939 = select_57 == 6'h2c; // @[Switch.scala 41:52:@32098.4]
  assign output_44_57 = io_outValid_57 & _T_70939; // @[Switch.scala 41:38:@32099.4]
  assign _T_70942 = select_58 == 6'h2c; // @[Switch.scala 41:52:@32101.4]
  assign output_44_58 = io_outValid_58 & _T_70942; // @[Switch.scala 41:38:@32102.4]
  assign _T_70945 = select_59 == 6'h2c; // @[Switch.scala 41:52:@32104.4]
  assign output_44_59 = io_outValid_59 & _T_70945; // @[Switch.scala 41:38:@32105.4]
  assign _T_70948 = select_60 == 6'h2c; // @[Switch.scala 41:52:@32107.4]
  assign output_44_60 = io_outValid_60 & _T_70948; // @[Switch.scala 41:38:@32108.4]
  assign _T_70951 = select_61 == 6'h2c; // @[Switch.scala 41:52:@32110.4]
  assign output_44_61 = io_outValid_61 & _T_70951; // @[Switch.scala 41:38:@32111.4]
  assign _T_70954 = select_62 == 6'h2c; // @[Switch.scala 41:52:@32113.4]
  assign output_44_62 = io_outValid_62 & _T_70954; // @[Switch.scala 41:38:@32114.4]
  assign _T_70957 = select_63 == 6'h2c; // @[Switch.scala 41:52:@32116.4]
  assign output_44_63 = io_outValid_63 & _T_70957; // @[Switch.scala 41:38:@32117.4]
  assign _T_70965 = {output_44_7,output_44_6,output_44_5,output_44_4,output_44_3,output_44_2,output_44_1,output_44_0}; // @[Switch.scala 43:31:@32125.4]
  assign _T_70973 = {output_44_15,output_44_14,output_44_13,output_44_12,output_44_11,output_44_10,output_44_9,output_44_8,_T_70965}; // @[Switch.scala 43:31:@32133.4]
  assign _T_70980 = {output_44_23,output_44_22,output_44_21,output_44_20,output_44_19,output_44_18,output_44_17,output_44_16}; // @[Switch.scala 43:31:@32140.4]
  assign _T_70989 = {output_44_31,output_44_30,output_44_29,output_44_28,output_44_27,output_44_26,output_44_25,output_44_24,_T_70980,_T_70973}; // @[Switch.scala 43:31:@32149.4]
  assign _T_70996 = {output_44_39,output_44_38,output_44_37,output_44_36,output_44_35,output_44_34,output_44_33,output_44_32}; // @[Switch.scala 43:31:@32156.4]
  assign _T_71004 = {output_44_47,output_44_46,output_44_45,output_44_44,output_44_43,output_44_42,output_44_41,output_44_40,_T_70996}; // @[Switch.scala 43:31:@32164.4]
  assign _T_71011 = {output_44_55,output_44_54,output_44_53,output_44_52,output_44_51,output_44_50,output_44_49,output_44_48}; // @[Switch.scala 43:31:@32171.4]
  assign _T_71020 = {output_44_63,output_44_62,output_44_61,output_44_60,output_44_59,output_44_58,output_44_57,output_44_56,_T_71011,_T_71004}; // @[Switch.scala 43:31:@32180.4]
  assign _T_71021 = {_T_71020,_T_70989}; // @[Switch.scala 43:31:@32181.4]
  assign _T_71025 = select_0 == 6'h2d; // @[Switch.scala 41:52:@32184.4]
  assign output_45_0 = io_outValid_0 & _T_71025; // @[Switch.scala 41:38:@32185.4]
  assign _T_71028 = select_1 == 6'h2d; // @[Switch.scala 41:52:@32187.4]
  assign output_45_1 = io_outValid_1 & _T_71028; // @[Switch.scala 41:38:@32188.4]
  assign _T_71031 = select_2 == 6'h2d; // @[Switch.scala 41:52:@32190.4]
  assign output_45_2 = io_outValid_2 & _T_71031; // @[Switch.scala 41:38:@32191.4]
  assign _T_71034 = select_3 == 6'h2d; // @[Switch.scala 41:52:@32193.4]
  assign output_45_3 = io_outValid_3 & _T_71034; // @[Switch.scala 41:38:@32194.4]
  assign _T_71037 = select_4 == 6'h2d; // @[Switch.scala 41:52:@32196.4]
  assign output_45_4 = io_outValid_4 & _T_71037; // @[Switch.scala 41:38:@32197.4]
  assign _T_71040 = select_5 == 6'h2d; // @[Switch.scala 41:52:@32199.4]
  assign output_45_5 = io_outValid_5 & _T_71040; // @[Switch.scala 41:38:@32200.4]
  assign _T_71043 = select_6 == 6'h2d; // @[Switch.scala 41:52:@32202.4]
  assign output_45_6 = io_outValid_6 & _T_71043; // @[Switch.scala 41:38:@32203.4]
  assign _T_71046 = select_7 == 6'h2d; // @[Switch.scala 41:52:@32205.4]
  assign output_45_7 = io_outValid_7 & _T_71046; // @[Switch.scala 41:38:@32206.4]
  assign _T_71049 = select_8 == 6'h2d; // @[Switch.scala 41:52:@32208.4]
  assign output_45_8 = io_outValid_8 & _T_71049; // @[Switch.scala 41:38:@32209.4]
  assign _T_71052 = select_9 == 6'h2d; // @[Switch.scala 41:52:@32211.4]
  assign output_45_9 = io_outValid_9 & _T_71052; // @[Switch.scala 41:38:@32212.4]
  assign _T_71055 = select_10 == 6'h2d; // @[Switch.scala 41:52:@32214.4]
  assign output_45_10 = io_outValid_10 & _T_71055; // @[Switch.scala 41:38:@32215.4]
  assign _T_71058 = select_11 == 6'h2d; // @[Switch.scala 41:52:@32217.4]
  assign output_45_11 = io_outValid_11 & _T_71058; // @[Switch.scala 41:38:@32218.4]
  assign _T_71061 = select_12 == 6'h2d; // @[Switch.scala 41:52:@32220.4]
  assign output_45_12 = io_outValid_12 & _T_71061; // @[Switch.scala 41:38:@32221.4]
  assign _T_71064 = select_13 == 6'h2d; // @[Switch.scala 41:52:@32223.4]
  assign output_45_13 = io_outValid_13 & _T_71064; // @[Switch.scala 41:38:@32224.4]
  assign _T_71067 = select_14 == 6'h2d; // @[Switch.scala 41:52:@32226.4]
  assign output_45_14 = io_outValid_14 & _T_71067; // @[Switch.scala 41:38:@32227.4]
  assign _T_71070 = select_15 == 6'h2d; // @[Switch.scala 41:52:@32229.4]
  assign output_45_15 = io_outValid_15 & _T_71070; // @[Switch.scala 41:38:@32230.4]
  assign _T_71073 = select_16 == 6'h2d; // @[Switch.scala 41:52:@32232.4]
  assign output_45_16 = io_outValid_16 & _T_71073; // @[Switch.scala 41:38:@32233.4]
  assign _T_71076 = select_17 == 6'h2d; // @[Switch.scala 41:52:@32235.4]
  assign output_45_17 = io_outValid_17 & _T_71076; // @[Switch.scala 41:38:@32236.4]
  assign _T_71079 = select_18 == 6'h2d; // @[Switch.scala 41:52:@32238.4]
  assign output_45_18 = io_outValid_18 & _T_71079; // @[Switch.scala 41:38:@32239.4]
  assign _T_71082 = select_19 == 6'h2d; // @[Switch.scala 41:52:@32241.4]
  assign output_45_19 = io_outValid_19 & _T_71082; // @[Switch.scala 41:38:@32242.4]
  assign _T_71085 = select_20 == 6'h2d; // @[Switch.scala 41:52:@32244.4]
  assign output_45_20 = io_outValid_20 & _T_71085; // @[Switch.scala 41:38:@32245.4]
  assign _T_71088 = select_21 == 6'h2d; // @[Switch.scala 41:52:@32247.4]
  assign output_45_21 = io_outValid_21 & _T_71088; // @[Switch.scala 41:38:@32248.4]
  assign _T_71091 = select_22 == 6'h2d; // @[Switch.scala 41:52:@32250.4]
  assign output_45_22 = io_outValid_22 & _T_71091; // @[Switch.scala 41:38:@32251.4]
  assign _T_71094 = select_23 == 6'h2d; // @[Switch.scala 41:52:@32253.4]
  assign output_45_23 = io_outValid_23 & _T_71094; // @[Switch.scala 41:38:@32254.4]
  assign _T_71097 = select_24 == 6'h2d; // @[Switch.scala 41:52:@32256.4]
  assign output_45_24 = io_outValid_24 & _T_71097; // @[Switch.scala 41:38:@32257.4]
  assign _T_71100 = select_25 == 6'h2d; // @[Switch.scala 41:52:@32259.4]
  assign output_45_25 = io_outValid_25 & _T_71100; // @[Switch.scala 41:38:@32260.4]
  assign _T_71103 = select_26 == 6'h2d; // @[Switch.scala 41:52:@32262.4]
  assign output_45_26 = io_outValid_26 & _T_71103; // @[Switch.scala 41:38:@32263.4]
  assign _T_71106 = select_27 == 6'h2d; // @[Switch.scala 41:52:@32265.4]
  assign output_45_27 = io_outValid_27 & _T_71106; // @[Switch.scala 41:38:@32266.4]
  assign _T_71109 = select_28 == 6'h2d; // @[Switch.scala 41:52:@32268.4]
  assign output_45_28 = io_outValid_28 & _T_71109; // @[Switch.scala 41:38:@32269.4]
  assign _T_71112 = select_29 == 6'h2d; // @[Switch.scala 41:52:@32271.4]
  assign output_45_29 = io_outValid_29 & _T_71112; // @[Switch.scala 41:38:@32272.4]
  assign _T_71115 = select_30 == 6'h2d; // @[Switch.scala 41:52:@32274.4]
  assign output_45_30 = io_outValid_30 & _T_71115; // @[Switch.scala 41:38:@32275.4]
  assign _T_71118 = select_31 == 6'h2d; // @[Switch.scala 41:52:@32277.4]
  assign output_45_31 = io_outValid_31 & _T_71118; // @[Switch.scala 41:38:@32278.4]
  assign _T_71121 = select_32 == 6'h2d; // @[Switch.scala 41:52:@32280.4]
  assign output_45_32 = io_outValid_32 & _T_71121; // @[Switch.scala 41:38:@32281.4]
  assign _T_71124 = select_33 == 6'h2d; // @[Switch.scala 41:52:@32283.4]
  assign output_45_33 = io_outValid_33 & _T_71124; // @[Switch.scala 41:38:@32284.4]
  assign _T_71127 = select_34 == 6'h2d; // @[Switch.scala 41:52:@32286.4]
  assign output_45_34 = io_outValid_34 & _T_71127; // @[Switch.scala 41:38:@32287.4]
  assign _T_71130 = select_35 == 6'h2d; // @[Switch.scala 41:52:@32289.4]
  assign output_45_35 = io_outValid_35 & _T_71130; // @[Switch.scala 41:38:@32290.4]
  assign _T_71133 = select_36 == 6'h2d; // @[Switch.scala 41:52:@32292.4]
  assign output_45_36 = io_outValid_36 & _T_71133; // @[Switch.scala 41:38:@32293.4]
  assign _T_71136 = select_37 == 6'h2d; // @[Switch.scala 41:52:@32295.4]
  assign output_45_37 = io_outValid_37 & _T_71136; // @[Switch.scala 41:38:@32296.4]
  assign _T_71139 = select_38 == 6'h2d; // @[Switch.scala 41:52:@32298.4]
  assign output_45_38 = io_outValid_38 & _T_71139; // @[Switch.scala 41:38:@32299.4]
  assign _T_71142 = select_39 == 6'h2d; // @[Switch.scala 41:52:@32301.4]
  assign output_45_39 = io_outValid_39 & _T_71142; // @[Switch.scala 41:38:@32302.4]
  assign _T_71145 = select_40 == 6'h2d; // @[Switch.scala 41:52:@32304.4]
  assign output_45_40 = io_outValid_40 & _T_71145; // @[Switch.scala 41:38:@32305.4]
  assign _T_71148 = select_41 == 6'h2d; // @[Switch.scala 41:52:@32307.4]
  assign output_45_41 = io_outValid_41 & _T_71148; // @[Switch.scala 41:38:@32308.4]
  assign _T_71151 = select_42 == 6'h2d; // @[Switch.scala 41:52:@32310.4]
  assign output_45_42 = io_outValid_42 & _T_71151; // @[Switch.scala 41:38:@32311.4]
  assign _T_71154 = select_43 == 6'h2d; // @[Switch.scala 41:52:@32313.4]
  assign output_45_43 = io_outValid_43 & _T_71154; // @[Switch.scala 41:38:@32314.4]
  assign _T_71157 = select_44 == 6'h2d; // @[Switch.scala 41:52:@32316.4]
  assign output_45_44 = io_outValid_44 & _T_71157; // @[Switch.scala 41:38:@32317.4]
  assign _T_71160 = select_45 == 6'h2d; // @[Switch.scala 41:52:@32319.4]
  assign output_45_45 = io_outValid_45 & _T_71160; // @[Switch.scala 41:38:@32320.4]
  assign _T_71163 = select_46 == 6'h2d; // @[Switch.scala 41:52:@32322.4]
  assign output_45_46 = io_outValid_46 & _T_71163; // @[Switch.scala 41:38:@32323.4]
  assign _T_71166 = select_47 == 6'h2d; // @[Switch.scala 41:52:@32325.4]
  assign output_45_47 = io_outValid_47 & _T_71166; // @[Switch.scala 41:38:@32326.4]
  assign _T_71169 = select_48 == 6'h2d; // @[Switch.scala 41:52:@32328.4]
  assign output_45_48 = io_outValid_48 & _T_71169; // @[Switch.scala 41:38:@32329.4]
  assign _T_71172 = select_49 == 6'h2d; // @[Switch.scala 41:52:@32331.4]
  assign output_45_49 = io_outValid_49 & _T_71172; // @[Switch.scala 41:38:@32332.4]
  assign _T_71175 = select_50 == 6'h2d; // @[Switch.scala 41:52:@32334.4]
  assign output_45_50 = io_outValid_50 & _T_71175; // @[Switch.scala 41:38:@32335.4]
  assign _T_71178 = select_51 == 6'h2d; // @[Switch.scala 41:52:@32337.4]
  assign output_45_51 = io_outValid_51 & _T_71178; // @[Switch.scala 41:38:@32338.4]
  assign _T_71181 = select_52 == 6'h2d; // @[Switch.scala 41:52:@32340.4]
  assign output_45_52 = io_outValid_52 & _T_71181; // @[Switch.scala 41:38:@32341.4]
  assign _T_71184 = select_53 == 6'h2d; // @[Switch.scala 41:52:@32343.4]
  assign output_45_53 = io_outValid_53 & _T_71184; // @[Switch.scala 41:38:@32344.4]
  assign _T_71187 = select_54 == 6'h2d; // @[Switch.scala 41:52:@32346.4]
  assign output_45_54 = io_outValid_54 & _T_71187; // @[Switch.scala 41:38:@32347.4]
  assign _T_71190 = select_55 == 6'h2d; // @[Switch.scala 41:52:@32349.4]
  assign output_45_55 = io_outValid_55 & _T_71190; // @[Switch.scala 41:38:@32350.4]
  assign _T_71193 = select_56 == 6'h2d; // @[Switch.scala 41:52:@32352.4]
  assign output_45_56 = io_outValid_56 & _T_71193; // @[Switch.scala 41:38:@32353.4]
  assign _T_71196 = select_57 == 6'h2d; // @[Switch.scala 41:52:@32355.4]
  assign output_45_57 = io_outValid_57 & _T_71196; // @[Switch.scala 41:38:@32356.4]
  assign _T_71199 = select_58 == 6'h2d; // @[Switch.scala 41:52:@32358.4]
  assign output_45_58 = io_outValid_58 & _T_71199; // @[Switch.scala 41:38:@32359.4]
  assign _T_71202 = select_59 == 6'h2d; // @[Switch.scala 41:52:@32361.4]
  assign output_45_59 = io_outValid_59 & _T_71202; // @[Switch.scala 41:38:@32362.4]
  assign _T_71205 = select_60 == 6'h2d; // @[Switch.scala 41:52:@32364.4]
  assign output_45_60 = io_outValid_60 & _T_71205; // @[Switch.scala 41:38:@32365.4]
  assign _T_71208 = select_61 == 6'h2d; // @[Switch.scala 41:52:@32367.4]
  assign output_45_61 = io_outValid_61 & _T_71208; // @[Switch.scala 41:38:@32368.4]
  assign _T_71211 = select_62 == 6'h2d; // @[Switch.scala 41:52:@32370.4]
  assign output_45_62 = io_outValid_62 & _T_71211; // @[Switch.scala 41:38:@32371.4]
  assign _T_71214 = select_63 == 6'h2d; // @[Switch.scala 41:52:@32373.4]
  assign output_45_63 = io_outValid_63 & _T_71214; // @[Switch.scala 41:38:@32374.4]
  assign _T_71222 = {output_45_7,output_45_6,output_45_5,output_45_4,output_45_3,output_45_2,output_45_1,output_45_0}; // @[Switch.scala 43:31:@32382.4]
  assign _T_71230 = {output_45_15,output_45_14,output_45_13,output_45_12,output_45_11,output_45_10,output_45_9,output_45_8,_T_71222}; // @[Switch.scala 43:31:@32390.4]
  assign _T_71237 = {output_45_23,output_45_22,output_45_21,output_45_20,output_45_19,output_45_18,output_45_17,output_45_16}; // @[Switch.scala 43:31:@32397.4]
  assign _T_71246 = {output_45_31,output_45_30,output_45_29,output_45_28,output_45_27,output_45_26,output_45_25,output_45_24,_T_71237,_T_71230}; // @[Switch.scala 43:31:@32406.4]
  assign _T_71253 = {output_45_39,output_45_38,output_45_37,output_45_36,output_45_35,output_45_34,output_45_33,output_45_32}; // @[Switch.scala 43:31:@32413.4]
  assign _T_71261 = {output_45_47,output_45_46,output_45_45,output_45_44,output_45_43,output_45_42,output_45_41,output_45_40,_T_71253}; // @[Switch.scala 43:31:@32421.4]
  assign _T_71268 = {output_45_55,output_45_54,output_45_53,output_45_52,output_45_51,output_45_50,output_45_49,output_45_48}; // @[Switch.scala 43:31:@32428.4]
  assign _T_71277 = {output_45_63,output_45_62,output_45_61,output_45_60,output_45_59,output_45_58,output_45_57,output_45_56,_T_71268,_T_71261}; // @[Switch.scala 43:31:@32437.4]
  assign _T_71278 = {_T_71277,_T_71246}; // @[Switch.scala 43:31:@32438.4]
  assign _T_71282 = select_0 == 6'h2e; // @[Switch.scala 41:52:@32441.4]
  assign output_46_0 = io_outValid_0 & _T_71282; // @[Switch.scala 41:38:@32442.4]
  assign _T_71285 = select_1 == 6'h2e; // @[Switch.scala 41:52:@32444.4]
  assign output_46_1 = io_outValid_1 & _T_71285; // @[Switch.scala 41:38:@32445.4]
  assign _T_71288 = select_2 == 6'h2e; // @[Switch.scala 41:52:@32447.4]
  assign output_46_2 = io_outValid_2 & _T_71288; // @[Switch.scala 41:38:@32448.4]
  assign _T_71291 = select_3 == 6'h2e; // @[Switch.scala 41:52:@32450.4]
  assign output_46_3 = io_outValid_3 & _T_71291; // @[Switch.scala 41:38:@32451.4]
  assign _T_71294 = select_4 == 6'h2e; // @[Switch.scala 41:52:@32453.4]
  assign output_46_4 = io_outValid_4 & _T_71294; // @[Switch.scala 41:38:@32454.4]
  assign _T_71297 = select_5 == 6'h2e; // @[Switch.scala 41:52:@32456.4]
  assign output_46_5 = io_outValid_5 & _T_71297; // @[Switch.scala 41:38:@32457.4]
  assign _T_71300 = select_6 == 6'h2e; // @[Switch.scala 41:52:@32459.4]
  assign output_46_6 = io_outValid_6 & _T_71300; // @[Switch.scala 41:38:@32460.4]
  assign _T_71303 = select_7 == 6'h2e; // @[Switch.scala 41:52:@32462.4]
  assign output_46_7 = io_outValid_7 & _T_71303; // @[Switch.scala 41:38:@32463.4]
  assign _T_71306 = select_8 == 6'h2e; // @[Switch.scala 41:52:@32465.4]
  assign output_46_8 = io_outValid_8 & _T_71306; // @[Switch.scala 41:38:@32466.4]
  assign _T_71309 = select_9 == 6'h2e; // @[Switch.scala 41:52:@32468.4]
  assign output_46_9 = io_outValid_9 & _T_71309; // @[Switch.scala 41:38:@32469.4]
  assign _T_71312 = select_10 == 6'h2e; // @[Switch.scala 41:52:@32471.4]
  assign output_46_10 = io_outValid_10 & _T_71312; // @[Switch.scala 41:38:@32472.4]
  assign _T_71315 = select_11 == 6'h2e; // @[Switch.scala 41:52:@32474.4]
  assign output_46_11 = io_outValid_11 & _T_71315; // @[Switch.scala 41:38:@32475.4]
  assign _T_71318 = select_12 == 6'h2e; // @[Switch.scala 41:52:@32477.4]
  assign output_46_12 = io_outValid_12 & _T_71318; // @[Switch.scala 41:38:@32478.4]
  assign _T_71321 = select_13 == 6'h2e; // @[Switch.scala 41:52:@32480.4]
  assign output_46_13 = io_outValid_13 & _T_71321; // @[Switch.scala 41:38:@32481.4]
  assign _T_71324 = select_14 == 6'h2e; // @[Switch.scala 41:52:@32483.4]
  assign output_46_14 = io_outValid_14 & _T_71324; // @[Switch.scala 41:38:@32484.4]
  assign _T_71327 = select_15 == 6'h2e; // @[Switch.scala 41:52:@32486.4]
  assign output_46_15 = io_outValid_15 & _T_71327; // @[Switch.scala 41:38:@32487.4]
  assign _T_71330 = select_16 == 6'h2e; // @[Switch.scala 41:52:@32489.4]
  assign output_46_16 = io_outValid_16 & _T_71330; // @[Switch.scala 41:38:@32490.4]
  assign _T_71333 = select_17 == 6'h2e; // @[Switch.scala 41:52:@32492.4]
  assign output_46_17 = io_outValid_17 & _T_71333; // @[Switch.scala 41:38:@32493.4]
  assign _T_71336 = select_18 == 6'h2e; // @[Switch.scala 41:52:@32495.4]
  assign output_46_18 = io_outValid_18 & _T_71336; // @[Switch.scala 41:38:@32496.4]
  assign _T_71339 = select_19 == 6'h2e; // @[Switch.scala 41:52:@32498.4]
  assign output_46_19 = io_outValid_19 & _T_71339; // @[Switch.scala 41:38:@32499.4]
  assign _T_71342 = select_20 == 6'h2e; // @[Switch.scala 41:52:@32501.4]
  assign output_46_20 = io_outValid_20 & _T_71342; // @[Switch.scala 41:38:@32502.4]
  assign _T_71345 = select_21 == 6'h2e; // @[Switch.scala 41:52:@32504.4]
  assign output_46_21 = io_outValid_21 & _T_71345; // @[Switch.scala 41:38:@32505.4]
  assign _T_71348 = select_22 == 6'h2e; // @[Switch.scala 41:52:@32507.4]
  assign output_46_22 = io_outValid_22 & _T_71348; // @[Switch.scala 41:38:@32508.4]
  assign _T_71351 = select_23 == 6'h2e; // @[Switch.scala 41:52:@32510.4]
  assign output_46_23 = io_outValid_23 & _T_71351; // @[Switch.scala 41:38:@32511.4]
  assign _T_71354 = select_24 == 6'h2e; // @[Switch.scala 41:52:@32513.4]
  assign output_46_24 = io_outValid_24 & _T_71354; // @[Switch.scala 41:38:@32514.4]
  assign _T_71357 = select_25 == 6'h2e; // @[Switch.scala 41:52:@32516.4]
  assign output_46_25 = io_outValid_25 & _T_71357; // @[Switch.scala 41:38:@32517.4]
  assign _T_71360 = select_26 == 6'h2e; // @[Switch.scala 41:52:@32519.4]
  assign output_46_26 = io_outValid_26 & _T_71360; // @[Switch.scala 41:38:@32520.4]
  assign _T_71363 = select_27 == 6'h2e; // @[Switch.scala 41:52:@32522.4]
  assign output_46_27 = io_outValid_27 & _T_71363; // @[Switch.scala 41:38:@32523.4]
  assign _T_71366 = select_28 == 6'h2e; // @[Switch.scala 41:52:@32525.4]
  assign output_46_28 = io_outValid_28 & _T_71366; // @[Switch.scala 41:38:@32526.4]
  assign _T_71369 = select_29 == 6'h2e; // @[Switch.scala 41:52:@32528.4]
  assign output_46_29 = io_outValid_29 & _T_71369; // @[Switch.scala 41:38:@32529.4]
  assign _T_71372 = select_30 == 6'h2e; // @[Switch.scala 41:52:@32531.4]
  assign output_46_30 = io_outValid_30 & _T_71372; // @[Switch.scala 41:38:@32532.4]
  assign _T_71375 = select_31 == 6'h2e; // @[Switch.scala 41:52:@32534.4]
  assign output_46_31 = io_outValid_31 & _T_71375; // @[Switch.scala 41:38:@32535.4]
  assign _T_71378 = select_32 == 6'h2e; // @[Switch.scala 41:52:@32537.4]
  assign output_46_32 = io_outValid_32 & _T_71378; // @[Switch.scala 41:38:@32538.4]
  assign _T_71381 = select_33 == 6'h2e; // @[Switch.scala 41:52:@32540.4]
  assign output_46_33 = io_outValid_33 & _T_71381; // @[Switch.scala 41:38:@32541.4]
  assign _T_71384 = select_34 == 6'h2e; // @[Switch.scala 41:52:@32543.4]
  assign output_46_34 = io_outValid_34 & _T_71384; // @[Switch.scala 41:38:@32544.4]
  assign _T_71387 = select_35 == 6'h2e; // @[Switch.scala 41:52:@32546.4]
  assign output_46_35 = io_outValid_35 & _T_71387; // @[Switch.scala 41:38:@32547.4]
  assign _T_71390 = select_36 == 6'h2e; // @[Switch.scala 41:52:@32549.4]
  assign output_46_36 = io_outValid_36 & _T_71390; // @[Switch.scala 41:38:@32550.4]
  assign _T_71393 = select_37 == 6'h2e; // @[Switch.scala 41:52:@32552.4]
  assign output_46_37 = io_outValid_37 & _T_71393; // @[Switch.scala 41:38:@32553.4]
  assign _T_71396 = select_38 == 6'h2e; // @[Switch.scala 41:52:@32555.4]
  assign output_46_38 = io_outValid_38 & _T_71396; // @[Switch.scala 41:38:@32556.4]
  assign _T_71399 = select_39 == 6'h2e; // @[Switch.scala 41:52:@32558.4]
  assign output_46_39 = io_outValid_39 & _T_71399; // @[Switch.scala 41:38:@32559.4]
  assign _T_71402 = select_40 == 6'h2e; // @[Switch.scala 41:52:@32561.4]
  assign output_46_40 = io_outValid_40 & _T_71402; // @[Switch.scala 41:38:@32562.4]
  assign _T_71405 = select_41 == 6'h2e; // @[Switch.scala 41:52:@32564.4]
  assign output_46_41 = io_outValid_41 & _T_71405; // @[Switch.scala 41:38:@32565.4]
  assign _T_71408 = select_42 == 6'h2e; // @[Switch.scala 41:52:@32567.4]
  assign output_46_42 = io_outValid_42 & _T_71408; // @[Switch.scala 41:38:@32568.4]
  assign _T_71411 = select_43 == 6'h2e; // @[Switch.scala 41:52:@32570.4]
  assign output_46_43 = io_outValid_43 & _T_71411; // @[Switch.scala 41:38:@32571.4]
  assign _T_71414 = select_44 == 6'h2e; // @[Switch.scala 41:52:@32573.4]
  assign output_46_44 = io_outValid_44 & _T_71414; // @[Switch.scala 41:38:@32574.4]
  assign _T_71417 = select_45 == 6'h2e; // @[Switch.scala 41:52:@32576.4]
  assign output_46_45 = io_outValid_45 & _T_71417; // @[Switch.scala 41:38:@32577.4]
  assign _T_71420 = select_46 == 6'h2e; // @[Switch.scala 41:52:@32579.4]
  assign output_46_46 = io_outValid_46 & _T_71420; // @[Switch.scala 41:38:@32580.4]
  assign _T_71423 = select_47 == 6'h2e; // @[Switch.scala 41:52:@32582.4]
  assign output_46_47 = io_outValid_47 & _T_71423; // @[Switch.scala 41:38:@32583.4]
  assign _T_71426 = select_48 == 6'h2e; // @[Switch.scala 41:52:@32585.4]
  assign output_46_48 = io_outValid_48 & _T_71426; // @[Switch.scala 41:38:@32586.4]
  assign _T_71429 = select_49 == 6'h2e; // @[Switch.scala 41:52:@32588.4]
  assign output_46_49 = io_outValid_49 & _T_71429; // @[Switch.scala 41:38:@32589.4]
  assign _T_71432 = select_50 == 6'h2e; // @[Switch.scala 41:52:@32591.4]
  assign output_46_50 = io_outValid_50 & _T_71432; // @[Switch.scala 41:38:@32592.4]
  assign _T_71435 = select_51 == 6'h2e; // @[Switch.scala 41:52:@32594.4]
  assign output_46_51 = io_outValid_51 & _T_71435; // @[Switch.scala 41:38:@32595.4]
  assign _T_71438 = select_52 == 6'h2e; // @[Switch.scala 41:52:@32597.4]
  assign output_46_52 = io_outValid_52 & _T_71438; // @[Switch.scala 41:38:@32598.4]
  assign _T_71441 = select_53 == 6'h2e; // @[Switch.scala 41:52:@32600.4]
  assign output_46_53 = io_outValid_53 & _T_71441; // @[Switch.scala 41:38:@32601.4]
  assign _T_71444 = select_54 == 6'h2e; // @[Switch.scala 41:52:@32603.4]
  assign output_46_54 = io_outValid_54 & _T_71444; // @[Switch.scala 41:38:@32604.4]
  assign _T_71447 = select_55 == 6'h2e; // @[Switch.scala 41:52:@32606.4]
  assign output_46_55 = io_outValid_55 & _T_71447; // @[Switch.scala 41:38:@32607.4]
  assign _T_71450 = select_56 == 6'h2e; // @[Switch.scala 41:52:@32609.4]
  assign output_46_56 = io_outValid_56 & _T_71450; // @[Switch.scala 41:38:@32610.4]
  assign _T_71453 = select_57 == 6'h2e; // @[Switch.scala 41:52:@32612.4]
  assign output_46_57 = io_outValid_57 & _T_71453; // @[Switch.scala 41:38:@32613.4]
  assign _T_71456 = select_58 == 6'h2e; // @[Switch.scala 41:52:@32615.4]
  assign output_46_58 = io_outValid_58 & _T_71456; // @[Switch.scala 41:38:@32616.4]
  assign _T_71459 = select_59 == 6'h2e; // @[Switch.scala 41:52:@32618.4]
  assign output_46_59 = io_outValid_59 & _T_71459; // @[Switch.scala 41:38:@32619.4]
  assign _T_71462 = select_60 == 6'h2e; // @[Switch.scala 41:52:@32621.4]
  assign output_46_60 = io_outValid_60 & _T_71462; // @[Switch.scala 41:38:@32622.4]
  assign _T_71465 = select_61 == 6'h2e; // @[Switch.scala 41:52:@32624.4]
  assign output_46_61 = io_outValid_61 & _T_71465; // @[Switch.scala 41:38:@32625.4]
  assign _T_71468 = select_62 == 6'h2e; // @[Switch.scala 41:52:@32627.4]
  assign output_46_62 = io_outValid_62 & _T_71468; // @[Switch.scala 41:38:@32628.4]
  assign _T_71471 = select_63 == 6'h2e; // @[Switch.scala 41:52:@32630.4]
  assign output_46_63 = io_outValid_63 & _T_71471; // @[Switch.scala 41:38:@32631.4]
  assign _T_71479 = {output_46_7,output_46_6,output_46_5,output_46_4,output_46_3,output_46_2,output_46_1,output_46_0}; // @[Switch.scala 43:31:@32639.4]
  assign _T_71487 = {output_46_15,output_46_14,output_46_13,output_46_12,output_46_11,output_46_10,output_46_9,output_46_8,_T_71479}; // @[Switch.scala 43:31:@32647.4]
  assign _T_71494 = {output_46_23,output_46_22,output_46_21,output_46_20,output_46_19,output_46_18,output_46_17,output_46_16}; // @[Switch.scala 43:31:@32654.4]
  assign _T_71503 = {output_46_31,output_46_30,output_46_29,output_46_28,output_46_27,output_46_26,output_46_25,output_46_24,_T_71494,_T_71487}; // @[Switch.scala 43:31:@32663.4]
  assign _T_71510 = {output_46_39,output_46_38,output_46_37,output_46_36,output_46_35,output_46_34,output_46_33,output_46_32}; // @[Switch.scala 43:31:@32670.4]
  assign _T_71518 = {output_46_47,output_46_46,output_46_45,output_46_44,output_46_43,output_46_42,output_46_41,output_46_40,_T_71510}; // @[Switch.scala 43:31:@32678.4]
  assign _T_71525 = {output_46_55,output_46_54,output_46_53,output_46_52,output_46_51,output_46_50,output_46_49,output_46_48}; // @[Switch.scala 43:31:@32685.4]
  assign _T_71534 = {output_46_63,output_46_62,output_46_61,output_46_60,output_46_59,output_46_58,output_46_57,output_46_56,_T_71525,_T_71518}; // @[Switch.scala 43:31:@32694.4]
  assign _T_71535 = {_T_71534,_T_71503}; // @[Switch.scala 43:31:@32695.4]
  assign _T_71539 = select_0 == 6'h2f; // @[Switch.scala 41:52:@32698.4]
  assign output_47_0 = io_outValid_0 & _T_71539; // @[Switch.scala 41:38:@32699.4]
  assign _T_71542 = select_1 == 6'h2f; // @[Switch.scala 41:52:@32701.4]
  assign output_47_1 = io_outValid_1 & _T_71542; // @[Switch.scala 41:38:@32702.4]
  assign _T_71545 = select_2 == 6'h2f; // @[Switch.scala 41:52:@32704.4]
  assign output_47_2 = io_outValid_2 & _T_71545; // @[Switch.scala 41:38:@32705.4]
  assign _T_71548 = select_3 == 6'h2f; // @[Switch.scala 41:52:@32707.4]
  assign output_47_3 = io_outValid_3 & _T_71548; // @[Switch.scala 41:38:@32708.4]
  assign _T_71551 = select_4 == 6'h2f; // @[Switch.scala 41:52:@32710.4]
  assign output_47_4 = io_outValid_4 & _T_71551; // @[Switch.scala 41:38:@32711.4]
  assign _T_71554 = select_5 == 6'h2f; // @[Switch.scala 41:52:@32713.4]
  assign output_47_5 = io_outValid_5 & _T_71554; // @[Switch.scala 41:38:@32714.4]
  assign _T_71557 = select_6 == 6'h2f; // @[Switch.scala 41:52:@32716.4]
  assign output_47_6 = io_outValid_6 & _T_71557; // @[Switch.scala 41:38:@32717.4]
  assign _T_71560 = select_7 == 6'h2f; // @[Switch.scala 41:52:@32719.4]
  assign output_47_7 = io_outValid_7 & _T_71560; // @[Switch.scala 41:38:@32720.4]
  assign _T_71563 = select_8 == 6'h2f; // @[Switch.scala 41:52:@32722.4]
  assign output_47_8 = io_outValid_8 & _T_71563; // @[Switch.scala 41:38:@32723.4]
  assign _T_71566 = select_9 == 6'h2f; // @[Switch.scala 41:52:@32725.4]
  assign output_47_9 = io_outValid_9 & _T_71566; // @[Switch.scala 41:38:@32726.4]
  assign _T_71569 = select_10 == 6'h2f; // @[Switch.scala 41:52:@32728.4]
  assign output_47_10 = io_outValid_10 & _T_71569; // @[Switch.scala 41:38:@32729.4]
  assign _T_71572 = select_11 == 6'h2f; // @[Switch.scala 41:52:@32731.4]
  assign output_47_11 = io_outValid_11 & _T_71572; // @[Switch.scala 41:38:@32732.4]
  assign _T_71575 = select_12 == 6'h2f; // @[Switch.scala 41:52:@32734.4]
  assign output_47_12 = io_outValid_12 & _T_71575; // @[Switch.scala 41:38:@32735.4]
  assign _T_71578 = select_13 == 6'h2f; // @[Switch.scala 41:52:@32737.4]
  assign output_47_13 = io_outValid_13 & _T_71578; // @[Switch.scala 41:38:@32738.4]
  assign _T_71581 = select_14 == 6'h2f; // @[Switch.scala 41:52:@32740.4]
  assign output_47_14 = io_outValid_14 & _T_71581; // @[Switch.scala 41:38:@32741.4]
  assign _T_71584 = select_15 == 6'h2f; // @[Switch.scala 41:52:@32743.4]
  assign output_47_15 = io_outValid_15 & _T_71584; // @[Switch.scala 41:38:@32744.4]
  assign _T_71587 = select_16 == 6'h2f; // @[Switch.scala 41:52:@32746.4]
  assign output_47_16 = io_outValid_16 & _T_71587; // @[Switch.scala 41:38:@32747.4]
  assign _T_71590 = select_17 == 6'h2f; // @[Switch.scala 41:52:@32749.4]
  assign output_47_17 = io_outValid_17 & _T_71590; // @[Switch.scala 41:38:@32750.4]
  assign _T_71593 = select_18 == 6'h2f; // @[Switch.scala 41:52:@32752.4]
  assign output_47_18 = io_outValid_18 & _T_71593; // @[Switch.scala 41:38:@32753.4]
  assign _T_71596 = select_19 == 6'h2f; // @[Switch.scala 41:52:@32755.4]
  assign output_47_19 = io_outValid_19 & _T_71596; // @[Switch.scala 41:38:@32756.4]
  assign _T_71599 = select_20 == 6'h2f; // @[Switch.scala 41:52:@32758.4]
  assign output_47_20 = io_outValid_20 & _T_71599; // @[Switch.scala 41:38:@32759.4]
  assign _T_71602 = select_21 == 6'h2f; // @[Switch.scala 41:52:@32761.4]
  assign output_47_21 = io_outValid_21 & _T_71602; // @[Switch.scala 41:38:@32762.4]
  assign _T_71605 = select_22 == 6'h2f; // @[Switch.scala 41:52:@32764.4]
  assign output_47_22 = io_outValid_22 & _T_71605; // @[Switch.scala 41:38:@32765.4]
  assign _T_71608 = select_23 == 6'h2f; // @[Switch.scala 41:52:@32767.4]
  assign output_47_23 = io_outValid_23 & _T_71608; // @[Switch.scala 41:38:@32768.4]
  assign _T_71611 = select_24 == 6'h2f; // @[Switch.scala 41:52:@32770.4]
  assign output_47_24 = io_outValid_24 & _T_71611; // @[Switch.scala 41:38:@32771.4]
  assign _T_71614 = select_25 == 6'h2f; // @[Switch.scala 41:52:@32773.4]
  assign output_47_25 = io_outValid_25 & _T_71614; // @[Switch.scala 41:38:@32774.4]
  assign _T_71617 = select_26 == 6'h2f; // @[Switch.scala 41:52:@32776.4]
  assign output_47_26 = io_outValid_26 & _T_71617; // @[Switch.scala 41:38:@32777.4]
  assign _T_71620 = select_27 == 6'h2f; // @[Switch.scala 41:52:@32779.4]
  assign output_47_27 = io_outValid_27 & _T_71620; // @[Switch.scala 41:38:@32780.4]
  assign _T_71623 = select_28 == 6'h2f; // @[Switch.scala 41:52:@32782.4]
  assign output_47_28 = io_outValid_28 & _T_71623; // @[Switch.scala 41:38:@32783.4]
  assign _T_71626 = select_29 == 6'h2f; // @[Switch.scala 41:52:@32785.4]
  assign output_47_29 = io_outValid_29 & _T_71626; // @[Switch.scala 41:38:@32786.4]
  assign _T_71629 = select_30 == 6'h2f; // @[Switch.scala 41:52:@32788.4]
  assign output_47_30 = io_outValid_30 & _T_71629; // @[Switch.scala 41:38:@32789.4]
  assign _T_71632 = select_31 == 6'h2f; // @[Switch.scala 41:52:@32791.4]
  assign output_47_31 = io_outValid_31 & _T_71632; // @[Switch.scala 41:38:@32792.4]
  assign _T_71635 = select_32 == 6'h2f; // @[Switch.scala 41:52:@32794.4]
  assign output_47_32 = io_outValid_32 & _T_71635; // @[Switch.scala 41:38:@32795.4]
  assign _T_71638 = select_33 == 6'h2f; // @[Switch.scala 41:52:@32797.4]
  assign output_47_33 = io_outValid_33 & _T_71638; // @[Switch.scala 41:38:@32798.4]
  assign _T_71641 = select_34 == 6'h2f; // @[Switch.scala 41:52:@32800.4]
  assign output_47_34 = io_outValid_34 & _T_71641; // @[Switch.scala 41:38:@32801.4]
  assign _T_71644 = select_35 == 6'h2f; // @[Switch.scala 41:52:@32803.4]
  assign output_47_35 = io_outValid_35 & _T_71644; // @[Switch.scala 41:38:@32804.4]
  assign _T_71647 = select_36 == 6'h2f; // @[Switch.scala 41:52:@32806.4]
  assign output_47_36 = io_outValid_36 & _T_71647; // @[Switch.scala 41:38:@32807.4]
  assign _T_71650 = select_37 == 6'h2f; // @[Switch.scala 41:52:@32809.4]
  assign output_47_37 = io_outValid_37 & _T_71650; // @[Switch.scala 41:38:@32810.4]
  assign _T_71653 = select_38 == 6'h2f; // @[Switch.scala 41:52:@32812.4]
  assign output_47_38 = io_outValid_38 & _T_71653; // @[Switch.scala 41:38:@32813.4]
  assign _T_71656 = select_39 == 6'h2f; // @[Switch.scala 41:52:@32815.4]
  assign output_47_39 = io_outValid_39 & _T_71656; // @[Switch.scala 41:38:@32816.4]
  assign _T_71659 = select_40 == 6'h2f; // @[Switch.scala 41:52:@32818.4]
  assign output_47_40 = io_outValid_40 & _T_71659; // @[Switch.scala 41:38:@32819.4]
  assign _T_71662 = select_41 == 6'h2f; // @[Switch.scala 41:52:@32821.4]
  assign output_47_41 = io_outValid_41 & _T_71662; // @[Switch.scala 41:38:@32822.4]
  assign _T_71665 = select_42 == 6'h2f; // @[Switch.scala 41:52:@32824.4]
  assign output_47_42 = io_outValid_42 & _T_71665; // @[Switch.scala 41:38:@32825.4]
  assign _T_71668 = select_43 == 6'h2f; // @[Switch.scala 41:52:@32827.4]
  assign output_47_43 = io_outValid_43 & _T_71668; // @[Switch.scala 41:38:@32828.4]
  assign _T_71671 = select_44 == 6'h2f; // @[Switch.scala 41:52:@32830.4]
  assign output_47_44 = io_outValid_44 & _T_71671; // @[Switch.scala 41:38:@32831.4]
  assign _T_71674 = select_45 == 6'h2f; // @[Switch.scala 41:52:@32833.4]
  assign output_47_45 = io_outValid_45 & _T_71674; // @[Switch.scala 41:38:@32834.4]
  assign _T_71677 = select_46 == 6'h2f; // @[Switch.scala 41:52:@32836.4]
  assign output_47_46 = io_outValid_46 & _T_71677; // @[Switch.scala 41:38:@32837.4]
  assign _T_71680 = select_47 == 6'h2f; // @[Switch.scala 41:52:@32839.4]
  assign output_47_47 = io_outValid_47 & _T_71680; // @[Switch.scala 41:38:@32840.4]
  assign _T_71683 = select_48 == 6'h2f; // @[Switch.scala 41:52:@32842.4]
  assign output_47_48 = io_outValid_48 & _T_71683; // @[Switch.scala 41:38:@32843.4]
  assign _T_71686 = select_49 == 6'h2f; // @[Switch.scala 41:52:@32845.4]
  assign output_47_49 = io_outValid_49 & _T_71686; // @[Switch.scala 41:38:@32846.4]
  assign _T_71689 = select_50 == 6'h2f; // @[Switch.scala 41:52:@32848.4]
  assign output_47_50 = io_outValid_50 & _T_71689; // @[Switch.scala 41:38:@32849.4]
  assign _T_71692 = select_51 == 6'h2f; // @[Switch.scala 41:52:@32851.4]
  assign output_47_51 = io_outValid_51 & _T_71692; // @[Switch.scala 41:38:@32852.4]
  assign _T_71695 = select_52 == 6'h2f; // @[Switch.scala 41:52:@32854.4]
  assign output_47_52 = io_outValid_52 & _T_71695; // @[Switch.scala 41:38:@32855.4]
  assign _T_71698 = select_53 == 6'h2f; // @[Switch.scala 41:52:@32857.4]
  assign output_47_53 = io_outValid_53 & _T_71698; // @[Switch.scala 41:38:@32858.4]
  assign _T_71701 = select_54 == 6'h2f; // @[Switch.scala 41:52:@32860.4]
  assign output_47_54 = io_outValid_54 & _T_71701; // @[Switch.scala 41:38:@32861.4]
  assign _T_71704 = select_55 == 6'h2f; // @[Switch.scala 41:52:@32863.4]
  assign output_47_55 = io_outValid_55 & _T_71704; // @[Switch.scala 41:38:@32864.4]
  assign _T_71707 = select_56 == 6'h2f; // @[Switch.scala 41:52:@32866.4]
  assign output_47_56 = io_outValid_56 & _T_71707; // @[Switch.scala 41:38:@32867.4]
  assign _T_71710 = select_57 == 6'h2f; // @[Switch.scala 41:52:@32869.4]
  assign output_47_57 = io_outValid_57 & _T_71710; // @[Switch.scala 41:38:@32870.4]
  assign _T_71713 = select_58 == 6'h2f; // @[Switch.scala 41:52:@32872.4]
  assign output_47_58 = io_outValid_58 & _T_71713; // @[Switch.scala 41:38:@32873.4]
  assign _T_71716 = select_59 == 6'h2f; // @[Switch.scala 41:52:@32875.4]
  assign output_47_59 = io_outValid_59 & _T_71716; // @[Switch.scala 41:38:@32876.4]
  assign _T_71719 = select_60 == 6'h2f; // @[Switch.scala 41:52:@32878.4]
  assign output_47_60 = io_outValid_60 & _T_71719; // @[Switch.scala 41:38:@32879.4]
  assign _T_71722 = select_61 == 6'h2f; // @[Switch.scala 41:52:@32881.4]
  assign output_47_61 = io_outValid_61 & _T_71722; // @[Switch.scala 41:38:@32882.4]
  assign _T_71725 = select_62 == 6'h2f; // @[Switch.scala 41:52:@32884.4]
  assign output_47_62 = io_outValid_62 & _T_71725; // @[Switch.scala 41:38:@32885.4]
  assign _T_71728 = select_63 == 6'h2f; // @[Switch.scala 41:52:@32887.4]
  assign output_47_63 = io_outValid_63 & _T_71728; // @[Switch.scala 41:38:@32888.4]
  assign _T_71736 = {output_47_7,output_47_6,output_47_5,output_47_4,output_47_3,output_47_2,output_47_1,output_47_0}; // @[Switch.scala 43:31:@32896.4]
  assign _T_71744 = {output_47_15,output_47_14,output_47_13,output_47_12,output_47_11,output_47_10,output_47_9,output_47_8,_T_71736}; // @[Switch.scala 43:31:@32904.4]
  assign _T_71751 = {output_47_23,output_47_22,output_47_21,output_47_20,output_47_19,output_47_18,output_47_17,output_47_16}; // @[Switch.scala 43:31:@32911.4]
  assign _T_71760 = {output_47_31,output_47_30,output_47_29,output_47_28,output_47_27,output_47_26,output_47_25,output_47_24,_T_71751,_T_71744}; // @[Switch.scala 43:31:@32920.4]
  assign _T_71767 = {output_47_39,output_47_38,output_47_37,output_47_36,output_47_35,output_47_34,output_47_33,output_47_32}; // @[Switch.scala 43:31:@32927.4]
  assign _T_71775 = {output_47_47,output_47_46,output_47_45,output_47_44,output_47_43,output_47_42,output_47_41,output_47_40,_T_71767}; // @[Switch.scala 43:31:@32935.4]
  assign _T_71782 = {output_47_55,output_47_54,output_47_53,output_47_52,output_47_51,output_47_50,output_47_49,output_47_48}; // @[Switch.scala 43:31:@32942.4]
  assign _T_71791 = {output_47_63,output_47_62,output_47_61,output_47_60,output_47_59,output_47_58,output_47_57,output_47_56,_T_71782,_T_71775}; // @[Switch.scala 43:31:@32951.4]
  assign _T_71792 = {_T_71791,_T_71760}; // @[Switch.scala 43:31:@32952.4]
  assign _T_71796 = select_0 == 6'h30; // @[Switch.scala 41:52:@32955.4]
  assign output_48_0 = io_outValid_0 & _T_71796; // @[Switch.scala 41:38:@32956.4]
  assign _T_71799 = select_1 == 6'h30; // @[Switch.scala 41:52:@32958.4]
  assign output_48_1 = io_outValid_1 & _T_71799; // @[Switch.scala 41:38:@32959.4]
  assign _T_71802 = select_2 == 6'h30; // @[Switch.scala 41:52:@32961.4]
  assign output_48_2 = io_outValid_2 & _T_71802; // @[Switch.scala 41:38:@32962.4]
  assign _T_71805 = select_3 == 6'h30; // @[Switch.scala 41:52:@32964.4]
  assign output_48_3 = io_outValid_3 & _T_71805; // @[Switch.scala 41:38:@32965.4]
  assign _T_71808 = select_4 == 6'h30; // @[Switch.scala 41:52:@32967.4]
  assign output_48_4 = io_outValid_4 & _T_71808; // @[Switch.scala 41:38:@32968.4]
  assign _T_71811 = select_5 == 6'h30; // @[Switch.scala 41:52:@32970.4]
  assign output_48_5 = io_outValid_5 & _T_71811; // @[Switch.scala 41:38:@32971.4]
  assign _T_71814 = select_6 == 6'h30; // @[Switch.scala 41:52:@32973.4]
  assign output_48_6 = io_outValid_6 & _T_71814; // @[Switch.scala 41:38:@32974.4]
  assign _T_71817 = select_7 == 6'h30; // @[Switch.scala 41:52:@32976.4]
  assign output_48_7 = io_outValid_7 & _T_71817; // @[Switch.scala 41:38:@32977.4]
  assign _T_71820 = select_8 == 6'h30; // @[Switch.scala 41:52:@32979.4]
  assign output_48_8 = io_outValid_8 & _T_71820; // @[Switch.scala 41:38:@32980.4]
  assign _T_71823 = select_9 == 6'h30; // @[Switch.scala 41:52:@32982.4]
  assign output_48_9 = io_outValid_9 & _T_71823; // @[Switch.scala 41:38:@32983.4]
  assign _T_71826 = select_10 == 6'h30; // @[Switch.scala 41:52:@32985.4]
  assign output_48_10 = io_outValid_10 & _T_71826; // @[Switch.scala 41:38:@32986.4]
  assign _T_71829 = select_11 == 6'h30; // @[Switch.scala 41:52:@32988.4]
  assign output_48_11 = io_outValid_11 & _T_71829; // @[Switch.scala 41:38:@32989.4]
  assign _T_71832 = select_12 == 6'h30; // @[Switch.scala 41:52:@32991.4]
  assign output_48_12 = io_outValid_12 & _T_71832; // @[Switch.scala 41:38:@32992.4]
  assign _T_71835 = select_13 == 6'h30; // @[Switch.scala 41:52:@32994.4]
  assign output_48_13 = io_outValid_13 & _T_71835; // @[Switch.scala 41:38:@32995.4]
  assign _T_71838 = select_14 == 6'h30; // @[Switch.scala 41:52:@32997.4]
  assign output_48_14 = io_outValid_14 & _T_71838; // @[Switch.scala 41:38:@32998.4]
  assign _T_71841 = select_15 == 6'h30; // @[Switch.scala 41:52:@33000.4]
  assign output_48_15 = io_outValid_15 & _T_71841; // @[Switch.scala 41:38:@33001.4]
  assign _T_71844 = select_16 == 6'h30; // @[Switch.scala 41:52:@33003.4]
  assign output_48_16 = io_outValid_16 & _T_71844; // @[Switch.scala 41:38:@33004.4]
  assign _T_71847 = select_17 == 6'h30; // @[Switch.scala 41:52:@33006.4]
  assign output_48_17 = io_outValid_17 & _T_71847; // @[Switch.scala 41:38:@33007.4]
  assign _T_71850 = select_18 == 6'h30; // @[Switch.scala 41:52:@33009.4]
  assign output_48_18 = io_outValid_18 & _T_71850; // @[Switch.scala 41:38:@33010.4]
  assign _T_71853 = select_19 == 6'h30; // @[Switch.scala 41:52:@33012.4]
  assign output_48_19 = io_outValid_19 & _T_71853; // @[Switch.scala 41:38:@33013.4]
  assign _T_71856 = select_20 == 6'h30; // @[Switch.scala 41:52:@33015.4]
  assign output_48_20 = io_outValid_20 & _T_71856; // @[Switch.scala 41:38:@33016.4]
  assign _T_71859 = select_21 == 6'h30; // @[Switch.scala 41:52:@33018.4]
  assign output_48_21 = io_outValid_21 & _T_71859; // @[Switch.scala 41:38:@33019.4]
  assign _T_71862 = select_22 == 6'h30; // @[Switch.scala 41:52:@33021.4]
  assign output_48_22 = io_outValid_22 & _T_71862; // @[Switch.scala 41:38:@33022.4]
  assign _T_71865 = select_23 == 6'h30; // @[Switch.scala 41:52:@33024.4]
  assign output_48_23 = io_outValid_23 & _T_71865; // @[Switch.scala 41:38:@33025.4]
  assign _T_71868 = select_24 == 6'h30; // @[Switch.scala 41:52:@33027.4]
  assign output_48_24 = io_outValid_24 & _T_71868; // @[Switch.scala 41:38:@33028.4]
  assign _T_71871 = select_25 == 6'h30; // @[Switch.scala 41:52:@33030.4]
  assign output_48_25 = io_outValid_25 & _T_71871; // @[Switch.scala 41:38:@33031.4]
  assign _T_71874 = select_26 == 6'h30; // @[Switch.scala 41:52:@33033.4]
  assign output_48_26 = io_outValid_26 & _T_71874; // @[Switch.scala 41:38:@33034.4]
  assign _T_71877 = select_27 == 6'h30; // @[Switch.scala 41:52:@33036.4]
  assign output_48_27 = io_outValid_27 & _T_71877; // @[Switch.scala 41:38:@33037.4]
  assign _T_71880 = select_28 == 6'h30; // @[Switch.scala 41:52:@33039.4]
  assign output_48_28 = io_outValid_28 & _T_71880; // @[Switch.scala 41:38:@33040.4]
  assign _T_71883 = select_29 == 6'h30; // @[Switch.scala 41:52:@33042.4]
  assign output_48_29 = io_outValid_29 & _T_71883; // @[Switch.scala 41:38:@33043.4]
  assign _T_71886 = select_30 == 6'h30; // @[Switch.scala 41:52:@33045.4]
  assign output_48_30 = io_outValid_30 & _T_71886; // @[Switch.scala 41:38:@33046.4]
  assign _T_71889 = select_31 == 6'h30; // @[Switch.scala 41:52:@33048.4]
  assign output_48_31 = io_outValid_31 & _T_71889; // @[Switch.scala 41:38:@33049.4]
  assign _T_71892 = select_32 == 6'h30; // @[Switch.scala 41:52:@33051.4]
  assign output_48_32 = io_outValid_32 & _T_71892; // @[Switch.scala 41:38:@33052.4]
  assign _T_71895 = select_33 == 6'h30; // @[Switch.scala 41:52:@33054.4]
  assign output_48_33 = io_outValid_33 & _T_71895; // @[Switch.scala 41:38:@33055.4]
  assign _T_71898 = select_34 == 6'h30; // @[Switch.scala 41:52:@33057.4]
  assign output_48_34 = io_outValid_34 & _T_71898; // @[Switch.scala 41:38:@33058.4]
  assign _T_71901 = select_35 == 6'h30; // @[Switch.scala 41:52:@33060.4]
  assign output_48_35 = io_outValid_35 & _T_71901; // @[Switch.scala 41:38:@33061.4]
  assign _T_71904 = select_36 == 6'h30; // @[Switch.scala 41:52:@33063.4]
  assign output_48_36 = io_outValid_36 & _T_71904; // @[Switch.scala 41:38:@33064.4]
  assign _T_71907 = select_37 == 6'h30; // @[Switch.scala 41:52:@33066.4]
  assign output_48_37 = io_outValid_37 & _T_71907; // @[Switch.scala 41:38:@33067.4]
  assign _T_71910 = select_38 == 6'h30; // @[Switch.scala 41:52:@33069.4]
  assign output_48_38 = io_outValid_38 & _T_71910; // @[Switch.scala 41:38:@33070.4]
  assign _T_71913 = select_39 == 6'h30; // @[Switch.scala 41:52:@33072.4]
  assign output_48_39 = io_outValid_39 & _T_71913; // @[Switch.scala 41:38:@33073.4]
  assign _T_71916 = select_40 == 6'h30; // @[Switch.scala 41:52:@33075.4]
  assign output_48_40 = io_outValid_40 & _T_71916; // @[Switch.scala 41:38:@33076.4]
  assign _T_71919 = select_41 == 6'h30; // @[Switch.scala 41:52:@33078.4]
  assign output_48_41 = io_outValid_41 & _T_71919; // @[Switch.scala 41:38:@33079.4]
  assign _T_71922 = select_42 == 6'h30; // @[Switch.scala 41:52:@33081.4]
  assign output_48_42 = io_outValid_42 & _T_71922; // @[Switch.scala 41:38:@33082.4]
  assign _T_71925 = select_43 == 6'h30; // @[Switch.scala 41:52:@33084.4]
  assign output_48_43 = io_outValid_43 & _T_71925; // @[Switch.scala 41:38:@33085.4]
  assign _T_71928 = select_44 == 6'h30; // @[Switch.scala 41:52:@33087.4]
  assign output_48_44 = io_outValid_44 & _T_71928; // @[Switch.scala 41:38:@33088.4]
  assign _T_71931 = select_45 == 6'h30; // @[Switch.scala 41:52:@33090.4]
  assign output_48_45 = io_outValid_45 & _T_71931; // @[Switch.scala 41:38:@33091.4]
  assign _T_71934 = select_46 == 6'h30; // @[Switch.scala 41:52:@33093.4]
  assign output_48_46 = io_outValid_46 & _T_71934; // @[Switch.scala 41:38:@33094.4]
  assign _T_71937 = select_47 == 6'h30; // @[Switch.scala 41:52:@33096.4]
  assign output_48_47 = io_outValid_47 & _T_71937; // @[Switch.scala 41:38:@33097.4]
  assign _T_71940 = select_48 == 6'h30; // @[Switch.scala 41:52:@33099.4]
  assign output_48_48 = io_outValid_48 & _T_71940; // @[Switch.scala 41:38:@33100.4]
  assign _T_71943 = select_49 == 6'h30; // @[Switch.scala 41:52:@33102.4]
  assign output_48_49 = io_outValid_49 & _T_71943; // @[Switch.scala 41:38:@33103.4]
  assign _T_71946 = select_50 == 6'h30; // @[Switch.scala 41:52:@33105.4]
  assign output_48_50 = io_outValid_50 & _T_71946; // @[Switch.scala 41:38:@33106.4]
  assign _T_71949 = select_51 == 6'h30; // @[Switch.scala 41:52:@33108.4]
  assign output_48_51 = io_outValid_51 & _T_71949; // @[Switch.scala 41:38:@33109.4]
  assign _T_71952 = select_52 == 6'h30; // @[Switch.scala 41:52:@33111.4]
  assign output_48_52 = io_outValid_52 & _T_71952; // @[Switch.scala 41:38:@33112.4]
  assign _T_71955 = select_53 == 6'h30; // @[Switch.scala 41:52:@33114.4]
  assign output_48_53 = io_outValid_53 & _T_71955; // @[Switch.scala 41:38:@33115.4]
  assign _T_71958 = select_54 == 6'h30; // @[Switch.scala 41:52:@33117.4]
  assign output_48_54 = io_outValid_54 & _T_71958; // @[Switch.scala 41:38:@33118.4]
  assign _T_71961 = select_55 == 6'h30; // @[Switch.scala 41:52:@33120.4]
  assign output_48_55 = io_outValid_55 & _T_71961; // @[Switch.scala 41:38:@33121.4]
  assign _T_71964 = select_56 == 6'h30; // @[Switch.scala 41:52:@33123.4]
  assign output_48_56 = io_outValid_56 & _T_71964; // @[Switch.scala 41:38:@33124.4]
  assign _T_71967 = select_57 == 6'h30; // @[Switch.scala 41:52:@33126.4]
  assign output_48_57 = io_outValid_57 & _T_71967; // @[Switch.scala 41:38:@33127.4]
  assign _T_71970 = select_58 == 6'h30; // @[Switch.scala 41:52:@33129.4]
  assign output_48_58 = io_outValid_58 & _T_71970; // @[Switch.scala 41:38:@33130.4]
  assign _T_71973 = select_59 == 6'h30; // @[Switch.scala 41:52:@33132.4]
  assign output_48_59 = io_outValid_59 & _T_71973; // @[Switch.scala 41:38:@33133.4]
  assign _T_71976 = select_60 == 6'h30; // @[Switch.scala 41:52:@33135.4]
  assign output_48_60 = io_outValid_60 & _T_71976; // @[Switch.scala 41:38:@33136.4]
  assign _T_71979 = select_61 == 6'h30; // @[Switch.scala 41:52:@33138.4]
  assign output_48_61 = io_outValid_61 & _T_71979; // @[Switch.scala 41:38:@33139.4]
  assign _T_71982 = select_62 == 6'h30; // @[Switch.scala 41:52:@33141.4]
  assign output_48_62 = io_outValid_62 & _T_71982; // @[Switch.scala 41:38:@33142.4]
  assign _T_71985 = select_63 == 6'h30; // @[Switch.scala 41:52:@33144.4]
  assign output_48_63 = io_outValid_63 & _T_71985; // @[Switch.scala 41:38:@33145.4]
  assign _T_71993 = {output_48_7,output_48_6,output_48_5,output_48_4,output_48_3,output_48_2,output_48_1,output_48_0}; // @[Switch.scala 43:31:@33153.4]
  assign _T_72001 = {output_48_15,output_48_14,output_48_13,output_48_12,output_48_11,output_48_10,output_48_9,output_48_8,_T_71993}; // @[Switch.scala 43:31:@33161.4]
  assign _T_72008 = {output_48_23,output_48_22,output_48_21,output_48_20,output_48_19,output_48_18,output_48_17,output_48_16}; // @[Switch.scala 43:31:@33168.4]
  assign _T_72017 = {output_48_31,output_48_30,output_48_29,output_48_28,output_48_27,output_48_26,output_48_25,output_48_24,_T_72008,_T_72001}; // @[Switch.scala 43:31:@33177.4]
  assign _T_72024 = {output_48_39,output_48_38,output_48_37,output_48_36,output_48_35,output_48_34,output_48_33,output_48_32}; // @[Switch.scala 43:31:@33184.4]
  assign _T_72032 = {output_48_47,output_48_46,output_48_45,output_48_44,output_48_43,output_48_42,output_48_41,output_48_40,_T_72024}; // @[Switch.scala 43:31:@33192.4]
  assign _T_72039 = {output_48_55,output_48_54,output_48_53,output_48_52,output_48_51,output_48_50,output_48_49,output_48_48}; // @[Switch.scala 43:31:@33199.4]
  assign _T_72048 = {output_48_63,output_48_62,output_48_61,output_48_60,output_48_59,output_48_58,output_48_57,output_48_56,_T_72039,_T_72032}; // @[Switch.scala 43:31:@33208.4]
  assign _T_72049 = {_T_72048,_T_72017}; // @[Switch.scala 43:31:@33209.4]
  assign _T_72053 = select_0 == 6'h31; // @[Switch.scala 41:52:@33212.4]
  assign output_49_0 = io_outValid_0 & _T_72053; // @[Switch.scala 41:38:@33213.4]
  assign _T_72056 = select_1 == 6'h31; // @[Switch.scala 41:52:@33215.4]
  assign output_49_1 = io_outValid_1 & _T_72056; // @[Switch.scala 41:38:@33216.4]
  assign _T_72059 = select_2 == 6'h31; // @[Switch.scala 41:52:@33218.4]
  assign output_49_2 = io_outValid_2 & _T_72059; // @[Switch.scala 41:38:@33219.4]
  assign _T_72062 = select_3 == 6'h31; // @[Switch.scala 41:52:@33221.4]
  assign output_49_3 = io_outValid_3 & _T_72062; // @[Switch.scala 41:38:@33222.4]
  assign _T_72065 = select_4 == 6'h31; // @[Switch.scala 41:52:@33224.4]
  assign output_49_4 = io_outValid_4 & _T_72065; // @[Switch.scala 41:38:@33225.4]
  assign _T_72068 = select_5 == 6'h31; // @[Switch.scala 41:52:@33227.4]
  assign output_49_5 = io_outValid_5 & _T_72068; // @[Switch.scala 41:38:@33228.4]
  assign _T_72071 = select_6 == 6'h31; // @[Switch.scala 41:52:@33230.4]
  assign output_49_6 = io_outValid_6 & _T_72071; // @[Switch.scala 41:38:@33231.4]
  assign _T_72074 = select_7 == 6'h31; // @[Switch.scala 41:52:@33233.4]
  assign output_49_7 = io_outValid_7 & _T_72074; // @[Switch.scala 41:38:@33234.4]
  assign _T_72077 = select_8 == 6'h31; // @[Switch.scala 41:52:@33236.4]
  assign output_49_8 = io_outValid_8 & _T_72077; // @[Switch.scala 41:38:@33237.4]
  assign _T_72080 = select_9 == 6'h31; // @[Switch.scala 41:52:@33239.4]
  assign output_49_9 = io_outValid_9 & _T_72080; // @[Switch.scala 41:38:@33240.4]
  assign _T_72083 = select_10 == 6'h31; // @[Switch.scala 41:52:@33242.4]
  assign output_49_10 = io_outValid_10 & _T_72083; // @[Switch.scala 41:38:@33243.4]
  assign _T_72086 = select_11 == 6'h31; // @[Switch.scala 41:52:@33245.4]
  assign output_49_11 = io_outValid_11 & _T_72086; // @[Switch.scala 41:38:@33246.4]
  assign _T_72089 = select_12 == 6'h31; // @[Switch.scala 41:52:@33248.4]
  assign output_49_12 = io_outValid_12 & _T_72089; // @[Switch.scala 41:38:@33249.4]
  assign _T_72092 = select_13 == 6'h31; // @[Switch.scala 41:52:@33251.4]
  assign output_49_13 = io_outValid_13 & _T_72092; // @[Switch.scala 41:38:@33252.4]
  assign _T_72095 = select_14 == 6'h31; // @[Switch.scala 41:52:@33254.4]
  assign output_49_14 = io_outValid_14 & _T_72095; // @[Switch.scala 41:38:@33255.4]
  assign _T_72098 = select_15 == 6'h31; // @[Switch.scala 41:52:@33257.4]
  assign output_49_15 = io_outValid_15 & _T_72098; // @[Switch.scala 41:38:@33258.4]
  assign _T_72101 = select_16 == 6'h31; // @[Switch.scala 41:52:@33260.4]
  assign output_49_16 = io_outValid_16 & _T_72101; // @[Switch.scala 41:38:@33261.4]
  assign _T_72104 = select_17 == 6'h31; // @[Switch.scala 41:52:@33263.4]
  assign output_49_17 = io_outValid_17 & _T_72104; // @[Switch.scala 41:38:@33264.4]
  assign _T_72107 = select_18 == 6'h31; // @[Switch.scala 41:52:@33266.4]
  assign output_49_18 = io_outValid_18 & _T_72107; // @[Switch.scala 41:38:@33267.4]
  assign _T_72110 = select_19 == 6'h31; // @[Switch.scala 41:52:@33269.4]
  assign output_49_19 = io_outValid_19 & _T_72110; // @[Switch.scala 41:38:@33270.4]
  assign _T_72113 = select_20 == 6'h31; // @[Switch.scala 41:52:@33272.4]
  assign output_49_20 = io_outValid_20 & _T_72113; // @[Switch.scala 41:38:@33273.4]
  assign _T_72116 = select_21 == 6'h31; // @[Switch.scala 41:52:@33275.4]
  assign output_49_21 = io_outValid_21 & _T_72116; // @[Switch.scala 41:38:@33276.4]
  assign _T_72119 = select_22 == 6'h31; // @[Switch.scala 41:52:@33278.4]
  assign output_49_22 = io_outValid_22 & _T_72119; // @[Switch.scala 41:38:@33279.4]
  assign _T_72122 = select_23 == 6'h31; // @[Switch.scala 41:52:@33281.4]
  assign output_49_23 = io_outValid_23 & _T_72122; // @[Switch.scala 41:38:@33282.4]
  assign _T_72125 = select_24 == 6'h31; // @[Switch.scala 41:52:@33284.4]
  assign output_49_24 = io_outValid_24 & _T_72125; // @[Switch.scala 41:38:@33285.4]
  assign _T_72128 = select_25 == 6'h31; // @[Switch.scala 41:52:@33287.4]
  assign output_49_25 = io_outValid_25 & _T_72128; // @[Switch.scala 41:38:@33288.4]
  assign _T_72131 = select_26 == 6'h31; // @[Switch.scala 41:52:@33290.4]
  assign output_49_26 = io_outValid_26 & _T_72131; // @[Switch.scala 41:38:@33291.4]
  assign _T_72134 = select_27 == 6'h31; // @[Switch.scala 41:52:@33293.4]
  assign output_49_27 = io_outValid_27 & _T_72134; // @[Switch.scala 41:38:@33294.4]
  assign _T_72137 = select_28 == 6'h31; // @[Switch.scala 41:52:@33296.4]
  assign output_49_28 = io_outValid_28 & _T_72137; // @[Switch.scala 41:38:@33297.4]
  assign _T_72140 = select_29 == 6'h31; // @[Switch.scala 41:52:@33299.4]
  assign output_49_29 = io_outValid_29 & _T_72140; // @[Switch.scala 41:38:@33300.4]
  assign _T_72143 = select_30 == 6'h31; // @[Switch.scala 41:52:@33302.4]
  assign output_49_30 = io_outValid_30 & _T_72143; // @[Switch.scala 41:38:@33303.4]
  assign _T_72146 = select_31 == 6'h31; // @[Switch.scala 41:52:@33305.4]
  assign output_49_31 = io_outValid_31 & _T_72146; // @[Switch.scala 41:38:@33306.4]
  assign _T_72149 = select_32 == 6'h31; // @[Switch.scala 41:52:@33308.4]
  assign output_49_32 = io_outValid_32 & _T_72149; // @[Switch.scala 41:38:@33309.4]
  assign _T_72152 = select_33 == 6'h31; // @[Switch.scala 41:52:@33311.4]
  assign output_49_33 = io_outValid_33 & _T_72152; // @[Switch.scala 41:38:@33312.4]
  assign _T_72155 = select_34 == 6'h31; // @[Switch.scala 41:52:@33314.4]
  assign output_49_34 = io_outValid_34 & _T_72155; // @[Switch.scala 41:38:@33315.4]
  assign _T_72158 = select_35 == 6'h31; // @[Switch.scala 41:52:@33317.4]
  assign output_49_35 = io_outValid_35 & _T_72158; // @[Switch.scala 41:38:@33318.4]
  assign _T_72161 = select_36 == 6'h31; // @[Switch.scala 41:52:@33320.4]
  assign output_49_36 = io_outValid_36 & _T_72161; // @[Switch.scala 41:38:@33321.4]
  assign _T_72164 = select_37 == 6'h31; // @[Switch.scala 41:52:@33323.4]
  assign output_49_37 = io_outValid_37 & _T_72164; // @[Switch.scala 41:38:@33324.4]
  assign _T_72167 = select_38 == 6'h31; // @[Switch.scala 41:52:@33326.4]
  assign output_49_38 = io_outValid_38 & _T_72167; // @[Switch.scala 41:38:@33327.4]
  assign _T_72170 = select_39 == 6'h31; // @[Switch.scala 41:52:@33329.4]
  assign output_49_39 = io_outValid_39 & _T_72170; // @[Switch.scala 41:38:@33330.4]
  assign _T_72173 = select_40 == 6'h31; // @[Switch.scala 41:52:@33332.4]
  assign output_49_40 = io_outValid_40 & _T_72173; // @[Switch.scala 41:38:@33333.4]
  assign _T_72176 = select_41 == 6'h31; // @[Switch.scala 41:52:@33335.4]
  assign output_49_41 = io_outValid_41 & _T_72176; // @[Switch.scala 41:38:@33336.4]
  assign _T_72179 = select_42 == 6'h31; // @[Switch.scala 41:52:@33338.4]
  assign output_49_42 = io_outValid_42 & _T_72179; // @[Switch.scala 41:38:@33339.4]
  assign _T_72182 = select_43 == 6'h31; // @[Switch.scala 41:52:@33341.4]
  assign output_49_43 = io_outValid_43 & _T_72182; // @[Switch.scala 41:38:@33342.4]
  assign _T_72185 = select_44 == 6'h31; // @[Switch.scala 41:52:@33344.4]
  assign output_49_44 = io_outValid_44 & _T_72185; // @[Switch.scala 41:38:@33345.4]
  assign _T_72188 = select_45 == 6'h31; // @[Switch.scala 41:52:@33347.4]
  assign output_49_45 = io_outValid_45 & _T_72188; // @[Switch.scala 41:38:@33348.4]
  assign _T_72191 = select_46 == 6'h31; // @[Switch.scala 41:52:@33350.4]
  assign output_49_46 = io_outValid_46 & _T_72191; // @[Switch.scala 41:38:@33351.4]
  assign _T_72194 = select_47 == 6'h31; // @[Switch.scala 41:52:@33353.4]
  assign output_49_47 = io_outValid_47 & _T_72194; // @[Switch.scala 41:38:@33354.4]
  assign _T_72197 = select_48 == 6'h31; // @[Switch.scala 41:52:@33356.4]
  assign output_49_48 = io_outValid_48 & _T_72197; // @[Switch.scala 41:38:@33357.4]
  assign _T_72200 = select_49 == 6'h31; // @[Switch.scala 41:52:@33359.4]
  assign output_49_49 = io_outValid_49 & _T_72200; // @[Switch.scala 41:38:@33360.4]
  assign _T_72203 = select_50 == 6'h31; // @[Switch.scala 41:52:@33362.4]
  assign output_49_50 = io_outValid_50 & _T_72203; // @[Switch.scala 41:38:@33363.4]
  assign _T_72206 = select_51 == 6'h31; // @[Switch.scala 41:52:@33365.4]
  assign output_49_51 = io_outValid_51 & _T_72206; // @[Switch.scala 41:38:@33366.4]
  assign _T_72209 = select_52 == 6'h31; // @[Switch.scala 41:52:@33368.4]
  assign output_49_52 = io_outValid_52 & _T_72209; // @[Switch.scala 41:38:@33369.4]
  assign _T_72212 = select_53 == 6'h31; // @[Switch.scala 41:52:@33371.4]
  assign output_49_53 = io_outValid_53 & _T_72212; // @[Switch.scala 41:38:@33372.4]
  assign _T_72215 = select_54 == 6'h31; // @[Switch.scala 41:52:@33374.4]
  assign output_49_54 = io_outValid_54 & _T_72215; // @[Switch.scala 41:38:@33375.4]
  assign _T_72218 = select_55 == 6'h31; // @[Switch.scala 41:52:@33377.4]
  assign output_49_55 = io_outValid_55 & _T_72218; // @[Switch.scala 41:38:@33378.4]
  assign _T_72221 = select_56 == 6'h31; // @[Switch.scala 41:52:@33380.4]
  assign output_49_56 = io_outValid_56 & _T_72221; // @[Switch.scala 41:38:@33381.4]
  assign _T_72224 = select_57 == 6'h31; // @[Switch.scala 41:52:@33383.4]
  assign output_49_57 = io_outValid_57 & _T_72224; // @[Switch.scala 41:38:@33384.4]
  assign _T_72227 = select_58 == 6'h31; // @[Switch.scala 41:52:@33386.4]
  assign output_49_58 = io_outValid_58 & _T_72227; // @[Switch.scala 41:38:@33387.4]
  assign _T_72230 = select_59 == 6'h31; // @[Switch.scala 41:52:@33389.4]
  assign output_49_59 = io_outValid_59 & _T_72230; // @[Switch.scala 41:38:@33390.4]
  assign _T_72233 = select_60 == 6'h31; // @[Switch.scala 41:52:@33392.4]
  assign output_49_60 = io_outValid_60 & _T_72233; // @[Switch.scala 41:38:@33393.4]
  assign _T_72236 = select_61 == 6'h31; // @[Switch.scala 41:52:@33395.4]
  assign output_49_61 = io_outValid_61 & _T_72236; // @[Switch.scala 41:38:@33396.4]
  assign _T_72239 = select_62 == 6'h31; // @[Switch.scala 41:52:@33398.4]
  assign output_49_62 = io_outValid_62 & _T_72239; // @[Switch.scala 41:38:@33399.4]
  assign _T_72242 = select_63 == 6'h31; // @[Switch.scala 41:52:@33401.4]
  assign output_49_63 = io_outValid_63 & _T_72242; // @[Switch.scala 41:38:@33402.4]
  assign _T_72250 = {output_49_7,output_49_6,output_49_5,output_49_4,output_49_3,output_49_2,output_49_1,output_49_0}; // @[Switch.scala 43:31:@33410.4]
  assign _T_72258 = {output_49_15,output_49_14,output_49_13,output_49_12,output_49_11,output_49_10,output_49_9,output_49_8,_T_72250}; // @[Switch.scala 43:31:@33418.4]
  assign _T_72265 = {output_49_23,output_49_22,output_49_21,output_49_20,output_49_19,output_49_18,output_49_17,output_49_16}; // @[Switch.scala 43:31:@33425.4]
  assign _T_72274 = {output_49_31,output_49_30,output_49_29,output_49_28,output_49_27,output_49_26,output_49_25,output_49_24,_T_72265,_T_72258}; // @[Switch.scala 43:31:@33434.4]
  assign _T_72281 = {output_49_39,output_49_38,output_49_37,output_49_36,output_49_35,output_49_34,output_49_33,output_49_32}; // @[Switch.scala 43:31:@33441.4]
  assign _T_72289 = {output_49_47,output_49_46,output_49_45,output_49_44,output_49_43,output_49_42,output_49_41,output_49_40,_T_72281}; // @[Switch.scala 43:31:@33449.4]
  assign _T_72296 = {output_49_55,output_49_54,output_49_53,output_49_52,output_49_51,output_49_50,output_49_49,output_49_48}; // @[Switch.scala 43:31:@33456.4]
  assign _T_72305 = {output_49_63,output_49_62,output_49_61,output_49_60,output_49_59,output_49_58,output_49_57,output_49_56,_T_72296,_T_72289}; // @[Switch.scala 43:31:@33465.4]
  assign _T_72306 = {_T_72305,_T_72274}; // @[Switch.scala 43:31:@33466.4]
  assign _T_72310 = select_0 == 6'h32; // @[Switch.scala 41:52:@33469.4]
  assign output_50_0 = io_outValid_0 & _T_72310; // @[Switch.scala 41:38:@33470.4]
  assign _T_72313 = select_1 == 6'h32; // @[Switch.scala 41:52:@33472.4]
  assign output_50_1 = io_outValid_1 & _T_72313; // @[Switch.scala 41:38:@33473.4]
  assign _T_72316 = select_2 == 6'h32; // @[Switch.scala 41:52:@33475.4]
  assign output_50_2 = io_outValid_2 & _T_72316; // @[Switch.scala 41:38:@33476.4]
  assign _T_72319 = select_3 == 6'h32; // @[Switch.scala 41:52:@33478.4]
  assign output_50_3 = io_outValid_3 & _T_72319; // @[Switch.scala 41:38:@33479.4]
  assign _T_72322 = select_4 == 6'h32; // @[Switch.scala 41:52:@33481.4]
  assign output_50_4 = io_outValid_4 & _T_72322; // @[Switch.scala 41:38:@33482.4]
  assign _T_72325 = select_5 == 6'h32; // @[Switch.scala 41:52:@33484.4]
  assign output_50_5 = io_outValid_5 & _T_72325; // @[Switch.scala 41:38:@33485.4]
  assign _T_72328 = select_6 == 6'h32; // @[Switch.scala 41:52:@33487.4]
  assign output_50_6 = io_outValid_6 & _T_72328; // @[Switch.scala 41:38:@33488.4]
  assign _T_72331 = select_7 == 6'h32; // @[Switch.scala 41:52:@33490.4]
  assign output_50_7 = io_outValid_7 & _T_72331; // @[Switch.scala 41:38:@33491.4]
  assign _T_72334 = select_8 == 6'h32; // @[Switch.scala 41:52:@33493.4]
  assign output_50_8 = io_outValid_8 & _T_72334; // @[Switch.scala 41:38:@33494.4]
  assign _T_72337 = select_9 == 6'h32; // @[Switch.scala 41:52:@33496.4]
  assign output_50_9 = io_outValid_9 & _T_72337; // @[Switch.scala 41:38:@33497.4]
  assign _T_72340 = select_10 == 6'h32; // @[Switch.scala 41:52:@33499.4]
  assign output_50_10 = io_outValid_10 & _T_72340; // @[Switch.scala 41:38:@33500.4]
  assign _T_72343 = select_11 == 6'h32; // @[Switch.scala 41:52:@33502.4]
  assign output_50_11 = io_outValid_11 & _T_72343; // @[Switch.scala 41:38:@33503.4]
  assign _T_72346 = select_12 == 6'h32; // @[Switch.scala 41:52:@33505.4]
  assign output_50_12 = io_outValid_12 & _T_72346; // @[Switch.scala 41:38:@33506.4]
  assign _T_72349 = select_13 == 6'h32; // @[Switch.scala 41:52:@33508.4]
  assign output_50_13 = io_outValid_13 & _T_72349; // @[Switch.scala 41:38:@33509.4]
  assign _T_72352 = select_14 == 6'h32; // @[Switch.scala 41:52:@33511.4]
  assign output_50_14 = io_outValid_14 & _T_72352; // @[Switch.scala 41:38:@33512.4]
  assign _T_72355 = select_15 == 6'h32; // @[Switch.scala 41:52:@33514.4]
  assign output_50_15 = io_outValid_15 & _T_72355; // @[Switch.scala 41:38:@33515.4]
  assign _T_72358 = select_16 == 6'h32; // @[Switch.scala 41:52:@33517.4]
  assign output_50_16 = io_outValid_16 & _T_72358; // @[Switch.scala 41:38:@33518.4]
  assign _T_72361 = select_17 == 6'h32; // @[Switch.scala 41:52:@33520.4]
  assign output_50_17 = io_outValid_17 & _T_72361; // @[Switch.scala 41:38:@33521.4]
  assign _T_72364 = select_18 == 6'h32; // @[Switch.scala 41:52:@33523.4]
  assign output_50_18 = io_outValid_18 & _T_72364; // @[Switch.scala 41:38:@33524.4]
  assign _T_72367 = select_19 == 6'h32; // @[Switch.scala 41:52:@33526.4]
  assign output_50_19 = io_outValid_19 & _T_72367; // @[Switch.scala 41:38:@33527.4]
  assign _T_72370 = select_20 == 6'h32; // @[Switch.scala 41:52:@33529.4]
  assign output_50_20 = io_outValid_20 & _T_72370; // @[Switch.scala 41:38:@33530.4]
  assign _T_72373 = select_21 == 6'h32; // @[Switch.scala 41:52:@33532.4]
  assign output_50_21 = io_outValid_21 & _T_72373; // @[Switch.scala 41:38:@33533.4]
  assign _T_72376 = select_22 == 6'h32; // @[Switch.scala 41:52:@33535.4]
  assign output_50_22 = io_outValid_22 & _T_72376; // @[Switch.scala 41:38:@33536.4]
  assign _T_72379 = select_23 == 6'h32; // @[Switch.scala 41:52:@33538.4]
  assign output_50_23 = io_outValid_23 & _T_72379; // @[Switch.scala 41:38:@33539.4]
  assign _T_72382 = select_24 == 6'h32; // @[Switch.scala 41:52:@33541.4]
  assign output_50_24 = io_outValid_24 & _T_72382; // @[Switch.scala 41:38:@33542.4]
  assign _T_72385 = select_25 == 6'h32; // @[Switch.scala 41:52:@33544.4]
  assign output_50_25 = io_outValid_25 & _T_72385; // @[Switch.scala 41:38:@33545.4]
  assign _T_72388 = select_26 == 6'h32; // @[Switch.scala 41:52:@33547.4]
  assign output_50_26 = io_outValid_26 & _T_72388; // @[Switch.scala 41:38:@33548.4]
  assign _T_72391 = select_27 == 6'h32; // @[Switch.scala 41:52:@33550.4]
  assign output_50_27 = io_outValid_27 & _T_72391; // @[Switch.scala 41:38:@33551.4]
  assign _T_72394 = select_28 == 6'h32; // @[Switch.scala 41:52:@33553.4]
  assign output_50_28 = io_outValid_28 & _T_72394; // @[Switch.scala 41:38:@33554.4]
  assign _T_72397 = select_29 == 6'h32; // @[Switch.scala 41:52:@33556.4]
  assign output_50_29 = io_outValid_29 & _T_72397; // @[Switch.scala 41:38:@33557.4]
  assign _T_72400 = select_30 == 6'h32; // @[Switch.scala 41:52:@33559.4]
  assign output_50_30 = io_outValid_30 & _T_72400; // @[Switch.scala 41:38:@33560.4]
  assign _T_72403 = select_31 == 6'h32; // @[Switch.scala 41:52:@33562.4]
  assign output_50_31 = io_outValid_31 & _T_72403; // @[Switch.scala 41:38:@33563.4]
  assign _T_72406 = select_32 == 6'h32; // @[Switch.scala 41:52:@33565.4]
  assign output_50_32 = io_outValid_32 & _T_72406; // @[Switch.scala 41:38:@33566.4]
  assign _T_72409 = select_33 == 6'h32; // @[Switch.scala 41:52:@33568.4]
  assign output_50_33 = io_outValid_33 & _T_72409; // @[Switch.scala 41:38:@33569.4]
  assign _T_72412 = select_34 == 6'h32; // @[Switch.scala 41:52:@33571.4]
  assign output_50_34 = io_outValid_34 & _T_72412; // @[Switch.scala 41:38:@33572.4]
  assign _T_72415 = select_35 == 6'h32; // @[Switch.scala 41:52:@33574.4]
  assign output_50_35 = io_outValid_35 & _T_72415; // @[Switch.scala 41:38:@33575.4]
  assign _T_72418 = select_36 == 6'h32; // @[Switch.scala 41:52:@33577.4]
  assign output_50_36 = io_outValid_36 & _T_72418; // @[Switch.scala 41:38:@33578.4]
  assign _T_72421 = select_37 == 6'h32; // @[Switch.scala 41:52:@33580.4]
  assign output_50_37 = io_outValid_37 & _T_72421; // @[Switch.scala 41:38:@33581.4]
  assign _T_72424 = select_38 == 6'h32; // @[Switch.scala 41:52:@33583.4]
  assign output_50_38 = io_outValid_38 & _T_72424; // @[Switch.scala 41:38:@33584.4]
  assign _T_72427 = select_39 == 6'h32; // @[Switch.scala 41:52:@33586.4]
  assign output_50_39 = io_outValid_39 & _T_72427; // @[Switch.scala 41:38:@33587.4]
  assign _T_72430 = select_40 == 6'h32; // @[Switch.scala 41:52:@33589.4]
  assign output_50_40 = io_outValid_40 & _T_72430; // @[Switch.scala 41:38:@33590.4]
  assign _T_72433 = select_41 == 6'h32; // @[Switch.scala 41:52:@33592.4]
  assign output_50_41 = io_outValid_41 & _T_72433; // @[Switch.scala 41:38:@33593.4]
  assign _T_72436 = select_42 == 6'h32; // @[Switch.scala 41:52:@33595.4]
  assign output_50_42 = io_outValid_42 & _T_72436; // @[Switch.scala 41:38:@33596.4]
  assign _T_72439 = select_43 == 6'h32; // @[Switch.scala 41:52:@33598.4]
  assign output_50_43 = io_outValid_43 & _T_72439; // @[Switch.scala 41:38:@33599.4]
  assign _T_72442 = select_44 == 6'h32; // @[Switch.scala 41:52:@33601.4]
  assign output_50_44 = io_outValid_44 & _T_72442; // @[Switch.scala 41:38:@33602.4]
  assign _T_72445 = select_45 == 6'h32; // @[Switch.scala 41:52:@33604.4]
  assign output_50_45 = io_outValid_45 & _T_72445; // @[Switch.scala 41:38:@33605.4]
  assign _T_72448 = select_46 == 6'h32; // @[Switch.scala 41:52:@33607.4]
  assign output_50_46 = io_outValid_46 & _T_72448; // @[Switch.scala 41:38:@33608.4]
  assign _T_72451 = select_47 == 6'h32; // @[Switch.scala 41:52:@33610.4]
  assign output_50_47 = io_outValid_47 & _T_72451; // @[Switch.scala 41:38:@33611.4]
  assign _T_72454 = select_48 == 6'h32; // @[Switch.scala 41:52:@33613.4]
  assign output_50_48 = io_outValid_48 & _T_72454; // @[Switch.scala 41:38:@33614.4]
  assign _T_72457 = select_49 == 6'h32; // @[Switch.scala 41:52:@33616.4]
  assign output_50_49 = io_outValid_49 & _T_72457; // @[Switch.scala 41:38:@33617.4]
  assign _T_72460 = select_50 == 6'h32; // @[Switch.scala 41:52:@33619.4]
  assign output_50_50 = io_outValid_50 & _T_72460; // @[Switch.scala 41:38:@33620.4]
  assign _T_72463 = select_51 == 6'h32; // @[Switch.scala 41:52:@33622.4]
  assign output_50_51 = io_outValid_51 & _T_72463; // @[Switch.scala 41:38:@33623.4]
  assign _T_72466 = select_52 == 6'h32; // @[Switch.scala 41:52:@33625.4]
  assign output_50_52 = io_outValid_52 & _T_72466; // @[Switch.scala 41:38:@33626.4]
  assign _T_72469 = select_53 == 6'h32; // @[Switch.scala 41:52:@33628.4]
  assign output_50_53 = io_outValid_53 & _T_72469; // @[Switch.scala 41:38:@33629.4]
  assign _T_72472 = select_54 == 6'h32; // @[Switch.scala 41:52:@33631.4]
  assign output_50_54 = io_outValid_54 & _T_72472; // @[Switch.scala 41:38:@33632.4]
  assign _T_72475 = select_55 == 6'h32; // @[Switch.scala 41:52:@33634.4]
  assign output_50_55 = io_outValid_55 & _T_72475; // @[Switch.scala 41:38:@33635.4]
  assign _T_72478 = select_56 == 6'h32; // @[Switch.scala 41:52:@33637.4]
  assign output_50_56 = io_outValid_56 & _T_72478; // @[Switch.scala 41:38:@33638.4]
  assign _T_72481 = select_57 == 6'h32; // @[Switch.scala 41:52:@33640.4]
  assign output_50_57 = io_outValid_57 & _T_72481; // @[Switch.scala 41:38:@33641.4]
  assign _T_72484 = select_58 == 6'h32; // @[Switch.scala 41:52:@33643.4]
  assign output_50_58 = io_outValid_58 & _T_72484; // @[Switch.scala 41:38:@33644.4]
  assign _T_72487 = select_59 == 6'h32; // @[Switch.scala 41:52:@33646.4]
  assign output_50_59 = io_outValid_59 & _T_72487; // @[Switch.scala 41:38:@33647.4]
  assign _T_72490 = select_60 == 6'h32; // @[Switch.scala 41:52:@33649.4]
  assign output_50_60 = io_outValid_60 & _T_72490; // @[Switch.scala 41:38:@33650.4]
  assign _T_72493 = select_61 == 6'h32; // @[Switch.scala 41:52:@33652.4]
  assign output_50_61 = io_outValid_61 & _T_72493; // @[Switch.scala 41:38:@33653.4]
  assign _T_72496 = select_62 == 6'h32; // @[Switch.scala 41:52:@33655.4]
  assign output_50_62 = io_outValid_62 & _T_72496; // @[Switch.scala 41:38:@33656.4]
  assign _T_72499 = select_63 == 6'h32; // @[Switch.scala 41:52:@33658.4]
  assign output_50_63 = io_outValid_63 & _T_72499; // @[Switch.scala 41:38:@33659.4]
  assign _T_72507 = {output_50_7,output_50_6,output_50_5,output_50_4,output_50_3,output_50_2,output_50_1,output_50_0}; // @[Switch.scala 43:31:@33667.4]
  assign _T_72515 = {output_50_15,output_50_14,output_50_13,output_50_12,output_50_11,output_50_10,output_50_9,output_50_8,_T_72507}; // @[Switch.scala 43:31:@33675.4]
  assign _T_72522 = {output_50_23,output_50_22,output_50_21,output_50_20,output_50_19,output_50_18,output_50_17,output_50_16}; // @[Switch.scala 43:31:@33682.4]
  assign _T_72531 = {output_50_31,output_50_30,output_50_29,output_50_28,output_50_27,output_50_26,output_50_25,output_50_24,_T_72522,_T_72515}; // @[Switch.scala 43:31:@33691.4]
  assign _T_72538 = {output_50_39,output_50_38,output_50_37,output_50_36,output_50_35,output_50_34,output_50_33,output_50_32}; // @[Switch.scala 43:31:@33698.4]
  assign _T_72546 = {output_50_47,output_50_46,output_50_45,output_50_44,output_50_43,output_50_42,output_50_41,output_50_40,_T_72538}; // @[Switch.scala 43:31:@33706.4]
  assign _T_72553 = {output_50_55,output_50_54,output_50_53,output_50_52,output_50_51,output_50_50,output_50_49,output_50_48}; // @[Switch.scala 43:31:@33713.4]
  assign _T_72562 = {output_50_63,output_50_62,output_50_61,output_50_60,output_50_59,output_50_58,output_50_57,output_50_56,_T_72553,_T_72546}; // @[Switch.scala 43:31:@33722.4]
  assign _T_72563 = {_T_72562,_T_72531}; // @[Switch.scala 43:31:@33723.4]
  assign _T_72567 = select_0 == 6'h33; // @[Switch.scala 41:52:@33726.4]
  assign output_51_0 = io_outValid_0 & _T_72567; // @[Switch.scala 41:38:@33727.4]
  assign _T_72570 = select_1 == 6'h33; // @[Switch.scala 41:52:@33729.4]
  assign output_51_1 = io_outValid_1 & _T_72570; // @[Switch.scala 41:38:@33730.4]
  assign _T_72573 = select_2 == 6'h33; // @[Switch.scala 41:52:@33732.4]
  assign output_51_2 = io_outValid_2 & _T_72573; // @[Switch.scala 41:38:@33733.4]
  assign _T_72576 = select_3 == 6'h33; // @[Switch.scala 41:52:@33735.4]
  assign output_51_3 = io_outValid_3 & _T_72576; // @[Switch.scala 41:38:@33736.4]
  assign _T_72579 = select_4 == 6'h33; // @[Switch.scala 41:52:@33738.4]
  assign output_51_4 = io_outValid_4 & _T_72579; // @[Switch.scala 41:38:@33739.4]
  assign _T_72582 = select_5 == 6'h33; // @[Switch.scala 41:52:@33741.4]
  assign output_51_5 = io_outValid_5 & _T_72582; // @[Switch.scala 41:38:@33742.4]
  assign _T_72585 = select_6 == 6'h33; // @[Switch.scala 41:52:@33744.4]
  assign output_51_6 = io_outValid_6 & _T_72585; // @[Switch.scala 41:38:@33745.4]
  assign _T_72588 = select_7 == 6'h33; // @[Switch.scala 41:52:@33747.4]
  assign output_51_7 = io_outValid_7 & _T_72588; // @[Switch.scala 41:38:@33748.4]
  assign _T_72591 = select_8 == 6'h33; // @[Switch.scala 41:52:@33750.4]
  assign output_51_8 = io_outValid_8 & _T_72591; // @[Switch.scala 41:38:@33751.4]
  assign _T_72594 = select_9 == 6'h33; // @[Switch.scala 41:52:@33753.4]
  assign output_51_9 = io_outValid_9 & _T_72594; // @[Switch.scala 41:38:@33754.4]
  assign _T_72597 = select_10 == 6'h33; // @[Switch.scala 41:52:@33756.4]
  assign output_51_10 = io_outValid_10 & _T_72597; // @[Switch.scala 41:38:@33757.4]
  assign _T_72600 = select_11 == 6'h33; // @[Switch.scala 41:52:@33759.4]
  assign output_51_11 = io_outValid_11 & _T_72600; // @[Switch.scala 41:38:@33760.4]
  assign _T_72603 = select_12 == 6'h33; // @[Switch.scala 41:52:@33762.4]
  assign output_51_12 = io_outValid_12 & _T_72603; // @[Switch.scala 41:38:@33763.4]
  assign _T_72606 = select_13 == 6'h33; // @[Switch.scala 41:52:@33765.4]
  assign output_51_13 = io_outValid_13 & _T_72606; // @[Switch.scala 41:38:@33766.4]
  assign _T_72609 = select_14 == 6'h33; // @[Switch.scala 41:52:@33768.4]
  assign output_51_14 = io_outValid_14 & _T_72609; // @[Switch.scala 41:38:@33769.4]
  assign _T_72612 = select_15 == 6'h33; // @[Switch.scala 41:52:@33771.4]
  assign output_51_15 = io_outValid_15 & _T_72612; // @[Switch.scala 41:38:@33772.4]
  assign _T_72615 = select_16 == 6'h33; // @[Switch.scala 41:52:@33774.4]
  assign output_51_16 = io_outValid_16 & _T_72615; // @[Switch.scala 41:38:@33775.4]
  assign _T_72618 = select_17 == 6'h33; // @[Switch.scala 41:52:@33777.4]
  assign output_51_17 = io_outValid_17 & _T_72618; // @[Switch.scala 41:38:@33778.4]
  assign _T_72621 = select_18 == 6'h33; // @[Switch.scala 41:52:@33780.4]
  assign output_51_18 = io_outValid_18 & _T_72621; // @[Switch.scala 41:38:@33781.4]
  assign _T_72624 = select_19 == 6'h33; // @[Switch.scala 41:52:@33783.4]
  assign output_51_19 = io_outValid_19 & _T_72624; // @[Switch.scala 41:38:@33784.4]
  assign _T_72627 = select_20 == 6'h33; // @[Switch.scala 41:52:@33786.4]
  assign output_51_20 = io_outValid_20 & _T_72627; // @[Switch.scala 41:38:@33787.4]
  assign _T_72630 = select_21 == 6'h33; // @[Switch.scala 41:52:@33789.4]
  assign output_51_21 = io_outValid_21 & _T_72630; // @[Switch.scala 41:38:@33790.4]
  assign _T_72633 = select_22 == 6'h33; // @[Switch.scala 41:52:@33792.4]
  assign output_51_22 = io_outValid_22 & _T_72633; // @[Switch.scala 41:38:@33793.4]
  assign _T_72636 = select_23 == 6'h33; // @[Switch.scala 41:52:@33795.4]
  assign output_51_23 = io_outValid_23 & _T_72636; // @[Switch.scala 41:38:@33796.4]
  assign _T_72639 = select_24 == 6'h33; // @[Switch.scala 41:52:@33798.4]
  assign output_51_24 = io_outValid_24 & _T_72639; // @[Switch.scala 41:38:@33799.4]
  assign _T_72642 = select_25 == 6'h33; // @[Switch.scala 41:52:@33801.4]
  assign output_51_25 = io_outValid_25 & _T_72642; // @[Switch.scala 41:38:@33802.4]
  assign _T_72645 = select_26 == 6'h33; // @[Switch.scala 41:52:@33804.4]
  assign output_51_26 = io_outValid_26 & _T_72645; // @[Switch.scala 41:38:@33805.4]
  assign _T_72648 = select_27 == 6'h33; // @[Switch.scala 41:52:@33807.4]
  assign output_51_27 = io_outValid_27 & _T_72648; // @[Switch.scala 41:38:@33808.4]
  assign _T_72651 = select_28 == 6'h33; // @[Switch.scala 41:52:@33810.4]
  assign output_51_28 = io_outValid_28 & _T_72651; // @[Switch.scala 41:38:@33811.4]
  assign _T_72654 = select_29 == 6'h33; // @[Switch.scala 41:52:@33813.4]
  assign output_51_29 = io_outValid_29 & _T_72654; // @[Switch.scala 41:38:@33814.4]
  assign _T_72657 = select_30 == 6'h33; // @[Switch.scala 41:52:@33816.4]
  assign output_51_30 = io_outValid_30 & _T_72657; // @[Switch.scala 41:38:@33817.4]
  assign _T_72660 = select_31 == 6'h33; // @[Switch.scala 41:52:@33819.4]
  assign output_51_31 = io_outValid_31 & _T_72660; // @[Switch.scala 41:38:@33820.4]
  assign _T_72663 = select_32 == 6'h33; // @[Switch.scala 41:52:@33822.4]
  assign output_51_32 = io_outValid_32 & _T_72663; // @[Switch.scala 41:38:@33823.4]
  assign _T_72666 = select_33 == 6'h33; // @[Switch.scala 41:52:@33825.4]
  assign output_51_33 = io_outValid_33 & _T_72666; // @[Switch.scala 41:38:@33826.4]
  assign _T_72669 = select_34 == 6'h33; // @[Switch.scala 41:52:@33828.4]
  assign output_51_34 = io_outValid_34 & _T_72669; // @[Switch.scala 41:38:@33829.4]
  assign _T_72672 = select_35 == 6'h33; // @[Switch.scala 41:52:@33831.4]
  assign output_51_35 = io_outValid_35 & _T_72672; // @[Switch.scala 41:38:@33832.4]
  assign _T_72675 = select_36 == 6'h33; // @[Switch.scala 41:52:@33834.4]
  assign output_51_36 = io_outValid_36 & _T_72675; // @[Switch.scala 41:38:@33835.4]
  assign _T_72678 = select_37 == 6'h33; // @[Switch.scala 41:52:@33837.4]
  assign output_51_37 = io_outValid_37 & _T_72678; // @[Switch.scala 41:38:@33838.4]
  assign _T_72681 = select_38 == 6'h33; // @[Switch.scala 41:52:@33840.4]
  assign output_51_38 = io_outValid_38 & _T_72681; // @[Switch.scala 41:38:@33841.4]
  assign _T_72684 = select_39 == 6'h33; // @[Switch.scala 41:52:@33843.4]
  assign output_51_39 = io_outValid_39 & _T_72684; // @[Switch.scala 41:38:@33844.4]
  assign _T_72687 = select_40 == 6'h33; // @[Switch.scala 41:52:@33846.4]
  assign output_51_40 = io_outValid_40 & _T_72687; // @[Switch.scala 41:38:@33847.4]
  assign _T_72690 = select_41 == 6'h33; // @[Switch.scala 41:52:@33849.4]
  assign output_51_41 = io_outValid_41 & _T_72690; // @[Switch.scala 41:38:@33850.4]
  assign _T_72693 = select_42 == 6'h33; // @[Switch.scala 41:52:@33852.4]
  assign output_51_42 = io_outValid_42 & _T_72693; // @[Switch.scala 41:38:@33853.4]
  assign _T_72696 = select_43 == 6'h33; // @[Switch.scala 41:52:@33855.4]
  assign output_51_43 = io_outValid_43 & _T_72696; // @[Switch.scala 41:38:@33856.4]
  assign _T_72699 = select_44 == 6'h33; // @[Switch.scala 41:52:@33858.4]
  assign output_51_44 = io_outValid_44 & _T_72699; // @[Switch.scala 41:38:@33859.4]
  assign _T_72702 = select_45 == 6'h33; // @[Switch.scala 41:52:@33861.4]
  assign output_51_45 = io_outValid_45 & _T_72702; // @[Switch.scala 41:38:@33862.4]
  assign _T_72705 = select_46 == 6'h33; // @[Switch.scala 41:52:@33864.4]
  assign output_51_46 = io_outValid_46 & _T_72705; // @[Switch.scala 41:38:@33865.4]
  assign _T_72708 = select_47 == 6'h33; // @[Switch.scala 41:52:@33867.4]
  assign output_51_47 = io_outValid_47 & _T_72708; // @[Switch.scala 41:38:@33868.4]
  assign _T_72711 = select_48 == 6'h33; // @[Switch.scala 41:52:@33870.4]
  assign output_51_48 = io_outValid_48 & _T_72711; // @[Switch.scala 41:38:@33871.4]
  assign _T_72714 = select_49 == 6'h33; // @[Switch.scala 41:52:@33873.4]
  assign output_51_49 = io_outValid_49 & _T_72714; // @[Switch.scala 41:38:@33874.4]
  assign _T_72717 = select_50 == 6'h33; // @[Switch.scala 41:52:@33876.4]
  assign output_51_50 = io_outValid_50 & _T_72717; // @[Switch.scala 41:38:@33877.4]
  assign _T_72720 = select_51 == 6'h33; // @[Switch.scala 41:52:@33879.4]
  assign output_51_51 = io_outValid_51 & _T_72720; // @[Switch.scala 41:38:@33880.4]
  assign _T_72723 = select_52 == 6'h33; // @[Switch.scala 41:52:@33882.4]
  assign output_51_52 = io_outValid_52 & _T_72723; // @[Switch.scala 41:38:@33883.4]
  assign _T_72726 = select_53 == 6'h33; // @[Switch.scala 41:52:@33885.4]
  assign output_51_53 = io_outValid_53 & _T_72726; // @[Switch.scala 41:38:@33886.4]
  assign _T_72729 = select_54 == 6'h33; // @[Switch.scala 41:52:@33888.4]
  assign output_51_54 = io_outValid_54 & _T_72729; // @[Switch.scala 41:38:@33889.4]
  assign _T_72732 = select_55 == 6'h33; // @[Switch.scala 41:52:@33891.4]
  assign output_51_55 = io_outValid_55 & _T_72732; // @[Switch.scala 41:38:@33892.4]
  assign _T_72735 = select_56 == 6'h33; // @[Switch.scala 41:52:@33894.4]
  assign output_51_56 = io_outValid_56 & _T_72735; // @[Switch.scala 41:38:@33895.4]
  assign _T_72738 = select_57 == 6'h33; // @[Switch.scala 41:52:@33897.4]
  assign output_51_57 = io_outValid_57 & _T_72738; // @[Switch.scala 41:38:@33898.4]
  assign _T_72741 = select_58 == 6'h33; // @[Switch.scala 41:52:@33900.4]
  assign output_51_58 = io_outValid_58 & _T_72741; // @[Switch.scala 41:38:@33901.4]
  assign _T_72744 = select_59 == 6'h33; // @[Switch.scala 41:52:@33903.4]
  assign output_51_59 = io_outValid_59 & _T_72744; // @[Switch.scala 41:38:@33904.4]
  assign _T_72747 = select_60 == 6'h33; // @[Switch.scala 41:52:@33906.4]
  assign output_51_60 = io_outValid_60 & _T_72747; // @[Switch.scala 41:38:@33907.4]
  assign _T_72750 = select_61 == 6'h33; // @[Switch.scala 41:52:@33909.4]
  assign output_51_61 = io_outValid_61 & _T_72750; // @[Switch.scala 41:38:@33910.4]
  assign _T_72753 = select_62 == 6'h33; // @[Switch.scala 41:52:@33912.4]
  assign output_51_62 = io_outValid_62 & _T_72753; // @[Switch.scala 41:38:@33913.4]
  assign _T_72756 = select_63 == 6'h33; // @[Switch.scala 41:52:@33915.4]
  assign output_51_63 = io_outValid_63 & _T_72756; // @[Switch.scala 41:38:@33916.4]
  assign _T_72764 = {output_51_7,output_51_6,output_51_5,output_51_4,output_51_3,output_51_2,output_51_1,output_51_0}; // @[Switch.scala 43:31:@33924.4]
  assign _T_72772 = {output_51_15,output_51_14,output_51_13,output_51_12,output_51_11,output_51_10,output_51_9,output_51_8,_T_72764}; // @[Switch.scala 43:31:@33932.4]
  assign _T_72779 = {output_51_23,output_51_22,output_51_21,output_51_20,output_51_19,output_51_18,output_51_17,output_51_16}; // @[Switch.scala 43:31:@33939.4]
  assign _T_72788 = {output_51_31,output_51_30,output_51_29,output_51_28,output_51_27,output_51_26,output_51_25,output_51_24,_T_72779,_T_72772}; // @[Switch.scala 43:31:@33948.4]
  assign _T_72795 = {output_51_39,output_51_38,output_51_37,output_51_36,output_51_35,output_51_34,output_51_33,output_51_32}; // @[Switch.scala 43:31:@33955.4]
  assign _T_72803 = {output_51_47,output_51_46,output_51_45,output_51_44,output_51_43,output_51_42,output_51_41,output_51_40,_T_72795}; // @[Switch.scala 43:31:@33963.4]
  assign _T_72810 = {output_51_55,output_51_54,output_51_53,output_51_52,output_51_51,output_51_50,output_51_49,output_51_48}; // @[Switch.scala 43:31:@33970.4]
  assign _T_72819 = {output_51_63,output_51_62,output_51_61,output_51_60,output_51_59,output_51_58,output_51_57,output_51_56,_T_72810,_T_72803}; // @[Switch.scala 43:31:@33979.4]
  assign _T_72820 = {_T_72819,_T_72788}; // @[Switch.scala 43:31:@33980.4]
  assign _T_72824 = select_0 == 6'h34; // @[Switch.scala 41:52:@33983.4]
  assign output_52_0 = io_outValid_0 & _T_72824; // @[Switch.scala 41:38:@33984.4]
  assign _T_72827 = select_1 == 6'h34; // @[Switch.scala 41:52:@33986.4]
  assign output_52_1 = io_outValid_1 & _T_72827; // @[Switch.scala 41:38:@33987.4]
  assign _T_72830 = select_2 == 6'h34; // @[Switch.scala 41:52:@33989.4]
  assign output_52_2 = io_outValid_2 & _T_72830; // @[Switch.scala 41:38:@33990.4]
  assign _T_72833 = select_3 == 6'h34; // @[Switch.scala 41:52:@33992.4]
  assign output_52_3 = io_outValid_3 & _T_72833; // @[Switch.scala 41:38:@33993.4]
  assign _T_72836 = select_4 == 6'h34; // @[Switch.scala 41:52:@33995.4]
  assign output_52_4 = io_outValid_4 & _T_72836; // @[Switch.scala 41:38:@33996.4]
  assign _T_72839 = select_5 == 6'h34; // @[Switch.scala 41:52:@33998.4]
  assign output_52_5 = io_outValid_5 & _T_72839; // @[Switch.scala 41:38:@33999.4]
  assign _T_72842 = select_6 == 6'h34; // @[Switch.scala 41:52:@34001.4]
  assign output_52_6 = io_outValid_6 & _T_72842; // @[Switch.scala 41:38:@34002.4]
  assign _T_72845 = select_7 == 6'h34; // @[Switch.scala 41:52:@34004.4]
  assign output_52_7 = io_outValid_7 & _T_72845; // @[Switch.scala 41:38:@34005.4]
  assign _T_72848 = select_8 == 6'h34; // @[Switch.scala 41:52:@34007.4]
  assign output_52_8 = io_outValid_8 & _T_72848; // @[Switch.scala 41:38:@34008.4]
  assign _T_72851 = select_9 == 6'h34; // @[Switch.scala 41:52:@34010.4]
  assign output_52_9 = io_outValid_9 & _T_72851; // @[Switch.scala 41:38:@34011.4]
  assign _T_72854 = select_10 == 6'h34; // @[Switch.scala 41:52:@34013.4]
  assign output_52_10 = io_outValid_10 & _T_72854; // @[Switch.scala 41:38:@34014.4]
  assign _T_72857 = select_11 == 6'h34; // @[Switch.scala 41:52:@34016.4]
  assign output_52_11 = io_outValid_11 & _T_72857; // @[Switch.scala 41:38:@34017.4]
  assign _T_72860 = select_12 == 6'h34; // @[Switch.scala 41:52:@34019.4]
  assign output_52_12 = io_outValid_12 & _T_72860; // @[Switch.scala 41:38:@34020.4]
  assign _T_72863 = select_13 == 6'h34; // @[Switch.scala 41:52:@34022.4]
  assign output_52_13 = io_outValid_13 & _T_72863; // @[Switch.scala 41:38:@34023.4]
  assign _T_72866 = select_14 == 6'h34; // @[Switch.scala 41:52:@34025.4]
  assign output_52_14 = io_outValid_14 & _T_72866; // @[Switch.scala 41:38:@34026.4]
  assign _T_72869 = select_15 == 6'h34; // @[Switch.scala 41:52:@34028.4]
  assign output_52_15 = io_outValid_15 & _T_72869; // @[Switch.scala 41:38:@34029.4]
  assign _T_72872 = select_16 == 6'h34; // @[Switch.scala 41:52:@34031.4]
  assign output_52_16 = io_outValid_16 & _T_72872; // @[Switch.scala 41:38:@34032.4]
  assign _T_72875 = select_17 == 6'h34; // @[Switch.scala 41:52:@34034.4]
  assign output_52_17 = io_outValid_17 & _T_72875; // @[Switch.scala 41:38:@34035.4]
  assign _T_72878 = select_18 == 6'h34; // @[Switch.scala 41:52:@34037.4]
  assign output_52_18 = io_outValid_18 & _T_72878; // @[Switch.scala 41:38:@34038.4]
  assign _T_72881 = select_19 == 6'h34; // @[Switch.scala 41:52:@34040.4]
  assign output_52_19 = io_outValid_19 & _T_72881; // @[Switch.scala 41:38:@34041.4]
  assign _T_72884 = select_20 == 6'h34; // @[Switch.scala 41:52:@34043.4]
  assign output_52_20 = io_outValid_20 & _T_72884; // @[Switch.scala 41:38:@34044.4]
  assign _T_72887 = select_21 == 6'h34; // @[Switch.scala 41:52:@34046.4]
  assign output_52_21 = io_outValid_21 & _T_72887; // @[Switch.scala 41:38:@34047.4]
  assign _T_72890 = select_22 == 6'h34; // @[Switch.scala 41:52:@34049.4]
  assign output_52_22 = io_outValid_22 & _T_72890; // @[Switch.scala 41:38:@34050.4]
  assign _T_72893 = select_23 == 6'h34; // @[Switch.scala 41:52:@34052.4]
  assign output_52_23 = io_outValid_23 & _T_72893; // @[Switch.scala 41:38:@34053.4]
  assign _T_72896 = select_24 == 6'h34; // @[Switch.scala 41:52:@34055.4]
  assign output_52_24 = io_outValid_24 & _T_72896; // @[Switch.scala 41:38:@34056.4]
  assign _T_72899 = select_25 == 6'h34; // @[Switch.scala 41:52:@34058.4]
  assign output_52_25 = io_outValid_25 & _T_72899; // @[Switch.scala 41:38:@34059.4]
  assign _T_72902 = select_26 == 6'h34; // @[Switch.scala 41:52:@34061.4]
  assign output_52_26 = io_outValid_26 & _T_72902; // @[Switch.scala 41:38:@34062.4]
  assign _T_72905 = select_27 == 6'h34; // @[Switch.scala 41:52:@34064.4]
  assign output_52_27 = io_outValid_27 & _T_72905; // @[Switch.scala 41:38:@34065.4]
  assign _T_72908 = select_28 == 6'h34; // @[Switch.scala 41:52:@34067.4]
  assign output_52_28 = io_outValid_28 & _T_72908; // @[Switch.scala 41:38:@34068.4]
  assign _T_72911 = select_29 == 6'h34; // @[Switch.scala 41:52:@34070.4]
  assign output_52_29 = io_outValid_29 & _T_72911; // @[Switch.scala 41:38:@34071.4]
  assign _T_72914 = select_30 == 6'h34; // @[Switch.scala 41:52:@34073.4]
  assign output_52_30 = io_outValid_30 & _T_72914; // @[Switch.scala 41:38:@34074.4]
  assign _T_72917 = select_31 == 6'h34; // @[Switch.scala 41:52:@34076.4]
  assign output_52_31 = io_outValid_31 & _T_72917; // @[Switch.scala 41:38:@34077.4]
  assign _T_72920 = select_32 == 6'h34; // @[Switch.scala 41:52:@34079.4]
  assign output_52_32 = io_outValid_32 & _T_72920; // @[Switch.scala 41:38:@34080.4]
  assign _T_72923 = select_33 == 6'h34; // @[Switch.scala 41:52:@34082.4]
  assign output_52_33 = io_outValid_33 & _T_72923; // @[Switch.scala 41:38:@34083.4]
  assign _T_72926 = select_34 == 6'h34; // @[Switch.scala 41:52:@34085.4]
  assign output_52_34 = io_outValid_34 & _T_72926; // @[Switch.scala 41:38:@34086.4]
  assign _T_72929 = select_35 == 6'h34; // @[Switch.scala 41:52:@34088.4]
  assign output_52_35 = io_outValid_35 & _T_72929; // @[Switch.scala 41:38:@34089.4]
  assign _T_72932 = select_36 == 6'h34; // @[Switch.scala 41:52:@34091.4]
  assign output_52_36 = io_outValid_36 & _T_72932; // @[Switch.scala 41:38:@34092.4]
  assign _T_72935 = select_37 == 6'h34; // @[Switch.scala 41:52:@34094.4]
  assign output_52_37 = io_outValid_37 & _T_72935; // @[Switch.scala 41:38:@34095.4]
  assign _T_72938 = select_38 == 6'h34; // @[Switch.scala 41:52:@34097.4]
  assign output_52_38 = io_outValid_38 & _T_72938; // @[Switch.scala 41:38:@34098.4]
  assign _T_72941 = select_39 == 6'h34; // @[Switch.scala 41:52:@34100.4]
  assign output_52_39 = io_outValid_39 & _T_72941; // @[Switch.scala 41:38:@34101.4]
  assign _T_72944 = select_40 == 6'h34; // @[Switch.scala 41:52:@34103.4]
  assign output_52_40 = io_outValid_40 & _T_72944; // @[Switch.scala 41:38:@34104.4]
  assign _T_72947 = select_41 == 6'h34; // @[Switch.scala 41:52:@34106.4]
  assign output_52_41 = io_outValid_41 & _T_72947; // @[Switch.scala 41:38:@34107.4]
  assign _T_72950 = select_42 == 6'h34; // @[Switch.scala 41:52:@34109.4]
  assign output_52_42 = io_outValid_42 & _T_72950; // @[Switch.scala 41:38:@34110.4]
  assign _T_72953 = select_43 == 6'h34; // @[Switch.scala 41:52:@34112.4]
  assign output_52_43 = io_outValid_43 & _T_72953; // @[Switch.scala 41:38:@34113.4]
  assign _T_72956 = select_44 == 6'h34; // @[Switch.scala 41:52:@34115.4]
  assign output_52_44 = io_outValid_44 & _T_72956; // @[Switch.scala 41:38:@34116.4]
  assign _T_72959 = select_45 == 6'h34; // @[Switch.scala 41:52:@34118.4]
  assign output_52_45 = io_outValid_45 & _T_72959; // @[Switch.scala 41:38:@34119.4]
  assign _T_72962 = select_46 == 6'h34; // @[Switch.scala 41:52:@34121.4]
  assign output_52_46 = io_outValid_46 & _T_72962; // @[Switch.scala 41:38:@34122.4]
  assign _T_72965 = select_47 == 6'h34; // @[Switch.scala 41:52:@34124.4]
  assign output_52_47 = io_outValid_47 & _T_72965; // @[Switch.scala 41:38:@34125.4]
  assign _T_72968 = select_48 == 6'h34; // @[Switch.scala 41:52:@34127.4]
  assign output_52_48 = io_outValid_48 & _T_72968; // @[Switch.scala 41:38:@34128.4]
  assign _T_72971 = select_49 == 6'h34; // @[Switch.scala 41:52:@34130.4]
  assign output_52_49 = io_outValid_49 & _T_72971; // @[Switch.scala 41:38:@34131.4]
  assign _T_72974 = select_50 == 6'h34; // @[Switch.scala 41:52:@34133.4]
  assign output_52_50 = io_outValid_50 & _T_72974; // @[Switch.scala 41:38:@34134.4]
  assign _T_72977 = select_51 == 6'h34; // @[Switch.scala 41:52:@34136.4]
  assign output_52_51 = io_outValid_51 & _T_72977; // @[Switch.scala 41:38:@34137.4]
  assign _T_72980 = select_52 == 6'h34; // @[Switch.scala 41:52:@34139.4]
  assign output_52_52 = io_outValid_52 & _T_72980; // @[Switch.scala 41:38:@34140.4]
  assign _T_72983 = select_53 == 6'h34; // @[Switch.scala 41:52:@34142.4]
  assign output_52_53 = io_outValid_53 & _T_72983; // @[Switch.scala 41:38:@34143.4]
  assign _T_72986 = select_54 == 6'h34; // @[Switch.scala 41:52:@34145.4]
  assign output_52_54 = io_outValid_54 & _T_72986; // @[Switch.scala 41:38:@34146.4]
  assign _T_72989 = select_55 == 6'h34; // @[Switch.scala 41:52:@34148.4]
  assign output_52_55 = io_outValid_55 & _T_72989; // @[Switch.scala 41:38:@34149.4]
  assign _T_72992 = select_56 == 6'h34; // @[Switch.scala 41:52:@34151.4]
  assign output_52_56 = io_outValid_56 & _T_72992; // @[Switch.scala 41:38:@34152.4]
  assign _T_72995 = select_57 == 6'h34; // @[Switch.scala 41:52:@34154.4]
  assign output_52_57 = io_outValid_57 & _T_72995; // @[Switch.scala 41:38:@34155.4]
  assign _T_72998 = select_58 == 6'h34; // @[Switch.scala 41:52:@34157.4]
  assign output_52_58 = io_outValid_58 & _T_72998; // @[Switch.scala 41:38:@34158.4]
  assign _T_73001 = select_59 == 6'h34; // @[Switch.scala 41:52:@34160.4]
  assign output_52_59 = io_outValid_59 & _T_73001; // @[Switch.scala 41:38:@34161.4]
  assign _T_73004 = select_60 == 6'h34; // @[Switch.scala 41:52:@34163.4]
  assign output_52_60 = io_outValid_60 & _T_73004; // @[Switch.scala 41:38:@34164.4]
  assign _T_73007 = select_61 == 6'h34; // @[Switch.scala 41:52:@34166.4]
  assign output_52_61 = io_outValid_61 & _T_73007; // @[Switch.scala 41:38:@34167.4]
  assign _T_73010 = select_62 == 6'h34; // @[Switch.scala 41:52:@34169.4]
  assign output_52_62 = io_outValid_62 & _T_73010; // @[Switch.scala 41:38:@34170.4]
  assign _T_73013 = select_63 == 6'h34; // @[Switch.scala 41:52:@34172.4]
  assign output_52_63 = io_outValid_63 & _T_73013; // @[Switch.scala 41:38:@34173.4]
  assign _T_73021 = {output_52_7,output_52_6,output_52_5,output_52_4,output_52_3,output_52_2,output_52_1,output_52_0}; // @[Switch.scala 43:31:@34181.4]
  assign _T_73029 = {output_52_15,output_52_14,output_52_13,output_52_12,output_52_11,output_52_10,output_52_9,output_52_8,_T_73021}; // @[Switch.scala 43:31:@34189.4]
  assign _T_73036 = {output_52_23,output_52_22,output_52_21,output_52_20,output_52_19,output_52_18,output_52_17,output_52_16}; // @[Switch.scala 43:31:@34196.4]
  assign _T_73045 = {output_52_31,output_52_30,output_52_29,output_52_28,output_52_27,output_52_26,output_52_25,output_52_24,_T_73036,_T_73029}; // @[Switch.scala 43:31:@34205.4]
  assign _T_73052 = {output_52_39,output_52_38,output_52_37,output_52_36,output_52_35,output_52_34,output_52_33,output_52_32}; // @[Switch.scala 43:31:@34212.4]
  assign _T_73060 = {output_52_47,output_52_46,output_52_45,output_52_44,output_52_43,output_52_42,output_52_41,output_52_40,_T_73052}; // @[Switch.scala 43:31:@34220.4]
  assign _T_73067 = {output_52_55,output_52_54,output_52_53,output_52_52,output_52_51,output_52_50,output_52_49,output_52_48}; // @[Switch.scala 43:31:@34227.4]
  assign _T_73076 = {output_52_63,output_52_62,output_52_61,output_52_60,output_52_59,output_52_58,output_52_57,output_52_56,_T_73067,_T_73060}; // @[Switch.scala 43:31:@34236.4]
  assign _T_73077 = {_T_73076,_T_73045}; // @[Switch.scala 43:31:@34237.4]
  assign _T_73081 = select_0 == 6'h35; // @[Switch.scala 41:52:@34240.4]
  assign output_53_0 = io_outValid_0 & _T_73081; // @[Switch.scala 41:38:@34241.4]
  assign _T_73084 = select_1 == 6'h35; // @[Switch.scala 41:52:@34243.4]
  assign output_53_1 = io_outValid_1 & _T_73084; // @[Switch.scala 41:38:@34244.4]
  assign _T_73087 = select_2 == 6'h35; // @[Switch.scala 41:52:@34246.4]
  assign output_53_2 = io_outValid_2 & _T_73087; // @[Switch.scala 41:38:@34247.4]
  assign _T_73090 = select_3 == 6'h35; // @[Switch.scala 41:52:@34249.4]
  assign output_53_3 = io_outValid_3 & _T_73090; // @[Switch.scala 41:38:@34250.4]
  assign _T_73093 = select_4 == 6'h35; // @[Switch.scala 41:52:@34252.4]
  assign output_53_4 = io_outValid_4 & _T_73093; // @[Switch.scala 41:38:@34253.4]
  assign _T_73096 = select_5 == 6'h35; // @[Switch.scala 41:52:@34255.4]
  assign output_53_5 = io_outValid_5 & _T_73096; // @[Switch.scala 41:38:@34256.4]
  assign _T_73099 = select_6 == 6'h35; // @[Switch.scala 41:52:@34258.4]
  assign output_53_6 = io_outValid_6 & _T_73099; // @[Switch.scala 41:38:@34259.4]
  assign _T_73102 = select_7 == 6'h35; // @[Switch.scala 41:52:@34261.4]
  assign output_53_7 = io_outValid_7 & _T_73102; // @[Switch.scala 41:38:@34262.4]
  assign _T_73105 = select_8 == 6'h35; // @[Switch.scala 41:52:@34264.4]
  assign output_53_8 = io_outValid_8 & _T_73105; // @[Switch.scala 41:38:@34265.4]
  assign _T_73108 = select_9 == 6'h35; // @[Switch.scala 41:52:@34267.4]
  assign output_53_9 = io_outValid_9 & _T_73108; // @[Switch.scala 41:38:@34268.4]
  assign _T_73111 = select_10 == 6'h35; // @[Switch.scala 41:52:@34270.4]
  assign output_53_10 = io_outValid_10 & _T_73111; // @[Switch.scala 41:38:@34271.4]
  assign _T_73114 = select_11 == 6'h35; // @[Switch.scala 41:52:@34273.4]
  assign output_53_11 = io_outValid_11 & _T_73114; // @[Switch.scala 41:38:@34274.4]
  assign _T_73117 = select_12 == 6'h35; // @[Switch.scala 41:52:@34276.4]
  assign output_53_12 = io_outValid_12 & _T_73117; // @[Switch.scala 41:38:@34277.4]
  assign _T_73120 = select_13 == 6'h35; // @[Switch.scala 41:52:@34279.4]
  assign output_53_13 = io_outValid_13 & _T_73120; // @[Switch.scala 41:38:@34280.4]
  assign _T_73123 = select_14 == 6'h35; // @[Switch.scala 41:52:@34282.4]
  assign output_53_14 = io_outValid_14 & _T_73123; // @[Switch.scala 41:38:@34283.4]
  assign _T_73126 = select_15 == 6'h35; // @[Switch.scala 41:52:@34285.4]
  assign output_53_15 = io_outValid_15 & _T_73126; // @[Switch.scala 41:38:@34286.4]
  assign _T_73129 = select_16 == 6'h35; // @[Switch.scala 41:52:@34288.4]
  assign output_53_16 = io_outValid_16 & _T_73129; // @[Switch.scala 41:38:@34289.4]
  assign _T_73132 = select_17 == 6'h35; // @[Switch.scala 41:52:@34291.4]
  assign output_53_17 = io_outValid_17 & _T_73132; // @[Switch.scala 41:38:@34292.4]
  assign _T_73135 = select_18 == 6'h35; // @[Switch.scala 41:52:@34294.4]
  assign output_53_18 = io_outValid_18 & _T_73135; // @[Switch.scala 41:38:@34295.4]
  assign _T_73138 = select_19 == 6'h35; // @[Switch.scala 41:52:@34297.4]
  assign output_53_19 = io_outValid_19 & _T_73138; // @[Switch.scala 41:38:@34298.4]
  assign _T_73141 = select_20 == 6'h35; // @[Switch.scala 41:52:@34300.4]
  assign output_53_20 = io_outValid_20 & _T_73141; // @[Switch.scala 41:38:@34301.4]
  assign _T_73144 = select_21 == 6'h35; // @[Switch.scala 41:52:@34303.4]
  assign output_53_21 = io_outValid_21 & _T_73144; // @[Switch.scala 41:38:@34304.4]
  assign _T_73147 = select_22 == 6'h35; // @[Switch.scala 41:52:@34306.4]
  assign output_53_22 = io_outValid_22 & _T_73147; // @[Switch.scala 41:38:@34307.4]
  assign _T_73150 = select_23 == 6'h35; // @[Switch.scala 41:52:@34309.4]
  assign output_53_23 = io_outValid_23 & _T_73150; // @[Switch.scala 41:38:@34310.4]
  assign _T_73153 = select_24 == 6'h35; // @[Switch.scala 41:52:@34312.4]
  assign output_53_24 = io_outValid_24 & _T_73153; // @[Switch.scala 41:38:@34313.4]
  assign _T_73156 = select_25 == 6'h35; // @[Switch.scala 41:52:@34315.4]
  assign output_53_25 = io_outValid_25 & _T_73156; // @[Switch.scala 41:38:@34316.4]
  assign _T_73159 = select_26 == 6'h35; // @[Switch.scala 41:52:@34318.4]
  assign output_53_26 = io_outValid_26 & _T_73159; // @[Switch.scala 41:38:@34319.4]
  assign _T_73162 = select_27 == 6'h35; // @[Switch.scala 41:52:@34321.4]
  assign output_53_27 = io_outValid_27 & _T_73162; // @[Switch.scala 41:38:@34322.4]
  assign _T_73165 = select_28 == 6'h35; // @[Switch.scala 41:52:@34324.4]
  assign output_53_28 = io_outValid_28 & _T_73165; // @[Switch.scala 41:38:@34325.4]
  assign _T_73168 = select_29 == 6'h35; // @[Switch.scala 41:52:@34327.4]
  assign output_53_29 = io_outValid_29 & _T_73168; // @[Switch.scala 41:38:@34328.4]
  assign _T_73171 = select_30 == 6'h35; // @[Switch.scala 41:52:@34330.4]
  assign output_53_30 = io_outValid_30 & _T_73171; // @[Switch.scala 41:38:@34331.4]
  assign _T_73174 = select_31 == 6'h35; // @[Switch.scala 41:52:@34333.4]
  assign output_53_31 = io_outValid_31 & _T_73174; // @[Switch.scala 41:38:@34334.4]
  assign _T_73177 = select_32 == 6'h35; // @[Switch.scala 41:52:@34336.4]
  assign output_53_32 = io_outValid_32 & _T_73177; // @[Switch.scala 41:38:@34337.4]
  assign _T_73180 = select_33 == 6'h35; // @[Switch.scala 41:52:@34339.4]
  assign output_53_33 = io_outValid_33 & _T_73180; // @[Switch.scala 41:38:@34340.4]
  assign _T_73183 = select_34 == 6'h35; // @[Switch.scala 41:52:@34342.4]
  assign output_53_34 = io_outValid_34 & _T_73183; // @[Switch.scala 41:38:@34343.4]
  assign _T_73186 = select_35 == 6'h35; // @[Switch.scala 41:52:@34345.4]
  assign output_53_35 = io_outValid_35 & _T_73186; // @[Switch.scala 41:38:@34346.4]
  assign _T_73189 = select_36 == 6'h35; // @[Switch.scala 41:52:@34348.4]
  assign output_53_36 = io_outValid_36 & _T_73189; // @[Switch.scala 41:38:@34349.4]
  assign _T_73192 = select_37 == 6'h35; // @[Switch.scala 41:52:@34351.4]
  assign output_53_37 = io_outValid_37 & _T_73192; // @[Switch.scala 41:38:@34352.4]
  assign _T_73195 = select_38 == 6'h35; // @[Switch.scala 41:52:@34354.4]
  assign output_53_38 = io_outValid_38 & _T_73195; // @[Switch.scala 41:38:@34355.4]
  assign _T_73198 = select_39 == 6'h35; // @[Switch.scala 41:52:@34357.4]
  assign output_53_39 = io_outValid_39 & _T_73198; // @[Switch.scala 41:38:@34358.4]
  assign _T_73201 = select_40 == 6'h35; // @[Switch.scala 41:52:@34360.4]
  assign output_53_40 = io_outValid_40 & _T_73201; // @[Switch.scala 41:38:@34361.4]
  assign _T_73204 = select_41 == 6'h35; // @[Switch.scala 41:52:@34363.4]
  assign output_53_41 = io_outValid_41 & _T_73204; // @[Switch.scala 41:38:@34364.4]
  assign _T_73207 = select_42 == 6'h35; // @[Switch.scala 41:52:@34366.4]
  assign output_53_42 = io_outValid_42 & _T_73207; // @[Switch.scala 41:38:@34367.4]
  assign _T_73210 = select_43 == 6'h35; // @[Switch.scala 41:52:@34369.4]
  assign output_53_43 = io_outValid_43 & _T_73210; // @[Switch.scala 41:38:@34370.4]
  assign _T_73213 = select_44 == 6'h35; // @[Switch.scala 41:52:@34372.4]
  assign output_53_44 = io_outValid_44 & _T_73213; // @[Switch.scala 41:38:@34373.4]
  assign _T_73216 = select_45 == 6'h35; // @[Switch.scala 41:52:@34375.4]
  assign output_53_45 = io_outValid_45 & _T_73216; // @[Switch.scala 41:38:@34376.4]
  assign _T_73219 = select_46 == 6'h35; // @[Switch.scala 41:52:@34378.4]
  assign output_53_46 = io_outValid_46 & _T_73219; // @[Switch.scala 41:38:@34379.4]
  assign _T_73222 = select_47 == 6'h35; // @[Switch.scala 41:52:@34381.4]
  assign output_53_47 = io_outValid_47 & _T_73222; // @[Switch.scala 41:38:@34382.4]
  assign _T_73225 = select_48 == 6'h35; // @[Switch.scala 41:52:@34384.4]
  assign output_53_48 = io_outValid_48 & _T_73225; // @[Switch.scala 41:38:@34385.4]
  assign _T_73228 = select_49 == 6'h35; // @[Switch.scala 41:52:@34387.4]
  assign output_53_49 = io_outValid_49 & _T_73228; // @[Switch.scala 41:38:@34388.4]
  assign _T_73231 = select_50 == 6'h35; // @[Switch.scala 41:52:@34390.4]
  assign output_53_50 = io_outValid_50 & _T_73231; // @[Switch.scala 41:38:@34391.4]
  assign _T_73234 = select_51 == 6'h35; // @[Switch.scala 41:52:@34393.4]
  assign output_53_51 = io_outValid_51 & _T_73234; // @[Switch.scala 41:38:@34394.4]
  assign _T_73237 = select_52 == 6'h35; // @[Switch.scala 41:52:@34396.4]
  assign output_53_52 = io_outValid_52 & _T_73237; // @[Switch.scala 41:38:@34397.4]
  assign _T_73240 = select_53 == 6'h35; // @[Switch.scala 41:52:@34399.4]
  assign output_53_53 = io_outValid_53 & _T_73240; // @[Switch.scala 41:38:@34400.4]
  assign _T_73243 = select_54 == 6'h35; // @[Switch.scala 41:52:@34402.4]
  assign output_53_54 = io_outValid_54 & _T_73243; // @[Switch.scala 41:38:@34403.4]
  assign _T_73246 = select_55 == 6'h35; // @[Switch.scala 41:52:@34405.4]
  assign output_53_55 = io_outValid_55 & _T_73246; // @[Switch.scala 41:38:@34406.4]
  assign _T_73249 = select_56 == 6'h35; // @[Switch.scala 41:52:@34408.4]
  assign output_53_56 = io_outValid_56 & _T_73249; // @[Switch.scala 41:38:@34409.4]
  assign _T_73252 = select_57 == 6'h35; // @[Switch.scala 41:52:@34411.4]
  assign output_53_57 = io_outValid_57 & _T_73252; // @[Switch.scala 41:38:@34412.4]
  assign _T_73255 = select_58 == 6'h35; // @[Switch.scala 41:52:@34414.4]
  assign output_53_58 = io_outValid_58 & _T_73255; // @[Switch.scala 41:38:@34415.4]
  assign _T_73258 = select_59 == 6'h35; // @[Switch.scala 41:52:@34417.4]
  assign output_53_59 = io_outValid_59 & _T_73258; // @[Switch.scala 41:38:@34418.4]
  assign _T_73261 = select_60 == 6'h35; // @[Switch.scala 41:52:@34420.4]
  assign output_53_60 = io_outValid_60 & _T_73261; // @[Switch.scala 41:38:@34421.4]
  assign _T_73264 = select_61 == 6'h35; // @[Switch.scala 41:52:@34423.4]
  assign output_53_61 = io_outValid_61 & _T_73264; // @[Switch.scala 41:38:@34424.4]
  assign _T_73267 = select_62 == 6'h35; // @[Switch.scala 41:52:@34426.4]
  assign output_53_62 = io_outValid_62 & _T_73267; // @[Switch.scala 41:38:@34427.4]
  assign _T_73270 = select_63 == 6'h35; // @[Switch.scala 41:52:@34429.4]
  assign output_53_63 = io_outValid_63 & _T_73270; // @[Switch.scala 41:38:@34430.4]
  assign _T_73278 = {output_53_7,output_53_6,output_53_5,output_53_4,output_53_3,output_53_2,output_53_1,output_53_0}; // @[Switch.scala 43:31:@34438.4]
  assign _T_73286 = {output_53_15,output_53_14,output_53_13,output_53_12,output_53_11,output_53_10,output_53_9,output_53_8,_T_73278}; // @[Switch.scala 43:31:@34446.4]
  assign _T_73293 = {output_53_23,output_53_22,output_53_21,output_53_20,output_53_19,output_53_18,output_53_17,output_53_16}; // @[Switch.scala 43:31:@34453.4]
  assign _T_73302 = {output_53_31,output_53_30,output_53_29,output_53_28,output_53_27,output_53_26,output_53_25,output_53_24,_T_73293,_T_73286}; // @[Switch.scala 43:31:@34462.4]
  assign _T_73309 = {output_53_39,output_53_38,output_53_37,output_53_36,output_53_35,output_53_34,output_53_33,output_53_32}; // @[Switch.scala 43:31:@34469.4]
  assign _T_73317 = {output_53_47,output_53_46,output_53_45,output_53_44,output_53_43,output_53_42,output_53_41,output_53_40,_T_73309}; // @[Switch.scala 43:31:@34477.4]
  assign _T_73324 = {output_53_55,output_53_54,output_53_53,output_53_52,output_53_51,output_53_50,output_53_49,output_53_48}; // @[Switch.scala 43:31:@34484.4]
  assign _T_73333 = {output_53_63,output_53_62,output_53_61,output_53_60,output_53_59,output_53_58,output_53_57,output_53_56,_T_73324,_T_73317}; // @[Switch.scala 43:31:@34493.4]
  assign _T_73334 = {_T_73333,_T_73302}; // @[Switch.scala 43:31:@34494.4]
  assign _T_73338 = select_0 == 6'h36; // @[Switch.scala 41:52:@34497.4]
  assign output_54_0 = io_outValid_0 & _T_73338; // @[Switch.scala 41:38:@34498.4]
  assign _T_73341 = select_1 == 6'h36; // @[Switch.scala 41:52:@34500.4]
  assign output_54_1 = io_outValid_1 & _T_73341; // @[Switch.scala 41:38:@34501.4]
  assign _T_73344 = select_2 == 6'h36; // @[Switch.scala 41:52:@34503.4]
  assign output_54_2 = io_outValid_2 & _T_73344; // @[Switch.scala 41:38:@34504.4]
  assign _T_73347 = select_3 == 6'h36; // @[Switch.scala 41:52:@34506.4]
  assign output_54_3 = io_outValid_3 & _T_73347; // @[Switch.scala 41:38:@34507.4]
  assign _T_73350 = select_4 == 6'h36; // @[Switch.scala 41:52:@34509.4]
  assign output_54_4 = io_outValid_4 & _T_73350; // @[Switch.scala 41:38:@34510.4]
  assign _T_73353 = select_5 == 6'h36; // @[Switch.scala 41:52:@34512.4]
  assign output_54_5 = io_outValid_5 & _T_73353; // @[Switch.scala 41:38:@34513.4]
  assign _T_73356 = select_6 == 6'h36; // @[Switch.scala 41:52:@34515.4]
  assign output_54_6 = io_outValid_6 & _T_73356; // @[Switch.scala 41:38:@34516.4]
  assign _T_73359 = select_7 == 6'h36; // @[Switch.scala 41:52:@34518.4]
  assign output_54_7 = io_outValid_7 & _T_73359; // @[Switch.scala 41:38:@34519.4]
  assign _T_73362 = select_8 == 6'h36; // @[Switch.scala 41:52:@34521.4]
  assign output_54_8 = io_outValid_8 & _T_73362; // @[Switch.scala 41:38:@34522.4]
  assign _T_73365 = select_9 == 6'h36; // @[Switch.scala 41:52:@34524.4]
  assign output_54_9 = io_outValid_9 & _T_73365; // @[Switch.scala 41:38:@34525.4]
  assign _T_73368 = select_10 == 6'h36; // @[Switch.scala 41:52:@34527.4]
  assign output_54_10 = io_outValid_10 & _T_73368; // @[Switch.scala 41:38:@34528.4]
  assign _T_73371 = select_11 == 6'h36; // @[Switch.scala 41:52:@34530.4]
  assign output_54_11 = io_outValid_11 & _T_73371; // @[Switch.scala 41:38:@34531.4]
  assign _T_73374 = select_12 == 6'h36; // @[Switch.scala 41:52:@34533.4]
  assign output_54_12 = io_outValid_12 & _T_73374; // @[Switch.scala 41:38:@34534.4]
  assign _T_73377 = select_13 == 6'h36; // @[Switch.scala 41:52:@34536.4]
  assign output_54_13 = io_outValid_13 & _T_73377; // @[Switch.scala 41:38:@34537.4]
  assign _T_73380 = select_14 == 6'h36; // @[Switch.scala 41:52:@34539.4]
  assign output_54_14 = io_outValid_14 & _T_73380; // @[Switch.scala 41:38:@34540.4]
  assign _T_73383 = select_15 == 6'h36; // @[Switch.scala 41:52:@34542.4]
  assign output_54_15 = io_outValid_15 & _T_73383; // @[Switch.scala 41:38:@34543.4]
  assign _T_73386 = select_16 == 6'h36; // @[Switch.scala 41:52:@34545.4]
  assign output_54_16 = io_outValid_16 & _T_73386; // @[Switch.scala 41:38:@34546.4]
  assign _T_73389 = select_17 == 6'h36; // @[Switch.scala 41:52:@34548.4]
  assign output_54_17 = io_outValid_17 & _T_73389; // @[Switch.scala 41:38:@34549.4]
  assign _T_73392 = select_18 == 6'h36; // @[Switch.scala 41:52:@34551.4]
  assign output_54_18 = io_outValid_18 & _T_73392; // @[Switch.scala 41:38:@34552.4]
  assign _T_73395 = select_19 == 6'h36; // @[Switch.scala 41:52:@34554.4]
  assign output_54_19 = io_outValid_19 & _T_73395; // @[Switch.scala 41:38:@34555.4]
  assign _T_73398 = select_20 == 6'h36; // @[Switch.scala 41:52:@34557.4]
  assign output_54_20 = io_outValid_20 & _T_73398; // @[Switch.scala 41:38:@34558.4]
  assign _T_73401 = select_21 == 6'h36; // @[Switch.scala 41:52:@34560.4]
  assign output_54_21 = io_outValid_21 & _T_73401; // @[Switch.scala 41:38:@34561.4]
  assign _T_73404 = select_22 == 6'h36; // @[Switch.scala 41:52:@34563.4]
  assign output_54_22 = io_outValid_22 & _T_73404; // @[Switch.scala 41:38:@34564.4]
  assign _T_73407 = select_23 == 6'h36; // @[Switch.scala 41:52:@34566.4]
  assign output_54_23 = io_outValid_23 & _T_73407; // @[Switch.scala 41:38:@34567.4]
  assign _T_73410 = select_24 == 6'h36; // @[Switch.scala 41:52:@34569.4]
  assign output_54_24 = io_outValid_24 & _T_73410; // @[Switch.scala 41:38:@34570.4]
  assign _T_73413 = select_25 == 6'h36; // @[Switch.scala 41:52:@34572.4]
  assign output_54_25 = io_outValid_25 & _T_73413; // @[Switch.scala 41:38:@34573.4]
  assign _T_73416 = select_26 == 6'h36; // @[Switch.scala 41:52:@34575.4]
  assign output_54_26 = io_outValid_26 & _T_73416; // @[Switch.scala 41:38:@34576.4]
  assign _T_73419 = select_27 == 6'h36; // @[Switch.scala 41:52:@34578.4]
  assign output_54_27 = io_outValid_27 & _T_73419; // @[Switch.scala 41:38:@34579.4]
  assign _T_73422 = select_28 == 6'h36; // @[Switch.scala 41:52:@34581.4]
  assign output_54_28 = io_outValid_28 & _T_73422; // @[Switch.scala 41:38:@34582.4]
  assign _T_73425 = select_29 == 6'h36; // @[Switch.scala 41:52:@34584.4]
  assign output_54_29 = io_outValid_29 & _T_73425; // @[Switch.scala 41:38:@34585.4]
  assign _T_73428 = select_30 == 6'h36; // @[Switch.scala 41:52:@34587.4]
  assign output_54_30 = io_outValid_30 & _T_73428; // @[Switch.scala 41:38:@34588.4]
  assign _T_73431 = select_31 == 6'h36; // @[Switch.scala 41:52:@34590.4]
  assign output_54_31 = io_outValid_31 & _T_73431; // @[Switch.scala 41:38:@34591.4]
  assign _T_73434 = select_32 == 6'h36; // @[Switch.scala 41:52:@34593.4]
  assign output_54_32 = io_outValid_32 & _T_73434; // @[Switch.scala 41:38:@34594.4]
  assign _T_73437 = select_33 == 6'h36; // @[Switch.scala 41:52:@34596.4]
  assign output_54_33 = io_outValid_33 & _T_73437; // @[Switch.scala 41:38:@34597.4]
  assign _T_73440 = select_34 == 6'h36; // @[Switch.scala 41:52:@34599.4]
  assign output_54_34 = io_outValid_34 & _T_73440; // @[Switch.scala 41:38:@34600.4]
  assign _T_73443 = select_35 == 6'h36; // @[Switch.scala 41:52:@34602.4]
  assign output_54_35 = io_outValid_35 & _T_73443; // @[Switch.scala 41:38:@34603.4]
  assign _T_73446 = select_36 == 6'h36; // @[Switch.scala 41:52:@34605.4]
  assign output_54_36 = io_outValid_36 & _T_73446; // @[Switch.scala 41:38:@34606.4]
  assign _T_73449 = select_37 == 6'h36; // @[Switch.scala 41:52:@34608.4]
  assign output_54_37 = io_outValid_37 & _T_73449; // @[Switch.scala 41:38:@34609.4]
  assign _T_73452 = select_38 == 6'h36; // @[Switch.scala 41:52:@34611.4]
  assign output_54_38 = io_outValid_38 & _T_73452; // @[Switch.scala 41:38:@34612.4]
  assign _T_73455 = select_39 == 6'h36; // @[Switch.scala 41:52:@34614.4]
  assign output_54_39 = io_outValid_39 & _T_73455; // @[Switch.scala 41:38:@34615.4]
  assign _T_73458 = select_40 == 6'h36; // @[Switch.scala 41:52:@34617.4]
  assign output_54_40 = io_outValid_40 & _T_73458; // @[Switch.scala 41:38:@34618.4]
  assign _T_73461 = select_41 == 6'h36; // @[Switch.scala 41:52:@34620.4]
  assign output_54_41 = io_outValid_41 & _T_73461; // @[Switch.scala 41:38:@34621.4]
  assign _T_73464 = select_42 == 6'h36; // @[Switch.scala 41:52:@34623.4]
  assign output_54_42 = io_outValid_42 & _T_73464; // @[Switch.scala 41:38:@34624.4]
  assign _T_73467 = select_43 == 6'h36; // @[Switch.scala 41:52:@34626.4]
  assign output_54_43 = io_outValid_43 & _T_73467; // @[Switch.scala 41:38:@34627.4]
  assign _T_73470 = select_44 == 6'h36; // @[Switch.scala 41:52:@34629.4]
  assign output_54_44 = io_outValid_44 & _T_73470; // @[Switch.scala 41:38:@34630.4]
  assign _T_73473 = select_45 == 6'h36; // @[Switch.scala 41:52:@34632.4]
  assign output_54_45 = io_outValid_45 & _T_73473; // @[Switch.scala 41:38:@34633.4]
  assign _T_73476 = select_46 == 6'h36; // @[Switch.scala 41:52:@34635.4]
  assign output_54_46 = io_outValid_46 & _T_73476; // @[Switch.scala 41:38:@34636.4]
  assign _T_73479 = select_47 == 6'h36; // @[Switch.scala 41:52:@34638.4]
  assign output_54_47 = io_outValid_47 & _T_73479; // @[Switch.scala 41:38:@34639.4]
  assign _T_73482 = select_48 == 6'h36; // @[Switch.scala 41:52:@34641.4]
  assign output_54_48 = io_outValid_48 & _T_73482; // @[Switch.scala 41:38:@34642.4]
  assign _T_73485 = select_49 == 6'h36; // @[Switch.scala 41:52:@34644.4]
  assign output_54_49 = io_outValid_49 & _T_73485; // @[Switch.scala 41:38:@34645.4]
  assign _T_73488 = select_50 == 6'h36; // @[Switch.scala 41:52:@34647.4]
  assign output_54_50 = io_outValid_50 & _T_73488; // @[Switch.scala 41:38:@34648.4]
  assign _T_73491 = select_51 == 6'h36; // @[Switch.scala 41:52:@34650.4]
  assign output_54_51 = io_outValid_51 & _T_73491; // @[Switch.scala 41:38:@34651.4]
  assign _T_73494 = select_52 == 6'h36; // @[Switch.scala 41:52:@34653.4]
  assign output_54_52 = io_outValid_52 & _T_73494; // @[Switch.scala 41:38:@34654.4]
  assign _T_73497 = select_53 == 6'h36; // @[Switch.scala 41:52:@34656.4]
  assign output_54_53 = io_outValid_53 & _T_73497; // @[Switch.scala 41:38:@34657.4]
  assign _T_73500 = select_54 == 6'h36; // @[Switch.scala 41:52:@34659.4]
  assign output_54_54 = io_outValid_54 & _T_73500; // @[Switch.scala 41:38:@34660.4]
  assign _T_73503 = select_55 == 6'h36; // @[Switch.scala 41:52:@34662.4]
  assign output_54_55 = io_outValid_55 & _T_73503; // @[Switch.scala 41:38:@34663.4]
  assign _T_73506 = select_56 == 6'h36; // @[Switch.scala 41:52:@34665.4]
  assign output_54_56 = io_outValid_56 & _T_73506; // @[Switch.scala 41:38:@34666.4]
  assign _T_73509 = select_57 == 6'h36; // @[Switch.scala 41:52:@34668.4]
  assign output_54_57 = io_outValid_57 & _T_73509; // @[Switch.scala 41:38:@34669.4]
  assign _T_73512 = select_58 == 6'h36; // @[Switch.scala 41:52:@34671.4]
  assign output_54_58 = io_outValid_58 & _T_73512; // @[Switch.scala 41:38:@34672.4]
  assign _T_73515 = select_59 == 6'h36; // @[Switch.scala 41:52:@34674.4]
  assign output_54_59 = io_outValid_59 & _T_73515; // @[Switch.scala 41:38:@34675.4]
  assign _T_73518 = select_60 == 6'h36; // @[Switch.scala 41:52:@34677.4]
  assign output_54_60 = io_outValid_60 & _T_73518; // @[Switch.scala 41:38:@34678.4]
  assign _T_73521 = select_61 == 6'h36; // @[Switch.scala 41:52:@34680.4]
  assign output_54_61 = io_outValid_61 & _T_73521; // @[Switch.scala 41:38:@34681.4]
  assign _T_73524 = select_62 == 6'h36; // @[Switch.scala 41:52:@34683.4]
  assign output_54_62 = io_outValid_62 & _T_73524; // @[Switch.scala 41:38:@34684.4]
  assign _T_73527 = select_63 == 6'h36; // @[Switch.scala 41:52:@34686.4]
  assign output_54_63 = io_outValid_63 & _T_73527; // @[Switch.scala 41:38:@34687.4]
  assign _T_73535 = {output_54_7,output_54_6,output_54_5,output_54_4,output_54_3,output_54_2,output_54_1,output_54_0}; // @[Switch.scala 43:31:@34695.4]
  assign _T_73543 = {output_54_15,output_54_14,output_54_13,output_54_12,output_54_11,output_54_10,output_54_9,output_54_8,_T_73535}; // @[Switch.scala 43:31:@34703.4]
  assign _T_73550 = {output_54_23,output_54_22,output_54_21,output_54_20,output_54_19,output_54_18,output_54_17,output_54_16}; // @[Switch.scala 43:31:@34710.4]
  assign _T_73559 = {output_54_31,output_54_30,output_54_29,output_54_28,output_54_27,output_54_26,output_54_25,output_54_24,_T_73550,_T_73543}; // @[Switch.scala 43:31:@34719.4]
  assign _T_73566 = {output_54_39,output_54_38,output_54_37,output_54_36,output_54_35,output_54_34,output_54_33,output_54_32}; // @[Switch.scala 43:31:@34726.4]
  assign _T_73574 = {output_54_47,output_54_46,output_54_45,output_54_44,output_54_43,output_54_42,output_54_41,output_54_40,_T_73566}; // @[Switch.scala 43:31:@34734.4]
  assign _T_73581 = {output_54_55,output_54_54,output_54_53,output_54_52,output_54_51,output_54_50,output_54_49,output_54_48}; // @[Switch.scala 43:31:@34741.4]
  assign _T_73590 = {output_54_63,output_54_62,output_54_61,output_54_60,output_54_59,output_54_58,output_54_57,output_54_56,_T_73581,_T_73574}; // @[Switch.scala 43:31:@34750.4]
  assign _T_73591 = {_T_73590,_T_73559}; // @[Switch.scala 43:31:@34751.4]
  assign _T_73595 = select_0 == 6'h37; // @[Switch.scala 41:52:@34754.4]
  assign output_55_0 = io_outValid_0 & _T_73595; // @[Switch.scala 41:38:@34755.4]
  assign _T_73598 = select_1 == 6'h37; // @[Switch.scala 41:52:@34757.4]
  assign output_55_1 = io_outValid_1 & _T_73598; // @[Switch.scala 41:38:@34758.4]
  assign _T_73601 = select_2 == 6'h37; // @[Switch.scala 41:52:@34760.4]
  assign output_55_2 = io_outValid_2 & _T_73601; // @[Switch.scala 41:38:@34761.4]
  assign _T_73604 = select_3 == 6'h37; // @[Switch.scala 41:52:@34763.4]
  assign output_55_3 = io_outValid_3 & _T_73604; // @[Switch.scala 41:38:@34764.4]
  assign _T_73607 = select_4 == 6'h37; // @[Switch.scala 41:52:@34766.4]
  assign output_55_4 = io_outValid_4 & _T_73607; // @[Switch.scala 41:38:@34767.4]
  assign _T_73610 = select_5 == 6'h37; // @[Switch.scala 41:52:@34769.4]
  assign output_55_5 = io_outValid_5 & _T_73610; // @[Switch.scala 41:38:@34770.4]
  assign _T_73613 = select_6 == 6'h37; // @[Switch.scala 41:52:@34772.4]
  assign output_55_6 = io_outValid_6 & _T_73613; // @[Switch.scala 41:38:@34773.4]
  assign _T_73616 = select_7 == 6'h37; // @[Switch.scala 41:52:@34775.4]
  assign output_55_7 = io_outValid_7 & _T_73616; // @[Switch.scala 41:38:@34776.4]
  assign _T_73619 = select_8 == 6'h37; // @[Switch.scala 41:52:@34778.4]
  assign output_55_8 = io_outValid_8 & _T_73619; // @[Switch.scala 41:38:@34779.4]
  assign _T_73622 = select_9 == 6'h37; // @[Switch.scala 41:52:@34781.4]
  assign output_55_9 = io_outValid_9 & _T_73622; // @[Switch.scala 41:38:@34782.4]
  assign _T_73625 = select_10 == 6'h37; // @[Switch.scala 41:52:@34784.4]
  assign output_55_10 = io_outValid_10 & _T_73625; // @[Switch.scala 41:38:@34785.4]
  assign _T_73628 = select_11 == 6'h37; // @[Switch.scala 41:52:@34787.4]
  assign output_55_11 = io_outValid_11 & _T_73628; // @[Switch.scala 41:38:@34788.4]
  assign _T_73631 = select_12 == 6'h37; // @[Switch.scala 41:52:@34790.4]
  assign output_55_12 = io_outValid_12 & _T_73631; // @[Switch.scala 41:38:@34791.4]
  assign _T_73634 = select_13 == 6'h37; // @[Switch.scala 41:52:@34793.4]
  assign output_55_13 = io_outValid_13 & _T_73634; // @[Switch.scala 41:38:@34794.4]
  assign _T_73637 = select_14 == 6'h37; // @[Switch.scala 41:52:@34796.4]
  assign output_55_14 = io_outValid_14 & _T_73637; // @[Switch.scala 41:38:@34797.4]
  assign _T_73640 = select_15 == 6'h37; // @[Switch.scala 41:52:@34799.4]
  assign output_55_15 = io_outValid_15 & _T_73640; // @[Switch.scala 41:38:@34800.4]
  assign _T_73643 = select_16 == 6'h37; // @[Switch.scala 41:52:@34802.4]
  assign output_55_16 = io_outValid_16 & _T_73643; // @[Switch.scala 41:38:@34803.4]
  assign _T_73646 = select_17 == 6'h37; // @[Switch.scala 41:52:@34805.4]
  assign output_55_17 = io_outValid_17 & _T_73646; // @[Switch.scala 41:38:@34806.4]
  assign _T_73649 = select_18 == 6'h37; // @[Switch.scala 41:52:@34808.4]
  assign output_55_18 = io_outValid_18 & _T_73649; // @[Switch.scala 41:38:@34809.4]
  assign _T_73652 = select_19 == 6'h37; // @[Switch.scala 41:52:@34811.4]
  assign output_55_19 = io_outValid_19 & _T_73652; // @[Switch.scala 41:38:@34812.4]
  assign _T_73655 = select_20 == 6'h37; // @[Switch.scala 41:52:@34814.4]
  assign output_55_20 = io_outValid_20 & _T_73655; // @[Switch.scala 41:38:@34815.4]
  assign _T_73658 = select_21 == 6'h37; // @[Switch.scala 41:52:@34817.4]
  assign output_55_21 = io_outValid_21 & _T_73658; // @[Switch.scala 41:38:@34818.4]
  assign _T_73661 = select_22 == 6'h37; // @[Switch.scala 41:52:@34820.4]
  assign output_55_22 = io_outValid_22 & _T_73661; // @[Switch.scala 41:38:@34821.4]
  assign _T_73664 = select_23 == 6'h37; // @[Switch.scala 41:52:@34823.4]
  assign output_55_23 = io_outValid_23 & _T_73664; // @[Switch.scala 41:38:@34824.4]
  assign _T_73667 = select_24 == 6'h37; // @[Switch.scala 41:52:@34826.4]
  assign output_55_24 = io_outValid_24 & _T_73667; // @[Switch.scala 41:38:@34827.4]
  assign _T_73670 = select_25 == 6'h37; // @[Switch.scala 41:52:@34829.4]
  assign output_55_25 = io_outValid_25 & _T_73670; // @[Switch.scala 41:38:@34830.4]
  assign _T_73673 = select_26 == 6'h37; // @[Switch.scala 41:52:@34832.4]
  assign output_55_26 = io_outValid_26 & _T_73673; // @[Switch.scala 41:38:@34833.4]
  assign _T_73676 = select_27 == 6'h37; // @[Switch.scala 41:52:@34835.4]
  assign output_55_27 = io_outValid_27 & _T_73676; // @[Switch.scala 41:38:@34836.4]
  assign _T_73679 = select_28 == 6'h37; // @[Switch.scala 41:52:@34838.4]
  assign output_55_28 = io_outValid_28 & _T_73679; // @[Switch.scala 41:38:@34839.4]
  assign _T_73682 = select_29 == 6'h37; // @[Switch.scala 41:52:@34841.4]
  assign output_55_29 = io_outValid_29 & _T_73682; // @[Switch.scala 41:38:@34842.4]
  assign _T_73685 = select_30 == 6'h37; // @[Switch.scala 41:52:@34844.4]
  assign output_55_30 = io_outValid_30 & _T_73685; // @[Switch.scala 41:38:@34845.4]
  assign _T_73688 = select_31 == 6'h37; // @[Switch.scala 41:52:@34847.4]
  assign output_55_31 = io_outValid_31 & _T_73688; // @[Switch.scala 41:38:@34848.4]
  assign _T_73691 = select_32 == 6'h37; // @[Switch.scala 41:52:@34850.4]
  assign output_55_32 = io_outValid_32 & _T_73691; // @[Switch.scala 41:38:@34851.4]
  assign _T_73694 = select_33 == 6'h37; // @[Switch.scala 41:52:@34853.4]
  assign output_55_33 = io_outValid_33 & _T_73694; // @[Switch.scala 41:38:@34854.4]
  assign _T_73697 = select_34 == 6'h37; // @[Switch.scala 41:52:@34856.4]
  assign output_55_34 = io_outValid_34 & _T_73697; // @[Switch.scala 41:38:@34857.4]
  assign _T_73700 = select_35 == 6'h37; // @[Switch.scala 41:52:@34859.4]
  assign output_55_35 = io_outValid_35 & _T_73700; // @[Switch.scala 41:38:@34860.4]
  assign _T_73703 = select_36 == 6'h37; // @[Switch.scala 41:52:@34862.4]
  assign output_55_36 = io_outValid_36 & _T_73703; // @[Switch.scala 41:38:@34863.4]
  assign _T_73706 = select_37 == 6'h37; // @[Switch.scala 41:52:@34865.4]
  assign output_55_37 = io_outValid_37 & _T_73706; // @[Switch.scala 41:38:@34866.4]
  assign _T_73709 = select_38 == 6'h37; // @[Switch.scala 41:52:@34868.4]
  assign output_55_38 = io_outValid_38 & _T_73709; // @[Switch.scala 41:38:@34869.4]
  assign _T_73712 = select_39 == 6'h37; // @[Switch.scala 41:52:@34871.4]
  assign output_55_39 = io_outValid_39 & _T_73712; // @[Switch.scala 41:38:@34872.4]
  assign _T_73715 = select_40 == 6'h37; // @[Switch.scala 41:52:@34874.4]
  assign output_55_40 = io_outValid_40 & _T_73715; // @[Switch.scala 41:38:@34875.4]
  assign _T_73718 = select_41 == 6'h37; // @[Switch.scala 41:52:@34877.4]
  assign output_55_41 = io_outValid_41 & _T_73718; // @[Switch.scala 41:38:@34878.4]
  assign _T_73721 = select_42 == 6'h37; // @[Switch.scala 41:52:@34880.4]
  assign output_55_42 = io_outValid_42 & _T_73721; // @[Switch.scala 41:38:@34881.4]
  assign _T_73724 = select_43 == 6'h37; // @[Switch.scala 41:52:@34883.4]
  assign output_55_43 = io_outValid_43 & _T_73724; // @[Switch.scala 41:38:@34884.4]
  assign _T_73727 = select_44 == 6'h37; // @[Switch.scala 41:52:@34886.4]
  assign output_55_44 = io_outValid_44 & _T_73727; // @[Switch.scala 41:38:@34887.4]
  assign _T_73730 = select_45 == 6'h37; // @[Switch.scala 41:52:@34889.4]
  assign output_55_45 = io_outValid_45 & _T_73730; // @[Switch.scala 41:38:@34890.4]
  assign _T_73733 = select_46 == 6'h37; // @[Switch.scala 41:52:@34892.4]
  assign output_55_46 = io_outValid_46 & _T_73733; // @[Switch.scala 41:38:@34893.4]
  assign _T_73736 = select_47 == 6'h37; // @[Switch.scala 41:52:@34895.4]
  assign output_55_47 = io_outValid_47 & _T_73736; // @[Switch.scala 41:38:@34896.4]
  assign _T_73739 = select_48 == 6'h37; // @[Switch.scala 41:52:@34898.4]
  assign output_55_48 = io_outValid_48 & _T_73739; // @[Switch.scala 41:38:@34899.4]
  assign _T_73742 = select_49 == 6'h37; // @[Switch.scala 41:52:@34901.4]
  assign output_55_49 = io_outValid_49 & _T_73742; // @[Switch.scala 41:38:@34902.4]
  assign _T_73745 = select_50 == 6'h37; // @[Switch.scala 41:52:@34904.4]
  assign output_55_50 = io_outValid_50 & _T_73745; // @[Switch.scala 41:38:@34905.4]
  assign _T_73748 = select_51 == 6'h37; // @[Switch.scala 41:52:@34907.4]
  assign output_55_51 = io_outValid_51 & _T_73748; // @[Switch.scala 41:38:@34908.4]
  assign _T_73751 = select_52 == 6'h37; // @[Switch.scala 41:52:@34910.4]
  assign output_55_52 = io_outValid_52 & _T_73751; // @[Switch.scala 41:38:@34911.4]
  assign _T_73754 = select_53 == 6'h37; // @[Switch.scala 41:52:@34913.4]
  assign output_55_53 = io_outValid_53 & _T_73754; // @[Switch.scala 41:38:@34914.4]
  assign _T_73757 = select_54 == 6'h37; // @[Switch.scala 41:52:@34916.4]
  assign output_55_54 = io_outValid_54 & _T_73757; // @[Switch.scala 41:38:@34917.4]
  assign _T_73760 = select_55 == 6'h37; // @[Switch.scala 41:52:@34919.4]
  assign output_55_55 = io_outValid_55 & _T_73760; // @[Switch.scala 41:38:@34920.4]
  assign _T_73763 = select_56 == 6'h37; // @[Switch.scala 41:52:@34922.4]
  assign output_55_56 = io_outValid_56 & _T_73763; // @[Switch.scala 41:38:@34923.4]
  assign _T_73766 = select_57 == 6'h37; // @[Switch.scala 41:52:@34925.4]
  assign output_55_57 = io_outValid_57 & _T_73766; // @[Switch.scala 41:38:@34926.4]
  assign _T_73769 = select_58 == 6'h37; // @[Switch.scala 41:52:@34928.4]
  assign output_55_58 = io_outValid_58 & _T_73769; // @[Switch.scala 41:38:@34929.4]
  assign _T_73772 = select_59 == 6'h37; // @[Switch.scala 41:52:@34931.4]
  assign output_55_59 = io_outValid_59 & _T_73772; // @[Switch.scala 41:38:@34932.4]
  assign _T_73775 = select_60 == 6'h37; // @[Switch.scala 41:52:@34934.4]
  assign output_55_60 = io_outValid_60 & _T_73775; // @[Switch.scala 41:38:@34935.4]
  assign _T_73778 = select_61 == 6'h37; // @[Switch.scala 41:52:@34937.4]
  assign output_55_61 = io_outValid_61 & _T_73778; // @[Switch.scala 41:38:@34938.4]
  assign _T_73781 = select_62 == 6'h37; // @[Switch.scala 41:52:@34940.4]
  assign output_55_62 = io_outValid_62 & _T_73781; // @[Switch.scala 41:38:@34941.4]
  assign _T_73784 = select_63 == 6'h37; // @[Switch.scala 41:52:@34943.4]
  assign output_55_63 = io_outValid_63 & _T_73784; // @[Switch.scala 41:38:@34944.4]
  assign _T_73792 = {output_55_7,output_55_6,output_55_5,output_55_4,output_55_3,output_55_2,output_55_1,output_55_0}; // @[Switch.scala 43:31:@34952.4]
  assign _T_73800 = {output_55_15,output_55_14,output_55_13,output_55_12,output_55_11,output_55_10,output_55_9,output_55_8,_T_73792}; // @[Switch.scala 43:31:@34960.4]
  assign _T_73807 = {output_55_23,output_55_22,output_55_21,output_55_20,output_55_19,output_55_18,output_55_17,output_55_16}; // @[Switch.scala 43:31:@34967.4]
  assign _T_73816 = {output_55_31,output_55_30,output_55_29,output_55_28,output_55_27,output_55_26,output_55_25,output_55_24,_T_73807,_T_73800}; // @[Switch.scala 43:31:@34976.4]
  assign _T_73823 = {output_55_39,output_55_38,output_55_37,output_55_36,output_55_35,output_55_34,output_55_33,output_55_32}; // @[Switch.scala 43:31:@34983.4]
  assign _T_73831 = {output_55_47,output_55_46,output_55_45,output_55_44,output_55_43,output_55_42,output_55_41,output_55_40,_T_73823}; // @[Switch.scala 43:31:@34991.4]
  assign _T_73838 = {output_55_55,output_55_54,output_55_53,output_55_52,output_55_51,output_55_50,output_55_49,output_55_48}; // @[Switch.scala 43:31:@34998.4]
  assign _T_73847 = {output_55_63,output_55_62,output_55_61,output_55_60,output_55_59,output_55_58,output_55_57,output_55_56,_T_73838,_T_73831}; // @[Switch.scala 43:31:@35007.4]
  assign _T_73848 = {_T_73847,_T_73816}; // @[Switch.scala 43:31:@35008.4]
  assign _T_73852 = select_0 == 6'h38; // @[Switch.scala 41:52:@35011.4]
  assign output_56_0 = io_outValid_0 & _T_73852; // @[Switch.scala 41:38:@35012.4]
  assign _T_73855 = select_1 == 6'h38; // @[Switch.scala 41:52:@35014.4]
  assign output_56_1 = io_outValid_1 & _T_73855; // @[Switch.scala 41:38:@35015.4]
  assign _T_73858 = select_2 == 6'h38; // @[Switch.scala 41:52:@35017.4]
  assign output_56_2 = io_outValid_2 & _T_73858; // @[Switch.scala 41:38:@35018.4]
  assign _T_73861 = select_3 == 6'h38; // @[Switch.scala 41:52:@35020.4]
  assign output_56_3 = io_outValid_3 & _T_73861; // @[Switch.scala 41:38:@35021.4]
  assign _T_73864 = select_4 == 6'h38; // @[Switch.scala 41:52:@35023.4]
  assign output_56_4 = io_outValid_4 & _T_73864; // @[Switch.scala 41:38:@35024.4]
  assign _T_73867 = select_5 == 6'h38; // @[Switch.scala 41:52:@35026.4]
  assign output_56_5 = io_outValid_5 & _T_73867; // @[Switch.scala 41:38:@35027.4]
  assign _T_73870 = select_6 == 6'h38; // @[Switch.scala 41:52:@35029.4]
  assign output_56_6 = io_outValid_6 & _T_73870; // @[Switch.scala 41:38:@35030.4]
  assign _T_73873 = select_7 == 6'h38; // @[Switch.scala 41:52:@35032.4]
  assign output_56_7 = io_outValid_7 & _T_73873; // @[Switch.scala 41:38:@35033.4]
  assign _T_73876 = select_8 == 6'h38; // @[Switch.scala 41:52:@35035.4]
  assign output_56_8 = io_outValid_8 & _T_73876; // @[Switch.scala 41:38:@35036.4]
  assign _T_73879 = select_9 == 6'h38; // @[Switch.scala 41:52:@35038.4]
  assign output_56_9 = io_outValid_9 & _T_73879; // @[Switch.scala 41:38:@35039.4]
  assign _T_73882 = select_10 == 6'h38; // @[Switch.scala 41:52:@35041.4]
  assign output_56_10 = io_outValid_10 & _T_73882; // @[Switch.scala 41:38:@35042.4]
  assign _T_73885 = select_11 == 6'h38; // @[Switch.scala 41:52:@35044.4]
  assign output_56_11 = io_outValid_11 & _T_73885; // @[Switch.scala 41:38:@35045.4]
  assign _T_73888 = select_12 == 6'h38; // @[Switch.scala 41:52:@35047.4]
  assign output_56_12 = io_outValid_12 & _T_73888; // @[Switch.scala 41:38:@35048.4]
  assign _T_73891 = select_13 == 6'h38; // @[Switch.scala 41:52:@35050.4]
  assign output_56_13 = io_outValid_13 & _T_73891; // @[Switch.scala 41:38:@35051.4]
  assign _T_73894 = select_14 == 6'h38; // @[Switch.scala 41:52:@35053.4]
  assign output_56_14 = io_outValid_14 & _T_73894; // @[Switch.scala 41:38:@35054.4]
  assign _T_73897 = select_15 == 6'h38; // @[Switch.scala 41:52:@35056.4]
  assign output_56_15 = io_outValid_15 & _T_73897; // @[Switch.scala 41:38:@35057.4]
  assign _T_73900 = select_16 == 6'h38; // @[Switch.scala 41:52:@35059.4]
  assign output_56_16 = io_outValid_16 & _T_73900; // @[Switch.scala 41:38:@35060.4]
  assign _T_73903 = select_17 == 6'h38; // @[Switch.scala 41:52:@35062.4]
  assign output_56_17 = io_outValid_17 & _T_73903; // @[Switch.scala 41:38:@35063.4]
  assign _T_73906 = select_18 == 6'h38; // @[Switch.scala 41:52:@35065.4]
  assign output_56_18 = io_outValid_18 & _T_73906; // @[Switch.scala 41:38:@35066.4]
  assign _T_73909 = select_19 == 6'h38; // @[Switch.scala 41:52:@35068.4]
  assign output_56_19 = io_outValid_19 & _T_73909; // @[Switch.scala 41:38:@35069.4]
  assign _T_73912 = select_20 == 6'h38; // @[Switch.scala 41:52:@35071.4]
  assign output_56_20 = io_outValid_20 & _T_73912; // @[Switch.scala 41:38:@35072.4]
  assign _T_73915 = select_21 == 6'h38; // @[Switch.scala 41:52:@35074.4]
  assign output_56_21 = io_outValid_21 & _T_73915; // @[Switch.scala 41:38:@35075.4]
  assign _T_73918 = select_22 == 6'h38; // @[Switch.scala 41:52:@35077.4]
  assign output_56_22 = io_outValid_22 & _T_73918; // @[Switch.scala 41:38:@35078.4]
  assign _T_73921 = select_23 == 6'h38; // @[Switch.scala 41:52:@35080.4]
  assign output_56_23 = io_outValid_23 & _T_73921; // @[Switch.scala 41:38:@35081.4]
  assign _T_73924 = select_24 == 6'h38; // @[Switch.scala 41:52:@35083.4]
  assign output_56_24 = io_outValid_24 & _T_73924; // @[Switch.scala 41:38:@35084.4]
  assign _T_73927 = select_25 == 6'h38; // @[Switch.scala 41:52:@35086.4]
  assign output_56_25 = io_outValid_25 & _T_73927; // @[Switch.scala 41:38:@35087.4]
  assign _T_73930 = select_26 == 6'h38; // @[Switch.scala 41:52:@35089.4]
  assign output_56_26 = io_outValid_26 & _T_73930; // @[Switch.scala 41:38:@35090.4]
  assign _T_73933 = select_27 == 6'h38; // @[Switch.scala 41:52:@35092.4]
  assign output_56_27 = io_outValid_27 & _T_73933; // @[Switch.scala 41:38:@35093.4]
  assign _T_73936 = select_28 == 6'h38; // @[Switch.scala 41:52:@35095.4]
  assign output_56_28 = io_outValid_28 & _T_73936; // @[Switch.scala 41:38:@35096.4]
  assign _T_73939 = select_29 == 6'h38; // @[Switch.scala 41:52:@35098.4]
  assign output_56_29 = io_outValid_29 & _T_73939; // @[Switch.scala 41:38:@35099.4]
  assign _T_73942 = select_30 == 6'h38; // @[Switch.scala 41:52:@35101.4]
  assign output_56_30 = io_outValid_30 & _T_73942; // @[Switch.scala 41:38:@35102.4]
  assign _T_73945 = select_31 == 6'h38; // @[Switch.scala 41:52:@35104.4]
  assign output_56_31 = io_outValid_31 & _T_73945; // @[Switch.scala 41:38:@35105.4]
  assign _T_73948 = select_32 == 6'h38; // @[Switch.scala 41:52:@35107.4]
  assign output_56_32 = io_outValid_32 & _T_73948; // @[Switch.scala 41:38:@35108.4]
  assign _T_73951 = select_33 == 6'h38; // @[Switch.scala 41:52:@35110.4]
  assign output_56_33 = io_outValid_33 & _T_73951; // @[Switch.scala 41:38:@35111.4]
  assign _T_73954 = select_34 == 6'h38; // @[Switch.scala 41:52:@35113.4]
  assign output_56_34 = io_outValid_34 & _T_73954; // @[Switch.scala 41:38:@35114.4]
  assign _T_73957 = select_35 == 6'h38; // @[Switch.scala 41:52:@35116.4]
  assign output_56_35 = io_outValid_35 & _T_73957; // @[Switch.scala 41:38:@35117.4]
  assign _T_73960 = select_36 == 6'h38; // @[Switch.scala 41:52:@35119.4]
  assign output_56_36 = io_outValid_36 & _T_73960; // @[Switch.scala 41:38:@35120.4]
  assign _T_73963 = select_37 == 6'h38; // @[Switch.scala 41:52:@35122.4]
  assign output_56_37 = io_outValid_37 & _T_73963; // @[Switch.scala 41:38:@35123.4]
  assign _T_73966 = select_38 == 6'h38; // @[Switch.scala 41:52:@35125.4]
  assign output_56_38 = io_outValid_38 & _T_73966; // @[Switch.scala 41:38:@35126.4]
  assign _T_73969 = select_39 == 6'h38; // @[Switch.scala 41:52:@35128.4]
  assign output_56_39 = io_outValid_39 & _T_73969; // @[Switch.scala 41:38:@35129.4]
  assign _T_73972 = select_40 == 6'h38; // @[Switch.scala 41:52:@35131.4]
  assign output_56_40 = io_outValid_40 & _T_73972; // @[Switch.scala 41:38:@35132.4]
  assign _T_73975 = select_41 == 6'h38; // @[Switch.scala 41:52:@35134.4]
  assign output_56_41 = io_outValid_41 & _T_73975; // @[Switch.scala 41:38:@35135.4]
  assign _T_73978 = select_42 == 6'h38; // @[Switch.scala 41:52:@35137.4]
  assign output_56_42 = io_outValid_42 & _T_73978; // @[Switch.scala 41:38:@35138.4]
  assign _T_73981 = select_43 == 6'h38; // @[Switch.scala 41:52:@35140.4]
  assign output_56_43 = io_outValid_43 & _T_73981; // @[Switch.scala 41:38:@35141.4]
  assign _T_73984 = select_44 == 6'h38; // @[Switch.scala 41:52:@35143.4]
  assign output_56_44 = io_outValid_44 & _T_73984; // @[Switch.scala 41:38:@35144.4]
  assign _T_73987 = select_45 == 6'h38; // @[Switch.scala 41:52:@35146.4]
  assign output_56_45 = io_outValid_45 & _T_73987; // @[Switch.scala 41:38:@35147.4]
  assign _T_73990 = select_46 == 6'h38; // @[Switch.scala 41:52:@35149.4]
  assign output_56_46 = io_outValid_46 & _T_73990; // @[Switch.scala 41:38:@35150.4]
  assign _T_73993 = select_47 == 6'h38; // @[Switch.scala 41:52:@35152.4]
  assign output_56_47 = io_outValid_47 & _T_73993; // @[Switch.scala 41:38:@35153.4]
  assign _T_73996 = select_48 == 6'h38; // @[Switch.scala 41:52:@35155.4]
  assign output_56_48 = io_outValid_48 & _T_73996; // @[Switch.scala 41:38:@35156.4]
  assign _T_73999 = select_49 == 6'h38; // @[Switch.scala 41:52:@35158.4]
  assign output_56_49 = io_outValid_49 & _T_73999; // @[Switch.scala 41:38:@35159.4]
  assign _T_74002 = select_50 == 6'h38; // @[Switch.scala 41:52:@35161.4]
  assign output_56_50 = io_outValid_50 & _T_74002; // @[Switch.scala 41:38:@35162.4]
  assign _T_74005 = select_51 == 6'h38; // @[Switch.scala 41:52:@35164.4]
  assign output_56_51 = io_outValid_51 & _T_74005; // @[Switch.scala 41:38:@35165.4]
  assign _T_74008 = select_52 == 6'h38; // @[Switch.scala 41:52:@35167.4]
  assign output_56_52 = io_outValid_52 & _T_74008; // @[Switch.scala 41:38:@35168.4]
  assign _T_74011 = select_53 == 6'h38; // @[Switch.scala 41:52:@35170.4]
  assign output_56_53 = io_outValid_53 & _T_74011; // @[Switch.scala 41:38:@35171.4]
  assign _T_74014 = select_54 == 6'h38; // @[Switch.scala 41:52:@35173.4]
  assign output_56_54 = io_outValid_54 & _T_74014; // @[Switch.scala 41:38:@35174.4]
  assign _T_74017 = select_55 == 6'h38; // @[Switch.scala 41:52:@35176.4]
  assign output_56_55 = io_outValid_55 & _T_74017; // @[Switch.scala 41:38:@35177.4]
  assign _T_74020 = select_56 == 6'h38; // @[Switch.scala 41:52:@35179.4]
  assign output_56_56 = io_outValid_56 & _T_74020; // @[Switch.scala 41:38:@35180.4]
  assign _T_74023 = select_57 == 6'h38; // @[Switch.scala 41:52:@35182.4]
  assign output_56_57 = io_outValid_57 & _T_74023; // @[Switch.scala 41:38:@35183.4]
  assign _T_74026 = select_58 == 6'h38; // @[Switch.scala 41:52:@35185.4]
  assign output_56_58 = io_outValid_58 & _T_74026; // @[Switch.scala 41:38:@35186.4]
  assign _T_74029 = select_59 == 6'h38; // @[Switch.scala 41:52:@35188.4]
  assign output_56_59 = io_outValid_59 & _T_74029; // @[Switch.scala 41:38:@35189.4]
  assign _T_74032 = select_60 == 6'h38; // @[Switch.scala 41:52:@35191.4]
  assign output_56_60 = io_outValid_60 & _T_74032; // @[Switch.scala 41:38:@35192.4]
  assign _T_74035 = select_61 == 6'h38; // @[Switch.scala 41:52:@35194.4]
  assign output_56_61 = io_outValid_61 & _T_74035; // @[Switch.scala 41:38:@35195.4]
  assign _T_74038 = select_62 == 6'h38; // @[Switch.scala 41:52:@35197.4]
  assign output_56_62 = io_outValid_62 & _T_74038; // @[Switch.scala 41:38:@35198.4]
  assign _T_74041 = select_63 == 6'h38; // @[Switch.scala 41:52:@35200.4]
  assign output_56_63 = io_outValid_63 & _T_74041; // @[Switch.scala 41:38:@35201.4]
  assign _T_74049 = {output_56_7,output_56_6,output_56_5,output_56_4,output_56_3,output_56_2,output_56_1,output_56_0}; // @[Switch.scala 43:31:@35209.4]
  assign _T_74057 = {output_56_15,output_56_14,output_56_13,output_56_12,output_56_11,output_56_10,output_56_9,output_56_8,_T_74049}; // @[Switch.scala 43:31:@35217.4]
  assign _T_74064 = {output_56_23,output_56_22,output_56_21,output_56_20,output_56_19,output_56_18,output_56_17,output_56_16}; // @[Switch.scala 43:31:@35224.4]
  assign _T_74073 = {output_56_31,output_56_30,output_56_29,output_56_28,output_56_27,output_56_26,output_56_25,output_56_24,_T_74064,_T_74057}; // @[Switch.scala 43:31:@35233.4]
  assign _T_74080 = {output_56_39,output_56_38,output_56_37,output_56_36,output_56_35,output_56_34,output_56_33,output_56_32}; // @[Switch.scala 43:31:@35240.4]
  assign _T_74088 = {output_56_47,output_56_46,output_56_45,output_56_44,output_56_43,output_56_42,output_56_41,output_56_40,_T_74080}; // @[Switch.scala 43:31:@35248.4]
  assign _T_74095 = {output_56_55,output_56_54,output_56_53,output_56_52,output_56_51,output_56_50,output_56_49,output_56_48}; // @[Switch.scala 43:31:@35255.4]
  assign _T_74104 = {output_56_63,output_56_62,output_56_61,output_56_60,output_56_59,output_56_58,output_56_57,output_56_56,_T_74095,_T_74088}; // @[Switch.scala 43:31:@35264.4]
  assign _T_74105 = {_T_74104,_T_74073}; // @[Switch.scala 43:31:@35265.4]
  assign _T_74109 = select_0 == 6'h39; // @[Switch.scala 41:52:@35268.4]
  assign output_57_0 = io_outValid_0 & _T_74109; // @[Switch.scala 41:38:@35269.4]
  assign _T_74112 = select_1 == 6'h39; // @[Switch.scala 41:52:@35271.4]
  assign output_57_1 = io_outValid_1 & _T_74112; // @[Switch.scala 41:38:@35272.4]
  assign _T_74115 = select_2 == 6'h39; // @[Switch.scala 41:52:@35274.4]
  assign output_57_2 = io_outValid_2 & _T_74115; // @[Switch.scala 41:38:@35275.4]
  assign _T_74118 = select_3 == 6'h39; // @[Switch.scala 41:52:@35277.4]
  assign output_57_3 = io_outValid_3 & _T_74118; // @[Switch.scala 41:38:@35278.4]
  assign _T_74121 = select_4 == 6'h39; // @[Switch.scala 41:52:@35280.4]
  assign output_57_4 = io_outValid_4 & _T_74121; // @[Switch.scala 41:38:@35281.4]
  assign _T_74124 = select_5 == 6'h39; // @[Switch.scala 41:52:@35283.4]
  assign output_57_5 = io_outValid_5 & _T_74124; // @[Switch.scala 41:38:@35284.4]
  assign _T_74127 = select_6 == 6'h39; // @[Switch.scala 41:52:@35286.4]
  assign output_57_6 = io_outValid_6 & _T_74127; // @[Switch.scala 41:38:@35287.4]
  assign _T_74130 = select_7 == 6'h39; // @[Switch.scala 41:52:@35289.4]
  assign output_57_7 = io_outValid_7 & _T_74130; // @[Switch.scala 41:38:@35290.4]
  assign _T_74133 = select_8 == 6'h39; // @[Switch.scala 41:52:@35292.4]
  assign output_57_8 = io_outValid_8 & _T_74133; // @[Switch.scala 41:38:@35293.4]
  assign _T_74136 = select_9 == 6'h39; // @[Switch.scala 41:52:@35295.4]
  assign output_57_9 = io_outValid_9 & _T_74136; // @[Switch.scala 41:38:@35296.4]
  assign _T_74139 = select_10 == 6'h39; // @[Switch.scala 41:52:@35298.4]
  assign output_57_10 = io_outValid_10 & _T_74139; // @[Switch.scala 41:38:@35299.4]
  assign _T_74142 = select_11 == 6'h39; // @[Switch.scala 41:52:@35301.4]
  assign output_57_11 = io_outValid_11 & _T_74142; // @[Switch.scala 41:38:@35302.4]
  assign _T_74145 = select_12 == 6'h39; // @[Switch.scala 41:52:@35304.4]
  assign output_57_12 = io_outValid_12 & _T_74145; // @[Switch.scala 41:38:@35305.4]
  assign _T_74148 = select_13 == 6'h39; // @[Switch.scala 41:52:@35307.4]
  assign output_57_13 = io_outValid_13 & _T_74148; // @[Switch.scala 41:38:@35308.4]
  assign _T_74151 = select_14 == 6'h39; // @[Switch.scala 41:52:@35310.4]
  assign output_57_14 = io_outValid_14 & _T_74151; // @[Switch.scala 41:38:@35311.4]
  assign _T_74154 = select_15 == 6'h39; // @[Switch.scala 41:52:@35313.4]
  assign output_57_15 = io_outValid_15 & _T_74154; // @[Switch.scala 41:38:@35314.4]
  assign _T_74157 = select_16 == 6'h39; // @[Switch.scala 41:52:@35316.4]
  assign output_57_16 = io_outValid_16 & _T_74157; // @[Switch.scala 41:38:@35317.4]
  assign _T_74160 = select_17 == 6'h39; // @[Switch.scala 41:52:@35319.4]
  assign output_57_17 = io_outValid_17 & _T_74160; // @[Switch.scala 41:38:@35320.4]
  assign _T_74163 = select_18 == 6'h39; // @[Switch.scala 41:52:@35322.4]
  assign output_57_18 = io_outValid_18 & _T_74163; // @[Switch.scala 41:38:@35323.4]
  assign _T_74166 = select_19 == 6'h39; // @[Switch.scala 41:52:@35325.4]
  assign output_57_19 = io_outValid_19 & _T_74166; // @[Switch.scala 41:38:@35326.4]
  assign _T_74169 = select_20 == 6'h39; // @[Switch.scala 41:52:@35328.4]
  assign output_57_20 = io_outValid_20 & _T_74169; // @[Switch.scala 41:38:@35329.4]
  assign _T_74172 = select_21 == 6'h39; // @[Switch.scala 41:52:@35331.4]
  assign output_57_21 = io_outValid_21 & _T_74172; // @[Switch.scala 41:38:@35332.4]
  assign _T_74175 = select_22 == 6'h39; // @[Switch.scala 41:52:@35334.4]
  assign output_57_22 = io_outValid_22 & _T_74175; // @[Switch.scala 41:38:@35335.4]
  assign _T_74178 = select_23 == 6'h39; // @[Switch.scala 41:52:@35337.4]
  assign output_57_23 = io_outValid_23 & _T_74178; // @[Switch.scala 41:38:@35338.4]
  assign _T_74181 = select_24 == 6'h39; // @[Switch.scala 41:52:@35340.4]
  assign output_57_24 = io_outValid_24 & _T_74181; // @[Switch.scala 41:38:@35341.4]
  assign _T_74184 = select_25 == 6'h39; // @[Switch.scala 41:52:@35343.4]
  assign output_57_25 = io_outValid_25 & _T_74184; // @[Switch.scala 41:38:@35344.4]
  assign _T_74187 = select_26 == 6'h39; // @[Switch.scala 41:52:@35346.4]
  assign output_57_26 = io_outValid_26 & _T_74187; // @[Switch.scala 41:38:@35347.4]
  assign _T_74190 = select_27 == 6'h39; // @[Switch.scala 41:52:@35349.4]
  assign output_57_27 = io_outValid_27 & _T_74190; // @[Switch.scala 41:38:@35350.4]
  assign _T_74193 = select_28 == 6'h39; // @[Switch.scala 41:52:@35352.4]
  assign output_57_28 = io_outValid_28 & _T_74193; // @[Switch.scala 41:38:@35353.4]
  assign _T_74196 = select_29 == 6'h39; // @[Switch.scala 41:52:@35355.4]
  assign output_57_29 = io_outValid_29 & _T_74196; // @[Switch.scala 41:38:@35356.4]
  assign _T_74199 = select_30 == 6'h39; // @[Switch.scala 41:52:@35358.4]
  assign output_57_30 = io_outValid_30 & _T_74199; // @[Switch.scala 41:38:@35359.4]
  assign _T_74202 = select_31 == 6'h39; // @[Switch.scala 41:52:@35361.4]
  assign output_57_31 = io_outValid_31 & _T_74202; // @[Switch.scala 41:38:@35362.4]
  assign _T_74205 = select_32 == 6'h39; // @[Switch.scala 41:52:@35364.4]
  assign output_57_32 = io_outValid_32 & _T_74205; // @[Switch.scala 41:38:@35365.4]
  assign _T_74208 = select_33 == 6'h39; // @[Switch.scala 41:52:@35367.4]
  assign output_57_33 = io_outValid_33 & _T_74208; // @[Switch.scala 41:38:@35368.4]
  assign _T_74211 = select_34 == 6'h39; // @[Switch.scala 41:52:@35370.4]
  assign output_57_34 = io_outValid_34 & _T_74211; // @[Switch.scala 41:38:@35371.4]
  assign _T_74214 = select_35 == 6'h39; // @[Switch.scala 41:52:@35373.4]
  assign output_57_35 = io_outValid_35 & _T_74214; // @[Switch.scala 41:38:@35374.4]
  assign _T_74217 = select_36 == 6'h39; // @[Switch.scala 41:52:@35376.4]
  assign output_57_36 = io_outValid_36 & _T_74217; // @[Switch.scala 41:38:@35377.4]
  assign _T_74220 = select_37 == 6'h39; // @[Switch.scala 41:52:@35379.4]
  assign output_57_37 = io_outValid_37 & _T_74220; // @[Switch.scala 41:38:@35380.4]
  assign _T_74223 = select_38 == 6'h39; // @[Switch.scala 41:52:@35382.4]
  assign output_57_38 = io_outValid_38 & _T_74223; // @[Switch.scala 41:38:@35383.4]
  assign _T_74226 = select_39 == 6'h39; // @[Switch.scala 41:52:@35385.4]
  assign output_57_39 = io_outValid_39 & _T_74226; // @[Switch.scala 41:38:@35386.4]
  assign _T_74229 = select_40 == 6'h39; // @[Switch.scala 41:52:@35388.4]
  assign output_57_40 = io_outValid_40 & _T_74229; // @[Switch.scala 41:38:@35389.4]
  assign _T_74232 = select_41 == 6'h39; // @[Switch.scala 41:52:@35391.4]
  assign output_57_41 = io_outValid_41 & _T_74232; // @[Switch.scala 41:38:@35392.4]
  assign _T_74235 = select_42 == 6'h39; // @[Switch.scala 41:52:@35394.4]
  assign output_57_42 = io_outValid_42 & _T_74235; // @[Switch.scala 41:38:@35395.4]
  assign _T_74238 = select_43 == 6'h39; // @[Switch.scala 41:52:@35397.4]
  assign output_57_43 = io_outValid_43 & _T_74238; // @[Switch.scala 41:38:@35398.4]
  assign _T_74241 = select_44 == 6'h39; // @[Switch.scala 41:52:@35400.4]
  assign output_57_44 = io_outValid_44 & _T_74241; // @[Switch.scala 41:38:@35401.4]
  assign _T_74244 = select_45 == 6'h39; // @[Switch.scala 41:52:@35403.4]
  assign output_57_45 = io_outValid_45 & _T_74244; // @[Switch.scala 41:38:@35404.4]
  assign _T_74247 = select_46 == 6'h39; // @[Switch.scala 41:52:@35406.4]
  assign output_57_46 = io_outValid_46 & _T_74247; // @[Switch.scala 41:38:@35407.4]
  assign _T_74250 = select_47 == 6'h39; // @[Switch.scala 41:52:@35409.4]
  assign output_57_47 = io_outValid_47 & _T_74250; // @[Switch.scala 41:38:@35410.4]
  assign _T_74253 = select_48 == 6'h39; // @[Switch.scala 41:52:@35412.4]
  assign output_57_48 = io_outValid_48 & _T_74253; // @[Switch.scala 41:38:@35413.4]
  assign _T_74256 = select_49 == 6'h39; // @[Switch.scala 41:52:@35415.4]
  assign output_57_49 = io_outValid_49 & _T_74256; // @[Switch.scala 41:38:@35416.4]
  assign _T_74259 = select_50 == 6'h39; // @[Switch.scala 41:52:@35418.4]
  assign output_57_50 = io_outValid_50 & _T_74259; // @[Switch.scala 41:38:@35419.4]
  assign _T_74262 = select_51 == 6'h39; // @[Switch.scala 41:52:@35421.4]
  assign output_57_51 = io_outValid_51 & _T_74262; // @[Switch.scala 41:38:@35422.4]
  assign _T_74265 = select_52 == 6'h39; // @[Switch.scala 41:52:@35424.4]
  assign output_57_52 = io_outValid_52 & _T_74265; // @[Switch.scala 41:38:@35425.4]
  assign _T_74268 = select_53 == 6'h39; // @[Switch.scala 41:52:@35427.4]
  assign output_57_53 = io_outValid_53 & _T_74268; // @[Switch.scala 41:38:@35428.4]
  assign _T_74271 = select_54 == 6'h39; // @[Switch.scala 41:52:@35430.4]
  assign output_57_54 = io_outValid_54 & _T_74271; // @[Switch.scala 41:38:@35431.4]
  assign _T_74274 = select_55 == 6'h39; // @[Switch.scala 41:52:@35433.4]
  assign output_57_55 = io_outValid_55 & _T_74274; // @[Switch.scala 41:38:@35434.4]
  assign _T_74277 = select_56 == 6'h39; // @[Switch.scala 41:52:@35436.4]
  assign output_57_56 = io_outValid_56 & _T_74277; // @[Switch.scala 41:38:@35437.4]
  assign _T_74280 = select_57 == 6'h39; // @[Switch.scala 41:52:@35439.4]
  assign output_57_57 = io_outValid_57 & _T_74280; // @[Switch.scala 41:38:@35440.4]
  assign _T_74283 = select_58 == 6'h39; // @[Switch.scala 41:52:@35442.4]
  assign output_57_58 = io_outValid_58 & _T_74283; // @[Switch.scala 41:38:@35443.4]
  assign _T_74286 = select_59 == 6'h39; // @[Switch.scala 41:52:@35445.4]
  assign output_57_59 = io_outValid_59 & _T_74286; // @[Switch.scala 41:38:@35446.4]
  assign _T_74289 = select_60 == 6'h39; // @[Switch.scala 41:52:@35448.4]
  assign output_57_60 = io_outValid_60 & _T_74289; // @[Switch.scala 41:38:@35449.4]
  assign _T_74292 = select_61 == 6'h39; // @[Switch.scala 41:52:@35451.4]
  assign output_57_61 = io_outValid_61 & _T_74292; // @[Switch.scala 41:38:@35452.4]
  assign _T_74295 = select_62 == 6'h39; // @[Switch.scala 41:52:@35454.4]
  assign output_57_62 = io_outValid_62 & _T_74295; // @[Switch.scala 41:38:@35455.4]
  assign _T_74298 = select_63 == 6'h39; // @[Switch.scala 41:52:@35457.4]
  assign output_57_63 = io_outValid_63 & _T_74298; // @[Switch.scala 41:38:@35458.4]
  assign _T_74306 = {output_57_7,output_57_6,output_57_5,output_57_4,output_57_3,output_57_2,output_57_1,output_57_0}; // @[Switch.scala 43:31:@35466.4]
  assign _T_74314 = {output_57_15,output_57_14,output_57_13,output_57_12,output_57_11,output_57_10,output_57_9,output_57_8,_T_74306}; // @[Switch.scala 43:31:@35474.4]
  assign _T_74321 = {output_57_23,output_57_22,output_57_21,output_57_20,output_57_19,output_57_18,output_57_17,output_57_16}; // @[Switch.scala 43:31:@35481.4]
  assign _T_74330 = {output_57_31,output_57_30,output_57_29,output_57_28,output_57_27,output_57_26,output_57_25,output_57_24,_T_74321,_T_74314}; // @[Switch.scala 43:31:@35490.4]
  assign _T_74337 = {output_57_39,output_57_38,output_57_37,output_57_36,output_57_35,output_57_34,output_57_33,output_57_32}; // @[Switch.scala 43:31:@35497.4]
  assign _T_74345 = {output_57_47,output_57_46,output_57_45,output_57_44,output_57_43,output_57_42,output_57_41,output_57_40,_T_74337}; // @[Switch.scala 43:31:@35505.4]
  assign _T_74352 = {output_57_55,output_57_54,output_57_53,output_57_52,output_57_51,output_57_50,output_57_49,output_57_48}; // @[Switch.scala 43:31:@35512.4]
  assign _T_74361 = {output_57_63,output_57_62,output_57_61,output_57_60,output_57_59,output_57_58,output_57_57,output_57_56,_T_74352,_T_74345}; // @[Switch.scala 43:31:@35521.4]
  assign _T_74362 = {_T_74361,_T_74330}; // @[Switch.scala 43:31:@35522.4]
  assign _T_74366 = select_0 == 6'h3a; // @[Switch.scala 41:52:@35525.4]
  assign output_58_0 = io_outValid_0 & _T_74366; // @[Switch.scala 41:38:@35526.4]
  assign _T_74369 = select_1 == 6'h3a; // @[Switch.scala 41:52:@35528.4]
  assign output_58_1 = io_outValid_1 & _T_74369; // @[Switch.scala 41:38:@35529.4]
  assign _T_74372 = select_2 == 6'h3a; // @[Switch.scala 41:52:@35531.4]
  assign output_58_2 = io_outValid_2 & _T_74372; // @[Switch.scala 41:38:@35532.4]
  assign _T_74375 = select_3 == 6'h3a; // @[Switch.scala 41:52:@35534.4]
  assign output_58_3 = io_outValid_3 & _T_74375; // @[Switch.scala 41:38:@35535.4]
  assign _T_74378 = select_4 == 6'h3a; // @[Switch.scala 41:52:@35537.4]
  assign output_58_4 = io_outValid_4 & _T_74378; // @[Switch.scala 41:38:@35538.4]
  assign _T_74381 = select_5 == 6'h3a; // @[Switch.scala 41:52:@35540.4]
  assign output_58_5 = io_outValid_5 & _T_74381; // @[Switch.scala 41:38:@35541.4]
  assign _T_74384 = select_6 == 6'h3a; // @[Switch.scala 41:52:@35543.4]
  assign output_58_6 = io_outValid_6 & _T_74384; // @[Switch.scala 41:38:@35544.4]
  assign _T_74387 = select_7 == 6'h3a; // @[Switch.scala 41:52:@35546.4]
  assign output_58_7 = io_outValid_7 & _T_74387; // @[Switch.scala 41:38:@35547.4]
  assign _T_74390 = select_8 == 6'h3a; // @[Switch.scala 41:52:@35549.4]
  assign output_58_8 = io_outValid_8 & _T_74390; // @[Switch.scala 41:38:@35550.4]
  assign _T_74393 = select_9 == 6'h3a; // @[Switch.scala 41:52:@35552.4]
  assign output_58_9 = io_outValid_9 & _T_74393; // @[Switch.scala 41:38:@35553.4]
  assign _T_74396 = select_10 == 6'h3a; // @[Switch.scala 41:52:@35555.4]
  assign output_58_10 = io_outValid_10 & _T_74396; // @[Switch.scala 41:38:@35556.4]
  assign _T_74399 = select_11 == 6'h3a; // @[Switch.scala 41:52:@35558.4]
  assign output_58_11 = io_outValid_11 & _T_74399; // @[Switch.scala 41:38:@35559.4]
  assign _T_74402 = select_12 == 6'h3a; // @[Switch.scala 41:52:@35561.4]
  assign output_58_12 = io_outValid_12 & _T_74402; // @[Switch.scala 41:38:@35562.4]
  assign _T_74405 = select_13 == 6'h3a; // @[Switch.scala 41:52:@35564.4]
  assign output_58_13 = io_outValid_13 & _T_74405; // @[Switch.scala 41:38:@35565.4]
  assign _T_74408 = select_14 == 6'h3a; // @[Switch.scala 41:52:@35567.4]
  assign output_58_14 = io_outValid_14 & _T_74408; // @[Switch.scala 41:38:@35568.4]
  assign _T_74411 = select_15 == 6'h3a; // @[Switch.scala 41:52:@35570.4]
  assign output_58_15 = io_outValid_15 & _T_74411; // @[Switch.scala 41:38:@35571.4]
  assign _T_74414 = select_16 == 6'h3a; // @[Switch.scala 41:52:@35573.4]
  assign output_58_16 = io_outValid_16 & _T_74414; // @[Switch.scala 41:38:@35574.4]
  assign _T_74417 = select_17 == 6'h3a; // @[Switch.scala 41:52:@35576.4]
  assign output_58_17 = io_outValid_17 & _T_74417; // @[Switch.scala 41:38:@35577.4]
  assign _T_74420 = select_18 == 6'h3a; // @[Switch.scala 41:52:@35579.4]
  assign output_58_18 = io_outValid_18 & _T_74420; // @[Switch.scala 41:38:@35580.4]
  assign _T_74423 = select_19 == 6'h3a; // @[Switch.scala 41:52:@35582.4]
  assign output_58_19 = io_outValid_19 & _T_74423; // @[Switch.scala 41:38:@35583.4]
  assign _T_74426 = select_20 == 6'h3a; // @[Switch.scala 41:52:@35585.4]
  assign output_58_20 = io_outValid_20 & _T_74426; // @[Switch.scala 41:38:@35586.4]
  assign _T_74429 = select_21 == 6'h3a; // @[Switch.scala 41:52:@35588.4]
  assign output_58_21 = io_outValid_21 & _T_74429; // @[Switch.scala 41:38:@35589.4]
  assign _T_74432 = select_22 == 6'h3a; // @[Switch.scala 41:52:@35591.4]
  assign output_58_22 = io_outValid_22 & _T_74432; // @[Switch.scala 41:38:@35592.4]
  assign _T_74435 = select_23 == 6'h3a; // @[Switch.scala 41:52:@35594.4]
  assign output_58_23 = io_outValid_23 & _T_74435; // @[Switch.scala 41:38:@35595.4]
  assign _T_74438 = select_24 == 6'h3a; // @[Switch.scala 41:52:@35597.4]
  assign output_58_24 = io_outValid_24 & _T_74438; // @[Switch.scala 41:38:@35598.4]
  assign _T_74441 = select_25 == 6'h3a; // @[Switch.scala 41:52:@35600.4]
  assign output_58_25 = io_outValid_25 & _T_74441; // @[Switch.scala 41:38:@35601.4]
  assign _T_74444 = select_26 == 6'h3a; // @[Switch.scala 41:52:@35603.4]
  assign output_58_26 = io_outValid_26 & _T_74444; // @[Switch.scala 41:38:@35604.4]
  assign _T_74447 = select_27 == 6'h3a; // @[Switch.scala 41:52:@35606.4]
  assign output_58_27 = io_outValid_27 & _T_74447; // @[Switch.scala 41:38:@35607.4]
  assign _T_74450 = select_28 == 6'h3a; // @[Switch.scala 41:52:@35609.4]
  assign output_58_28 = io_outValid_28 & _T_74450; // @[Switch.scala 41:38:@35610.4]
  assign _T_74453 = select_29 == 6'h3a; // @[Switch.scala 41:52:@35612.4]
  assign output_58_29 = io_outValid_29 & _T_74453; // @[Switch.scala 41:38:@35613.4]
  assign _T_74456 = select_30 == 6'h3a; // @[Switch.scala 41:52:@35615.4]
  assign output_58_30 = io_outValid_30 & _T_74456; // @[Switch.scala 41:38:@35616.4]
  assign _T_74459 = select_31 == 6'h3a; // @[Switch.scala 41:52:@35618.4]
  assign output_58_31 = io_outValid_31 & _T_74459; // @[Switch.scala 41:38:@35619.4]
  assign _T_74462 = select_32 == 6'h3a; // @[Switch.scala 41:52:@35621.4]
  assign output_58_32 = io_outValid_32 & _T_74462; // @[Switch.scala 41:38:@35622.4]
  assign _T_74465 = select_33 == 6'h3a; // @[Switch.scala 41:52:@35624.4]
  assign output_58_33 = io_outValid_33 & _T_74465; // @[Switch.scala 41:38:@35625.4]
  assign _T_74468 = select_34 == 6'h3a; // @[Switch.scala 41:52:@35627.4]
  assign output_58_34 = io_outValid_34 & _T_74468; // @[Switch.scala 41:38:@35628.4]
  assign _T_74471 = select_35 == 6'h3a; // @[Switch.scala 41:52:@35630.4]
  assign output_58_35 = io_outValid_35 & _T_74471; // @[Switch.scala 41:38:@35631.4]
  assign _T_74474 = select_36 == 6'h3a; // @[Switch.scala 41:52:@35633.4]
  assign output_58_36 = io_outValid_36 & _T_74474; // @[Switch.scala 41:38:@35634.4]
  assign _T_74477 = select_37 == 6'h3a; // @[Switch.scala 41:52:@35636.4]
  assign output_58_37 = io_outValid_37 & _T_74477; // @[Switch.scala 41:38:@35637.4]
  assign _T_74480 = select_38 == 6'h3a; // @[Switch.scala 41:52:@35639.4]
  assign output_58_38 = io_outValid_38 & _T_74480; // @[Switch.scala 41:38:@35640.4]
  assign _T_74483 = select_39 == 6'h3a; // @[Switch.scala 41:52:@35642.4]
  assign output_58_39 = io_outValid_39 & _T_74483; // @[Switch.scala 41:38:@35643.4]
  assign _T_74486 = select_40 == 6'h3a; // @[Switch.scala 41:52:@35645.4]
  assign output_58_40 = io_outValid_40 & _T_74486; // @[Switch.scala 41:38:@35646.4]
  assign _T_74489 = select_41 == 6'h3a; // @[Switch.scala 41:52:@35648.4]
  assign output_58_41 = io_outValid_41 & _T_74489; // @[Switch.scala 41:38:@35649.4]
  assign _T_74492 = select_42 == 6'h3a; // @[Switch.scala 41:52:@35651.4]
  assign output_58_42 = io_outValid_42 & _T_74492; // @[Switch.scala 41:38:@35652.4]
  assign _T_74495 = select_43 == 6'h3a; // @[Switch.scala 41:52:@35654.4]
  assign output_58_43 = io_outValid_43 & _T_74495; // @[Switch.scala 41:38:@35655.4]
  assign _T_74498 = select_44 == 6'h3a; // @[Switch.scala 41:52:@35657.4]
  assign output_58_44 = io_outValid_44 & _T_74498; // @[Switch.scala 41:38:@35658.4]
  assign _T_74501 = select_45 == 6'h3a; // @[Switch.scala 41:52:@35660.4]
  assign output_58_45 = io_outValid_45 & _T_74501; // @[Switch.scala 41:38:@35661.4]
  assign _T_74504 = select_46 == 6'h3a; // @[Switch.scala 41:52:@35663.4]
  assign output_58_46 = io_outValid_46 & _T_74504; // @[Switch.scala 41:38:@35664.4]
  assign _T_74507 = select_47 == 6'h3a; // @[Switch.scala 41:52:@35666.4]
  assign output_58_47 = io_outValid_47 & _T_74507; // @[Switch.scala 41:38:@35667.4]
  assign _T_74510 = select_48 == 6'h3a; // @[Switch.scala 41:52:@35669.4]
  assign output_58_48 = io_outValid_48 & _T_74510; // @[Switch.scala 41:38:@35670.4]
  assign _T_74513 = select_49 == 6'h3a; // @[Switch.scala 41:52:@35672.4]
  assign output_58_49 = io_outValid_49 & _T_74513; // @[Switch.scala 41:38:@35673.4]
  assign _T_74516 = select_50 == 6'h3a; // @[Switch.scala 41:52:@35675.4]
  assign output_58_50 = io_outValid_50 & _T_74516; // @[Switch.scala 41:38:@35676.4]
  assign _T_74519 = select_51 == 6'h3a; // @[Switch.scala 41:52:@35678.4]
  assign output_58_51 = io_outValid_51 & _T_74519; // @[Switch.scala 41:38:@35679.4]
  assign _T_74522 = select_52 == 6'h3a; // @[Switch.scala 41:52:@35681.4]
  assign output_58_52 = io_outValid_52 & _T_74522; // @[Switch.scala 41:38:@35682.4]
  assign _T_74525 = select_53 == 6'h3a; // @[Switch.scala 41:52:@35684.4]
  assign output_58_53 = io_outValid_53 & _T_74525; // @[Switch.scala 41:38:@35685.4]
  assign _T_74528 = select_54 == 6'h3a; // @[Switch.scala 41:52:@35687.4]
  assign output_58_54 = io_outValid_54 & _T_74528; // @[Switch.scala 41:38:@35688.4]
  assign _T_74531 = select_55 == 6'h3a; // @[Switch.scala 41:52:@35690.4]
  assign output_58_55 = io_outValid_55 & _T_74531; // @[Switch.scala 41:38:@35691.4]
  assign _T_74534 = select_56 == 6'h3a; // @[Switch.scala 41:52:@35693.4]
  assign output_58_56 = io_outValid_56 & _T_74534; // @[Switch.scala 41:38:@35694.4]
  assign _T_74537 = select_57 == 6'h3a; // @[Switch.scala 41:52:@35696.4]
  assign output_58_57 = io_outValid_57 & _T_74537; // @[Switch.scala 41:38:@35697.4]
  assign _T_74540 = select_58 == 6'h3a; // @[Switch.scala 41:52:@35699.4]
  assign output_58_58 = io_outValid_58 & _T_74540; // @[Switch.scala 41:38:@35700.4]
  assign _T_74543 = select_59 == 6'h3a; // @[Switch.scala 41:52:@35702.4]
  assign output_58_59 = io_outValid_59 & _T_74543; // @[Switch.scala 41:38:@35703.4]
  assign _T_74546 = select_60 == 6'h3a; // @[Switch.scala 41:52:@35705.4]
  assign output_58_60 = io_outValid_60 & _T_74546; // @[Switch.scala 41:38:@35706.4]
  assign _T_74549 = select_61 == 6'h3a; // @[Switch.scala 41:52:@35708.4]
  assign output_58_61 = io_outValid_61 & _T_74549; // @[Switch.scala 41:38:@35709.4]
  assign _T_74552 = select_62 == 6'h3a; // @[Switch.scala 41:52:@35711.4]
  assign output_58_62 = io_outValid_62 & _T_74552; // @[Switch.scala 41:38:@35712.4]
  assign _T_74555 = select_63 == 6'h3a; // @[Switch.scala 41:52:@35714.4]
  assign output_58_63 = io_outValid_63 & _T_74555; // @[Switch.scala 41:38:@35715.4]
  assign _T_74563 = {output_58_7,output_58_6,output_58_5,output_58_4,output_58_3,output_58_2,output_58_1,output_58_0}; // @[Switch.scala 43:31:@35723.4]
  assign _T_74571 = {output_58_15,output_58_14,output_58_13,output_58_12,output_58_11,output_58_10,output_58_9,output_58_8,_T_74563}; // @[Switch.scala 43:31:@35731.4]
  assign _T_74578 = {output_58_23,output_58_22,output_58_21,output_58_20,output_58_19,output_58_18,output_58_17,output_58_16}; // @[Switch.scala 43:31:@35738.4]
  assign _T_74587 = {output_58_31,output_58_30,output_58_29,output_58_28,output_58_27,output_58_26,output_58_25,output_58_24,_T_74578,_T_74571}; // @[Switch.scala 43:31:@35747.4]
  assign _T_74594 = {output_58_39,output_58_38,output_58_37,output_58_36,output_58_35,output_58_34,output_58_33,output_58_32}; // @[Switch.scala 43:31:@35754.4]
  assign _T_74602 = {output_58_47,output_58_46,output_58_45,output_58_44,output_58_43,output_58_42,output_58_41,output_58_40,_T_74594}; // @[Switch.scala 43:31:@35762.4]
  assign _T_74609 = {output_58_55,output_58_54,output_58_53,output_58_52,output_58_51,output_58_50,output_58_49,output_58_48}; // @[Switch.scala 43:31:@35769.4]
  assign _T_74618 = {output_58_63,output_58_62,output_58_61,output_58_60,output_58_59,output_58_58,output_58_57,output_58_56,_T_74609,_T_74602}; // @[Switch.scala 43:31:@35778.4]
  assign _T_74619 = {_T_74618,_T_74587}; // @[Switch.scala 43:31:@35779.4]
  assign _T_74623 = select_0 == 6'h3b; // @[Switch.scala 41:52:@35782.4]
  assign output_59_0 = io_outValid_0 & _T_74623; // @[Switch.scala 41:38:@35783.4]
  assign _T_74626 = select_1 == 6'h3b; // @[Switch.scala 41:52:@35785.4]
  assign output_59_1 = io_outValid_1 & _T_74626; // @[Switch.scala 41:38:@35786.4]
  assign _T_74629 = select_2 == 6'h3b; // @[Switch.scala 41:52:@35788.4]
  assign output_59_2 = io_outValid_2 & _T_74629; // @[Switch.scala 41:38:@35789.4]
  assign _T_74632 = select_3 == 6'h3b; // @[Switch.scala 41:52:@35791.4]
  assign output_59_3 = io_outValid_3 & _T_74632; // @[Switch.scala 41:38:@35792.4]
  assign _T_74635 = select_4 == 6'h3b; // @[Switch.scala 41:52:@35794.4]
  assign output_59_4 = io_outValid_4 & _T_74635; // @[Switch.scala 41:38:@35795.4]
  assign _T_74638 = select_5 == 6'h3b; // @[Switch.scala 41:52:@35797.4]
  assign output_59_5 = io_outValid_5 & _T_74638; // @[Switch.scala 41:38:@35798.4]
  assign _T_74641 = select_6 == 6'h3b; // @[Switch.scala 41:52:@35800.4]
  assign output_59_6 = io_outValid_6 & _T_74641; // @[Switch.scala 41:38:@35801.4]
  assign _T_74644 = select_7 == 6'h3b; // @[Switch.scala 41:52:@35803.4]
  assign output_59_7 = io_outValid_7 & _T_74644; // @[Switch.scala 41:38:@35804.4]
  assign _T_74647 = select_8 == 6'h3b; // @[Switch.scala 41:52:@35806.4]
  assign output_59_8 = io_outValid_8 & _T_74647; // @[Switch.scala 41:38:@35807.4]
  assign _T_74650 = select_9 == 6'h3b; // @[Switch.scala 41:52:@35809.4]
  assign output_59_9 = io_outValid_9 & _T_74650; // @[Switch.scala 41:38:@35810.4]
  assign _T_74653 = select_10 == 6'h3b; // @[Switch.scala 41:52:@35812.4]
  assign output_59_10 = io_outValid_10 & _T_74653; // @[Switch.scala 41:38:@35813.4]
  assign _T_74656 = select_11 == 6'h3b; // @[Switch.scala 41:52:@35815.4]
  assign output_59_11 = io_outValid_11 & _T_74656; // @[Switch.scala 41:38:@35816.4]
  assign _T_74659 = select_12 == 6'h3b; // @[Switch.scala 41:52:@35818.4]
  assign output_59_12 = io_outValid_12 & _T_74659; // @[Switch.scala 41:38:@35819.4]
  assign _T_74662 = select_13 == 6'h3b; // @[Switch.scala 41:52:@35821.4]
  assign output_59_13 = io_outValid_13 & _T_74662; // @[Switch.scala 41:38:@35822.4]
  assign _T_74665 = select_14 == 6'h3b; // @[Switch.scala 41:52:@35824.4]
  assign output_59_14 = io_outValid_14 & _T_74665; // @[Switch.scala 41:38:@35825.4]
  assign _T_74668 = select_15 == 6'h3b; // @[Switch.scala 41:52:@35827.4]
  assign output_59_15 = io_outValid_15 & _T_74668; // @[Switch.scala 41:38:@35828.4]
  assign _T_74671 = select_16 == 6'h3b; // @[Switch.scala 41:52:@35830.4]
  assign output_59_16 = io_outValid_16 & _T_74671; // @[Switch.scala 41:38:@35831.4]
  assign _T_74674 = select_17 == 6'h3b; // @[Switch.scala 41:52:@35833.4]
  assign output_59_17 = io_outValid_17 & _T_74674; // @[Switch.scala 41:38:@35834.4]
  assign _T_74677 = select_18 == 6'h3b; // @[Switch.scala 41:52:@35836.4]
  assign output_59_18 = io_outValid_18 & _T_74677; // @[Switch.scala 41:38:@35837.4]
  assign _T_74680 = select_19 == 6'h3b; // @[Switch.scala 41:52:@35839.4]
  assign output_59_19 = io_outValid_19 & _T_74680; // @[Switch.scala 41:38:@35840.4]
  assign _T_74683 = select_20 == 6'h3b; // @[Switch.scala 41:52:@35842.4]
  assign output_59_20 = io_outValid_20 & _T_74683; // @[Switch.scala 41:38:@35843.4]
  assign _T_74686 = select_21 == 6'h3b; // @[Switch.scala 41:52:@35845.4]
  assign output_59_21 = io_outValid_21 & _T_74686; // @[Switch.scala 41:38:@35846.4]
  assign _T_74689 = select_22 == 6'h3b; // @[Switch.scala 41:52:@35848.4]
  assign output_59_22 = io_outValid_22 & _T_74689; // @[Switch.scala 41:38:@35849.4]
  assign _T_74692 = select_23 == 6'h3b; // @[Switch.scala 41:52:@35851.4]
  assign output_59_23 = io_outValid_23 & _T_74692; // @[Switch.scala 41:38:@35852.4]
  assign _T_74695 = select_24 == 6'h3b; // @[Switch.scala 41:52:@35854.4]
  assign output_59_24 = io_outValid_24 & _T_74695; // @[Switch.scala 41:38:@35855.4]
  assign _T_74698 = select_25 == 6'h3b; // @[Switch.scala 41:52:@35857.4]
  assign output_59_25 = io_outValid_25 & _T_74698; // @[Switch.scala 41:38:@35858.4]
  assign _T_74701 = select_26 == 6'h3b; // @[Switch.scala 41:52:@35860.4]
  assign output_59_26 = io_outValid_26 & _T_74701; // @[Switch.scala 41:38:@35861.4]
  assign _T_74704 = select_27 == 6'h3b; // @[Switch.scala 41:52:@35863.4]
  assign output_59_27 = io_outValid_27 & _T_74704; // @[Switch.scala 41:38:@35864.4]
  assign _T_74707 = select_28 == 6'h3b; // @[Switch.scala 41:52:@35866.4]
  assign output_59_28 = io_outValid_28 & _T_74707; // @[Switch.scala 41:38:@35867.4]
  assign _T_74710 = select_29 == 6'h3b; // @[Switch.scala 41:52:@35869.4]
  assign output_59_29 = io_outValid_29 & _T_74710; // @[Switch.scala 41:38:@35870.4]
  assign _T_74713 = select_30 == 6'h3b; // @[Switch.scala 41:52:@35872.4]
  assign output_59_30 = io_outValid_30 & _T_74713; // @[Switch.scala 41:38:@35873.4]
  assign _T_74716 = select_31 == 6'h3b; // @[Switch.scala 41:52:@35875.4]
  assign output_59_31 = io_outValid_31 & _T_74716; // @[Switch.scala 41:38:@35876.4]
  assign _T_74719 = select_32 == 6'h3b; // @[Switch.scala 41:52:@35878.4]
  assign output_59_32 = io_outValid_32 & _T_74719; // @[Switch.scala 41:38:@35879.4]
  assign _T_74722 = select_33 == 6'h3b; // @[Switch.scala 41:52:@35881.4]
  assign output_59_33 = io_outValid_33 & _T_74722; // @[Switch.scala 41:38:@35882.4]
  assign _T_74725 = select_34 == 6'h3b; // @[Switch.scala 41:52:@35884.4]
  assign output_59_34 = io_outValid_34 & _T_74725; // @[Switch.scala 41:38:@35885.4]
  assign _T_74728 = select_35 == 6'h3b; // @[Switch.scala 41:52:@35887.4]
  assign output_59_35 = io_outValid_35 & _T_74728; // @[Switch.scala 41:38:@35888.4]
  assign _T_74731 = select_36 == 6'h3b; // @[Switch.scala 41:52:@35890.4]
  assign output_59_36 = io_outValid_36 & _T_74731; // @[Switch.scala 41:38:@35891.4]
  assign _T_74734 = select_37 == 6'h3b; // @[Switch.scala 41:52:@35893.4]
  assign output_59_37 = io_outValid_37 & _T_74734; // @[Switch.scala 41:38:@35894.4]
  assign _T_74737 = select_38 == 6'h3b; // @[Switch.scala 41:52:@35896.4]
  assign output_59_38 = io_outValid_38 & _T_74737; // @[Switch.scala 41:38:@35897.4]
  assign _T_74740 = select_39 == 6'h3b; // @[Switch.scala 41:52:@35899.4]
  assign output_59_39 = io_outValid_39 & _T_74740; // @[Switch.scala 41:38:@35900.4]
  assign _T_74743 = select_40 == 6'h3b; // @[Switch.scala 41:52:@35902.4]
  assign output_59_40 = io_outValid_40 & _T_74743; // @[Switch.scala 41:38:@35903.4]
  assign _T_74746 = select_41 == 6'h3b; // @[Switch.scala 41:52:@35905.4]
  assign output_59_41 = io_outValid_41 & _T_74746; // @[Switch.scala 41:38:@35906.4]
  assign _T_74749 = select_42 == 6'h3b; // @[Switch.scala 41:52:@35908.4]
  assign output_59_42 = io_outValid_42 & _T_74749; // @[Switch.scala 41:38:@35909.4]
  assign _T_74752 = select_43 == 6'h3b; // @[Switch.scala 41:52:@35911.4]
  assign output_59_43 = io_outValid_43 & _T_74752; // @[Switch.scala 41:38:@35912.4]
  assign _T_74755 = select_44 == 6'h3b; // @[Switch.scala 41:52:@35914.4]
  assign output_59_44 = io_outValid_44 & _T_74755; // @[Switch.scala 41:38:@35915.4]
  assign _T_74758 = select_45 == 6'h3b; // @[Switch.scala 41:52:@35917.4]
  assign output_59_45 = io_outValid_45 & _T_74758; // @[Switch.scala 41:38:@35918.4]
  assign _T_74761 = select_46 == 6'h3b; // @[Switch.scala 41:52:@35920.4]
  assign output_59_46 = io_outValid_46 & _T_74761; // @[Switch.scala 41:38:@35921.4]
  assign _T_74764 = select_47 == 6'h3b; // @[Switch.scala 41:52:@35923.4]
  assign output_59_47 = io_outValid_47 & _T_74764; // @[Switch.scala 41:38:@35924.4]
  assign _T_74767 = select_48 == 6'h3b; // @[Switch.scala 41:52:@35926.4]
  assign output_59_48 = io_outValid_48 & _T_74767; // @[Switch.scala 41:38:@35927.4]
  assign _T_74770 = select_49 == 6'h3b; // @[Switch.scala 41:52:@35929.4]
  assign output_59_49 = io_outValid_49 & _T_74770; // @[Switch.scala 41:38:@35930.4]
  assign _T_74773 = select_50 == 6'h3b; // @[Switch.scala 41:52:@35932.4]
  assign output_59_50 = io_outValid_50 & _T_74773; // @[Switch.scala 41:38:@35933.4]
  assign _T_74776 = select_51 == 6'h3b; // @[Switch.scala 41:52:@35935.4]
  assign output_59_51 = io_outValid_51 & _T_74776; // @[Switch.scala 41:38:@35936.4]
  assign _T_74779 = select_52 == 6'h3b; // @[Switch.scala 41:52:@35938.4]
  assign output_59_52 = io_outValid_52 & _T_74779; // @[Switch.scala 41:38:@35939.4]
  assign _T_74782 = select_53 == 6'h3b; // @[Switch.scala 41:52:@35941.4]
  assign output_59_53 = io_outValid_53 & _T_74782; // @[Switch.scala 41:38:@35942.4]
  assign _T_74785 = select_54 == 6'h3b; // @[Switch.scala 41:52:@35944.4]
  assign output_59_54 = io_outValid_54 & _T_74785; // @[Switch.scala 41:38:@35945.4]
  assign _T_74788 = select_55 == 6'h3b; // @[Switch.scala 41:52:@35947.4]
  assign output_59_55 = io_outValid_55 & _T_74788; // @[Switch.scala 41:38:@35948.4]
  assign _T_74791 = select_56 == 6'h3b; // @[Switch.scala 41:52:@35950.4]
  assign output_59_56 = io_outValid_56 & _T_74791; // @[Switch.scala 41:38:@35951.4]
  assign _T_74794 = select_57 == 6'h3b; // @[Switch.scala 41:52:@35953.4]
  assign output_59_57 = io_outValid_57 & _T_74794; // @[Switch.scala 41:38:@35954.4]
  assign _T_74797 = select_58 == 6'h3b; // @[Switch.scala 41:52:@35956.4]
  assign output_59_58 = io_outValid_58 & _T_74797; // @[Switch.scala 41:38:@35957.4]
  assign _T_74800 = select_59 == 6'h3b; // @[Switch.scala 41:52:@35959.4]
  assign output_59_59 = io_outValid_59 & _T_74800; // @[Switch.scala 41:38:@35960.4]
  assign _T_74803 = select_60 == 6'h3b; // @[Switch.scala 41:52:@35962.4]
  assign output_59_60 = io_outValid_60 & _T_74803; // @[Switch.scala 41:38:@35963.4]
  assign _T_74806 = select_61 == 6'h3b; // @[Switch.scala 41:52:@35965.4]
  assign output_59_61 = io_outValid_61 & _T_74806; // @[Switch.scala 41:38:@35966.4]
  assign _T_74809 = select_62 == 6'h3b; // @[Switch.scala 41:52:@35968.4]
  assign output_59_62 = io_outValid_62 & _T_74809; // @[Switch.scala 41:38:@35969.4]
  assign _T_74812 = select_63 == 6'h3b; // @[Switch.scala 41:52:@35971.4]
  assign output_59_63 = io_outValid_63 & _T_74812; // @[Switch.scala 41:38:@35972.4]
  assign _T_74820 = {output_59_7,output_59_6,output_59_5,output_59_4,output_59_3,output_59_2,output_59_1,output_59_0}; // @[Switch.scala 43:31:@35980.4]
  assign _T_74828 = {output_59_15,output_59_14,output_59_13,output_59_12,output_59_11,output_59_10,output_59_9,output_59_8,_T_74820}; // @[Switch.scala 43:31:@35988.4]
  assign _T_74835 = {output_59_23,output_59_22,output_59_21,output_59_20,output_59_19,output_59_18,output_59_17,output_59_16}; // @[Switch.scala 43:31:@35995.4]
  assign _T_74844 = {output_59_31,output_59_30,output_59_29,output_59_28,output_59_27,output_59_26,output_59_25,output_59_24,_T_74835,_T_74828}; // @[Switch.scala 43:31:@36004.4]
  assign _T_74851 = {output_59_39,output_59_38,output_59_37,output_59_36,output_59_35,output_59_34,output_59_33,output_59_32}; // @[Switch.scala 43:31:@36011.4]
  assign _T_74859 = {output_59_47,output_59_46,output_59_45,output_59_44,output_59_43,output_59_42,output_59_41,output_59_40,_T_74851}; // @[Switch.scala 43:31:@36019.4]
  assign _T_74866 = {output_59_55,output_59_54,output_59_53,output_59_52,output_59_51,output_59_50,output_59_49,output_59_48}; // @[Switch.scala 43:31:@36026.4]
  assign _T_74875 = {output_59_63,output_59_62,output_59_61,output_59_60,output_59_59,output_59_58,output_59_57,output_59_56,_T_74866,_T_74859}; // @[Switch.scala 43:31:@36035.4]
  assign _T_74876 = {_T_74875,_T_74844}; // @[Switch.scala 43:31:@36036.4]
  assign _T_74880 = select_0 == 6'h3c; // @[Switch.scala 41:52:@36039.4]
  assign output_60_0 = io_outValid_0 & _T_74880; // @[Switch.scala 41:38:@36040.4]
  assign _T_74883 = select_1 == 6'h3c; // @[Switch.scala 41:52:@36042.4]
  assign output_60_1 = io_outValid_1 & _T_74883; // @[Switch.scala 41:38:@36043.4]
  assign _T_74886 = select_2 == 6'h3c; // @[Switch.scala 41:52:@36045.4]
  assign output_60_2 = io_outValid_2 & _T_74886; // @[Switch.scala 41:38:@36046.4]
  assign _T_74889 = select_3 == 6'h3c; // @[Switch.scala 41:52:@36048.4]
  assign output_60_3 = io_outValid_3 & _T_74889; // @[Switch.scala 41:38:@36049.4]
  assign _T_74892 = select_4 == 6'h3c; // @[Switch.scala 41:52:@36051.4]
  assign output_60_4 = io_outValid_4 & _T_74892; // @[Switch.scala 41:38:@36052.4]
  assign _T_74895 = select_5 == 6'h3c; // @[Switch.scala 41:52:@36054.4]
  assign output_60_5 = io_outValid_5 & _T_74895; // @[Switch.scala 41:38:@36055.4]
  assign _T_74898 = select_6 == 6'h3c; // @[Switch.scala 41:52:@36057.4]
  assign output_60_6 = io_outValid_6 & _T_74898; // @[Switch.scala 41:38:@36058.4]
  assign _T_74901 = select_7 == 6'h3c; // @[Switch.scala 41:52:@36060.4]
  assign output_60_7 = io_outValid_7 & _T_74901; // @[Switch.scala 41:38:@36061.4]
  assign _T_74904 = select_8 == 6'h3c; // @[Switch.scala 41:52:@36063.4]
  assign output_60_8 = io_outValid_8 & _T_74904; // @[Switch.scala 41:38:@36064.4]
  assign _T_74907 = select_9 == 6'h3c; // @[Switch.scala 41:52:@36066.4]
  assign output_60_9 = io_outValid_9 & _T_74907; // @[Switch.scala 41:38:@36067.4]
  assign _T_74910 = select_10 == 6'h3c; // @[Switch.scala 41:52:@36069.4]
  assign output_60_10 = io_outValid_10 & _T_74910; // @[Switch.scala 41:38:@36070.4]
  assign _T_74913 = select_11 == 6'h3c; // @[Switch.scala 41:52:@36072.4]
  assign output_60_11 = io_outValid_11 & _T_74913; // @[Switch.scala 41:38:@36073.4]
  assign _T_74916 = select_12 == 6'h3c; // @[Switch.scala 41:52:@36075.4]
  assign output_60_12 = io_outValid_12 & _T_74916; // @[Switch.scala 41:38:@36076.4]
  assign _T_74919 = select_13 == 6'h3c; // @[Switch.scala 41:52:@36078.4]
  assign output_60_13 = io_outValid_13 & _T_74919; // @[Switch.scala 41:38:@36079.4]
  assign _T_74922 = select_14 == 6'h3c; // @[Switch.scala 41:52:@36081.4]
  assign output_60_14 = io_outValid_14 & _T_74922; // @[Switch.scala 41:38:@36082.4]
  assign _T_74925 = select_15 == 6'h3c; // @[Switch.scala 41:52:@36084.4]
  assign output_60_15 = io_outValid_15 & _T_74925; // @[Switch.scala 41:38:@36085.4]
  assign _T_74928 = select_16 == 6'h3c; // @[Switch.scala 41:52:@36087.4]
  assign output_60_16 = io_outValid_16 & _T_74928; // @[Switch.scala 41:38:@36088.4]
  assign _T_74931 = select_17 == 6'h3c; // @[Switch.scala 41:52:@36090.4]
  assign output_60_17 = io_outValid_17 & _T_74931; // @[Switch.scala 41:38:@36091.4]
  assign _T_74934 = select_18 == 6'h3c; // @[Switch.scala 41:52:@36093.4]
  assign output_60_18 = io_outValid_18 & _T_74934; // @[Switch.scala 41:38:@36094.4]
  assign _T_74937 = select_19 == 6'h3c; // @[Switch.scala 41:52:@36096.4]
  assign output_60_19 = io_outValid_19 & _T_74937; // @[Switch.scala 41:38:@36097.4]
  assign _T_74940 = select_20 == 6'h3c; // @[Switch.scala 41:52:@36099.4]
  assign output_60_20 = io_outValid_20 & _T_74940; // @[Switch.scala 41:38:@36100.4]
  assign _T_74943 = select_21 == 6'h3c; // @[Switch.scala 41:52:@36102.4]
  assign output_60_21 = io_outValid_21 & _T_74943; // @[Switch.scala 41:38:@36103.4]
  assign _T_74946 = select_22 == 6'h3c; // @[Switch.scala 41:52:@36105.4]
  assign output_60_22 = io_outValid_22 & _T_74946; // @[Switch.scala 41:38:@36106.4]
  assign _T_74949 = select_23 == 6'h3c; // @[Switch.scala 41:52:@36108.4]
  assign output_60_23 = io_outValid_23 & _T_74949; // @[Switch.scala 41:38:@36109.4]
  assign _T_74952 = select_24 == 6'h3c; // @[Switch.scala 41:52:@36111.4]
  assign output_60_24 = io_outValid_24 & _T_74952; // @[Switch.scala 41:38:@36112.4]
  assign _T_74955 = select_25 == 6'h3c; // @[Switch.scala 41:52:@36114.4]
  assign output_60_25 = io_outValid_25 & _T_74955; // @[Switch.scala 41:38:@36115.4]
  assign _T_74958 = select_26 == 6'h3c; // @[Switch.scala 41:52:@36117.4]
  assign output_60_26 = io_outValid_26 & _T_74958; // @[Switch.scala 41:38:@36118.4]
  assign _T_74961 = select_27 == 6'h3c; // @[Switch.scala 41:52:@36120.4]
  assign output_60_27 = io_outValid_27 & _T_74961; // @[Switch.scala 41:38:@36121.4]
  assign _T_74964 = select_28 == 6'h3c; // @[Switch.scala 41:52:@36123.4]
  assign output_60_28 = io_outValid_28 & _T_74964; // @[Switch.scala 41:38:@36124.4]
  assign _T_74967 = select_29 == 6'h3c; // @[Switch.scala 41:52:@36126.4]
  assign output_60_29 = io_outValid_29 & _T_74967; // @[Switch.scala 41:38:@36127.4]
  assign _T_74970 = select_30 == 6'h3c; // @[Switch.scala 41:52:@36129.4]
  assign output_60_30 = io_outValid_30 & _T_74970; // @[Switch.scala 41:38:@36130.4]
  assign _T_74973 = select_31 == 6'h3c; // @[Switch.scala 41:52:@36132.4]
  assign output_60_31 = io_outValid_31 & _T_74973; // @[Switch.scala 41:38:@36133.4]
  assign _T_74976 = select_32 == 6'h3c; // @[Switch.scala 41:52:@36135.4]
  assign output_60_32 = io_outValid_32 & _T_74976; // @[Switch.scala 41:38:@36136.4]
  assign _T_74979 = select_33 == 6'h3c; // @[Switch.scala 41:52:@36138.4]
  assign output_60_33 = io_outValid_33 & _T_74979; // @[Switch.scala 41:38:@36139.4]
  assign _T_74982 = select_34 == 6'h3c; // @[Switch.scala 41:52:@36141.4]
  assign output_60_34 = io_outValid_34 & _T_74982; // @[Switch.scala 41:38:@36142.4]
  assign _T_74985 = select_35 == 6'h3c; // @[Switch.scala 41:52:@36144.4]
  assign output_60_35 = io_outValid_35 & _T_74985; // @[Switch.scala 41:38:@36145.4]
  assign _T_74988 = select_36 == 6'h3c; // @[Switch.scala 41:52:@36147.4]
  assign output_60_36 = io_outValid_36 & _T_74988; // @[Switch.scala 41:38:@36148.4]
  assign _T_74991 = select_37 == 6'h3c; // @[Switch.scala 41:52:@36150.4]
  assign output_60_37 = io_outValid_37 & _T_74991; // @[Switch.scala 41:38:@36151.4]
  assign _T_74994 = select_38 == 6'h3c; // @[Switch.scala 41:52:@36153.4]
  assign output_60_38 = io_outValid_38 & _T_74994; // @[Switch.scala 41:38:@36154.4]
  assign _T_74997 = select_39 == 6'h3c; // @[Switch.scala 41:52:@36156.4]
  assign output_60_39 = io_outValid_39 & _T_74997; // @[Switch.scala 41:38:@36157.4]
  assign _T_75000 = select_40 == 6'h3c; // @[Switch.scala 41:52:@36159.4]
  assign output_60_40 = io_outValid_40 & _T_75000; // @[Switch.scala 41:38:@36160.4]
  assign _T_75003 = select_41 == 6'h3c; // @[Switch.scala 41:52:@36162.4]
  assign output_60_41 = io_outValid_41 & _T_75003; // @[Switch.scala 41:38:@36163.4]
  assign _T_75006 = select_42 == 6'h3c; // @[Switch.scala 41:52:@36165.4]
  assign output_60_42 = io_outValid_42 & _T_75006; // @[Switch.scala 41:38:@36166.4]
  assign _T_75009 = select_43 == 6'h3c; // @[Switch.scala 41:52:@36168.4]
  assign output_60_43 = io_outValid_43 & _T_75009; // @[Switch.scala 41:38:@36169.4]
  assign _T_75012 = select_44 == 6'h3c; // @[Switch.scala 41:52:@36171.4]
  assign output_60_44 = io_outValid_44 & _T_75012; // @[Switch.scala 41:38:@36172.4]
  assign _T_75015 = select_45 == 6'h3c; // @[Switch.scala 41:52:@36174.4]
  assign output_60_45 = io_outValid_45 & _T_75015; // @[Switch.scala 41:38:@36175.4]
  assign _T_75018 = select_46 == 6'h3c; // @[Switch.scala 41:52:@36177.4]
  assign output_60_46 = io_outValid_46 & _T_75018; // @[Switch.scala 41:38:@36178.4]
  assign _T_75021 = select_47 == 6'h3c; // @[Switch.scala 41:52:@36180.4]
  assign output_60_47 = io_outValid_47 & _T_75021; // @[Switch.scala 41:38:@36181.4]
  assign _T_75024 = select_48 == 6'h3c; // @[Switch.scala 41:52:@36183.4]
  assign output_60_48 = io_outValid_48 & _T_75024; // @[Switch.scala 41:38:@36184.4]
  assign _T_75027 = select_49 == 6'h3c; // @[Switch.scala 41:52:@36186.4]
  assign output_60_49 = io_outValid_49 & _T_75027; // @[Switch.scala 41:38:@36187.4]
  assign _T_75030 = select_50 == 6'h3c; // @[Switch.scala 41:52:@36189.4]
  assign output_60_50 = io_outValid_50 & _T_75030; // @[Switch.scala 41:38:@36190.4]
  assign _T_75033 = select_51 == 6'h3c; // @[Switch.scala 41:52:@36192.4]
  assign output_60_51 = io_outValid_51 & _T_75033; // @[Switch.scala 41:38:@36193.4]
  assign _T_75036 = select_52 == 6'h3c; // @[Switch.scala 41:52:@36195.4]
  assign output_60_52 = io_outValid_52 & _T_75036; // @[Switch.scala 41:38:@36196.4]
  assign _T_75039 = select_53 == 6'h3c; // @[Switch.scala 41:52:@36198.4]
  assign output_60_53 = io_outValid_53 & _T_75039; // @[Switch.scala 41:38:@36199.4]
  assign _T_75042 = select_54 == 6'h3c; // @[Switch.scala 41:52:@36201.4]
  assign output_60_54 = io_outValid_54 & _T_75042; // @[Switch.scala 41:38:@36202.4]
  assign _T_75045 = select_55 == 6'h3c; // @[Switch.scala 41:52:@36204.4]
  assign output_60_55 = io_outValid_55 & _T_75045; // @[Switch.scala 41:38:@36205.4]
  assign _T_75048 = select_56 == 6'h3c; // @[Switch.scala 41:52:@36207.4]
  assign output_60_56 = io_outValid_56 & _T_75048; // @[Switch.scala 41:38:@36208.4]
  assign _T_75051 = select_57 == 6'h3c; // @[Switch.scala 41:52:@36210.4]
  assign output_60_57 = io_outValid_57 & _T_75051; // @[Switch.scala 41:38:@36211.4]
  assign _T_75054 = select_58 == 6'h3c; // @[Switch.scala 41:52:@36213.4]
  assign output_60_58 = io_outValid_58 & _T_75054; // @[Switch.scala 41:38:@36214.4]
  assign _T_75057 = select_59 == 6'h3c; // @[Switch.scala 41:52:@36216.4]
  assign output_60_59 = io_outValid_59 & _T_75057; // @[Switch.scala 41:38:@36217.4]
  assign _T_75060 = select_60 == 6'h3c; // @[Switch.scala 41:52:@36219.4]
  assign output_60_60 = io_outValid_60 & _T_75060; // @[Switch.scala 41:38:@36220.4]
  assign _T_75063 = select_61 == 6'h3c; // @[Switch.scala 41:52:@36222.4]
  assign output_60_61 = io_outValid_61 & _T_75063; // @[Switch.scala 41:38:@36223.4]
  assign _T_75066 = select_62 == 6'h3c; // @[Switch.scala 41:52:@36225.4]
  assign output_60_62 = io_outValid_62 & _T_75066; // @[Switch.scala 41:38:@36226.4]
  assign _T_75069 = select_63 == 6'h3c; // @[Switch.scala 41:52:@36228.4]
  assign output_60_63 = io_outValid_63 & _T_75069; // @[Switch.scala 41:38:@36229.4]
  assign _T_75077 = {output_60_7,output_60_6,output_60_5,output_60_4,output_60_3,output_60_2,output_60_1,output_60_0}; // @[Switch.scala 43:31:@36237.4]
  assign _T_75085 = {output_60_15,output_60_14,output_60_13,output_60_12,output_60_11,output_60_10,output_60_9,output_60_8,_T_75077}; // @[Switch.scala 43:31:@36245.4]
  assign _T_75092 = {output_60_23,output_60_22,output_60_21,output_60_20,output_60_19,output_60_18,output_60_17,output_60_16}; // @[Switch.scala 43:31:@36252.4]
  assign _T_75101 = {output_60_31,output_60_30,output_60_29,output_60_28,output_60_27,output_60_26,output_60_25,output_60_24,_T_75092,_T_75085}; // @[Switch.scala 43:31:@36261.4]
  assign _T_75108 = {output_60_39,output_60_38,output_60_37,output_60_36,output_60_35,output_60_34,output_60_33,output_60_32}; // @[Switch.scala 43:31:@36268.4]
  assign _T_75116 = {output_60_47,output_60_46,output_60_45,output_60_44,output_60_43,output_60_42,output_60_41,output_60_40,_T_75108}; // @[Switch.scala 43:31:@36276.4]
  assign _T_75123 = {output_60_55,output_60_54,output_60_53,output_60_52,output_60_51,output_60_50,output_60_49,output_60_48}; // @[Switch.scala 43:31:@36283.4]
  assign _T_75132 = {output_60_63,output_60_62,output_60_61,output_60_60,output_60_59,output_60_58,output_60_57,output_60_56,_T_75123,_T_75116}; // @[Switch.scala 43:31:@36292.4]
  assign _T_75133 = {_T_75132,_T_75101}; // @[Switch.scala 43:31:@36293.4]
  assign _T_75137 = select_0 == 6'h3d; // @[Switch.scala 41:52:@36296.4]
  assign output_61_0 = io_outValid_0 & _T_75137; // @[Switch.scala 41:38:@36297.4]
  assign _T_75140 = select_1 == 6'h3d; // @[Switch.scala 41:52:@36299.4]
  assign output_61_1 = io_outValid_1 & _T_75140; // @[Switch.scala 41:38:@36300.4]
  assign _T_75143 = select_2 == 6'h3d; // @[Switch.scala 41:52:@36302.4]
  assign output_61_2 = io_outValid_2 & _T_75143; // @[Switch.scala 41:38:@36303.4]
  assign _T_75146 = select_3 == 6'h3d; // @[Switch.scala 41:52:@36305.4]
  assign output_61_3 = io_outValid_3 & _T_75146; // @[Switch.scala 41:38:@36306.4]
  assign _T_75149 = select_4 == 6'h3d; // @[Switch.scala 41:52:@36308.4]
  assign output_61_4 = io_outValid_4 & _T_75149; // @[Switch.scala 41:38:@36309.4]
  assign _T_75152 = select_5 == 6'h3d; // @[Switch.scala 41:52:@36311.4]
  assign output_61_5 = io_outValid_5 & _T_75152; // @[Switch.scala 41:38:@36312.4]
  assign _T_75155 = select_6 == 6'h3d; // @[Switch.scala 41:52:@36314.4]
  assign output_61_6 = io_outValid_6 & _T_75155; // @[Switch.scala 41:38:@36315.4]
  assign _T_75158 = select_7 == 6'h3d; // @[Switch.scala 41:52:@36317.4]
  assign output_61_7 = io_outValid_7 & _T_75158; // @[Switch.scala 41:38:@36318.4]
  assign _T_75161 = select_8 == 6'h3d; // @[Switch.scala 41:52:@36320.4]
  assign output_61_8 = io_outValid_8 & _T_75161; // @[Switch.scala 41:38:@36321.4]
  assign _T_75164 = select_9 == 6'h3d; // @[Switch.scala 41:52:@36323.4]
  assign output_61_9 = io_outValid_9 & _T_75164; // @[Switch.scala 41:38:@36324.4]
  assign _T_75167 = select_10 == 6'h3d; // @[Switch.scala 41:52:@36326.4]
  assign output_61_10 = io_outValid_10 & _T_75167; // @[Switch.scala 41:38:@36327.4]
  assign _T_75170 = select_11 == 6'h3d; // @[Switch.scala 41:52:@36329.4]
  assign output_61_11 = io_outValid_11 & _T_75170; // @[Switch.scala 41:38:@36330.4]
  assign _T_75173 = select_12 == 6'h3d; // @[Switch.scala 41:52:@36332.4]
  assign output_61_12 = io_outValid_12 & _T_75173; // @[Switch.scala 41:38:@36333.4]
  assign _T_75176 = select_13 == 6'h3d; // @[Switch.scala 41:52:@36335.4]
  assign output_61_13 = io_outValid_13 & _T_75176; // @[Switch.scala 41:38:@36336.4]
  assign _T_75179 = select_14 == 6'h3d; // @[Switch.scala 41:52:@36338.4]
  assign output_61_14 = io_outValid_14 & _T_75179; // @[Switch.scala 41:38:@36339.4]
  assign _T_75182 = select_15 == 6'h3d; // @[Switch.scala 41:52:@36341.4]
  assign output_61_15 = io_outValid_15 & _T_75182; // @[Switch.scala 41:38:@36342.4]
  assign _T_75185 = select_16 == 6'h3d; // @[Switch.scala 41:52:@36344.4]
  assign output_61_16 = io_outValid_16 & _T_75185; // @[Switch.scala 41:38:@36345.4]
  assign _T_75188 = select_17 == 6'h3d; // @[Switch.scala 41:52:@36347.4]
  assign output_61_17 = io_outValid_17 & _T_75188; // @[Switch.scala 41:38:@36348.4]
  assign _T_75191 = select_18 == 6'h3d; // @[Switch.scala 41:52:@36350.4]
  assign output_61_18 = io_outValid_18 & _T_75191; // @[Switch.scala 41:38:@36351.4]
  assign _T_75194 = select_19 == 6'h3d; // @[Switch.scala 41:52:@36353.4]
  assign output_61_19 = io_outValid_19 & _T_75194; // @[Switch.scala 41:38:@36354.4]
  assign _T_75197 = select_20 == 6'h3d; // @[Switch.scala 41:52:@36356.4]
  assign output_61_20 = io_outValid_20 & _T_75197; // @[Switch.scala 41:38:@36357.4]
  assign _T_75200 = select_21 == 6'h3d; // @[Switch.scala 41:52:@36359.4]
  assign output_61_21 = io_outValid_21 & _T_75200; // @[Switch.scala 41:38:@36360.4]
  assign _T_75203 = select_22 == 6'h3d; // @[Switch.scala 41:52:@36362.4]
  assign output_61_22 = io_outValid_22 & _T_75203; // @[Switch.scala 41:38:@36363.4]
  assign _T_75206 = select_23 == 6'h3d; // @[Switch.scala 41:52:@36365.4]
  assign output_61_23 = io_outValid_23 & _T_75206; // @[Switch.scala 41:38:@36366.4]
  assign _T_75209 = select_24 == 6'h3d; // @[Switch.scala 41:52:@36368.4]
  assign output_61_24 = io_outValid_24 & _T_75209; // @[Switch.scala 41:38:@36369.4]
  assign _T_75212 = select_25 == 6'h3d; // @[Switch.scala 41:52:@36371.4]
  assign output_61_25 = io_outValid_25 & _T_75212; // @[Switch.scala 41:38:@36372.4]
  assign _T_75215 = select_26 == 6'h3d; // @[Switch.scala 41:52:@36374.4]
  assign output_61_26 = io_outValid_26 & _T_75215; // @[Switch.scala 41:38:@36375.4]
  assign _T_75218 = select_27 == 6'h3d; // @[Switch.scala 41:52:@36377.4]
  assign output_61_27 = io_outValid_27 & _T_75218; // @[Switch.scala 41:38:@36378.4]
  assign _T_75221 = select_28 == 6'h3d; // @[Switch.scala 41:52:@36380.4]
  assign output_61_28 = io_outValid_28 & _T_75221; // @[Switch.scala 41:38:@36381.4]
  assign _T_75224 = select_29 == 6'h3d; // @[Switch.scala 41:52:@36383.4]
  assign output_61_29 = io_outValid_29 & _T_75224; // @[Switch.scala 41:38:@36384.4]
  assign _T_75227 = select_30 == 6'h3d; // @[Switch.scala 41:52:@36386.4]
  assign output_61_30 = io_outValid_30 & _T_75227; // @[Switch.scala 41:38:@36387.4]
  assign _T_75230 = select_31 == 6'h3d; // @[Switch.scala 41:52:@36389.4]
  assign output_61_31 = io_outValid_31 & _T_75230; // @[Switch.scala 41:38:@36390.4]
  assign _T_75233 = select_32 == 6'h3d; // @[Switch.scala 41:52:@36392.4]
  assign output_61_32 = io_outValid_32 & _T_75233; // @[Switch.scala 41:38:@36393.4]
  assign _T_75236 = select_33 == 6'h3d; // @[Switch.scala 41:52:@36395.4]
  assign output_61_33 = io_outValid_33 & _T_75236; // @[Switch.scala 41:38:@36396.4]
  assign _T_75239 = select_34 == 6'h3d; // @[Switch.scala 41:52:@36398.4]
  assign output_61_34 = io_outValid_34 & _T_75239; // @[Switch.scala 41:38:@36399.4]
  assign _T_75242 = select_35 == 6'h3d; // @[Switch.scala 41:52:@36401.4]
  assign output_61_35 = io_outValid_35 & _T_75242; // @[Switch.scala 41:38:@36402.4]
  assign _T_75245 = select_36 == 6'h3d; // @[Switch.scala 41:52:@36404.4]
  assign output_61_36 = io_outValid_36 & _T_75245; // @[Switch.scala 41:38:@36405.4]
  assign _T_75248 = select_37 == 6'h3d; // @[Switch.scala 41:52:@36407.4]
  assign output_61_37 = io_outValid_37 & _T_75248; // @[Switch.scala 41:38:@36408.4]
  assign _T_75251 = select_38 == 6'h3d; // @[Switch.scala 41:52:@36410.4]
  assign output_61_38 = io_outValid_38 & _T_75251; // @[Switch.scala 41:38:@36411.4]
  assign _T_75254 = select_39 == 6'h3d; // @[Switch.scala 41:52:@36413.4]
  assign output_61_39 = io_outValid_39 & _T_75254; // @[Switch.scala 41:38:@36414.4]
  assign _T_75257 = select_40 == 6'h3d; // @[Switch.scala 41:52:@36416.4]
  assign output_61_40 = io_outValid_40 & _T_75257; // @[Switch.scala 41:38:@36417.4]
  assign _T_75260 = select_41 == 6'h3d; // @[Switch.scala 41:52:@36419.4]
  assign output_61_41 = io_outValid_41 & _T_75260; // @[Switch.scala 41:38:@36420.4]
  assign _T_75263 = select_42 == 6'h3d; // @[Switch.scala 41:52:@36422.4]
  assign output_61_42 = io_outValid_42 & _T_75263; // @[Switch.scala 41:38:@36423.4]
  assign _T_75266 = select_43 == 6'h3d; // @[Switch.scala 41:52:@36425.4]
  assign output_61_43 = io_outValid_43 & _T_75266; // @[Switch.scala 41:38:@36426.4]
  assign _T_75269 = select_44 == 6'h3d; // @[Switch.scala 41:52:@36428.4]
  assign output_61_44 = io_outValid_44 & _T_75269; // @[Switch.scala 41:38:@36429.4]
  assign _T_75272 = select_45 == 6'h3d; // @[Switch.scala 41:52:@36431.4]
  assign output_61_45 = io_outValid_45 & _T_75272; // @[Switch.scala 41:38:@36432.4]
  assign _T_75275 = select_46 == 6'h3d; // @[Switch.scala 41:52:@36434.4]
  assign output_61_46 = io_outValid_46 & _T_75275; // @[Switch.scala 41:38:@36435.4]
  assign _T_75278 = select_47 == 6'h3d; // @[Switch.scala 41:52:@36437.4]
  assign output_61_47 = io_outValid_47 & _T_75278; // @[Switch.scala 41:38:@36438.4]
  assign _T_75281 = select_48 == 6'h3d; // @[Switch.scala 41:52:@36440.4]
  assign output_61_48 = io_outValid_48 & _T_75281; // @[Switch.scala 41:38:@36441.4]
  assign _T_75284 = select_49 == 6'h3d; // @[Switch.scala 41:52:@36443.4]
  assign output_61_49 = io_outValid_49 & _T_75284; // @[Switch.scala 41:38:@36444.4]
  assign _T_75287 = select_50 == 6'h3d; // @[Switch.scala 41:52:@36446.4]
  assign output_61_50 = io_outValid_50 & _T_75287; // @[Switch.scala 41:38:@36447.4]
  assign _T_75290 = select_51 == 6'h3d; // @[Switch.scala 41:52:@36449.4]
  assign output_61_51 = io_outValid_51 & _T_75290; // @[Switch.scala 41:38:@36450.4]
  assign _T_75293 = select_52 == 6'h3d; // @[Switch.scala 41:52:@36452.4]
  assign output_61_52 = io_outValid_52 & _T_75293; // @[Switch.scala 41:38:@36453.4]
  assign _T_75296 = select_53 == 6'h3d; // @[Switch.scala 41:52:@36455.4]
  assign output_61_53 = io_outValid_53 & _T_75296; // @[Switch.scala 41:38:@36456.4]
  assign _T_75299 = select_54 == 6'h3d; // @[Switch.scala 41:52:@36458.4]
  assign output_61_54 = io_outValid_54 & _T_75299; // @[Switch.scala 41:38:@36459.4]
  assign _T_75302 = select_55 == 6'h3d; // @[Switch.scala 41:52:@36461.4]
  assign output_61_55 = io_outValid_55 & _T_75302; // @[Switch.scala 41:38:@36462.4]
  assign _T_75305 = select_56 == 6'h3d; // @[Switch.scala 41:52:@36464.4]
  assign output_61_56 = io_outValid_56 & _T_75305; // @[Switch.scala 41:38:@36465.4]
  assign _T_75308 = select_57 == 6'h3d; // @[Switch.scala 41:52:@36467.4]
  assign output_61_57 = io_outValid_57 & _T_75308; // @[Switch.scala 41:38:@36468.4]
  assign _T_75311 = select_58 == 6'h3d; // @[Switch.scala 41:52:@36470.4]
  assign output_61_58 = io_outValid_58 & _T_75311; // @[Switch.scala 41:38:@36471.4]
  assign _T_75314 = select_59 == 6'h3d; // @[Switch.scala 41:52:@36473.4]
  assign output_61_59 = io_outValid_59 & _T_75314; // @[Switch.scala 41:38:@36474.4]
  assign _T_75317 = select_60 == 6'h3d; // @[Switch.scala 41:52:@36476.4]
  assign output_61_60 = io_outValid_60 & _T_75317; // @[Switch.scala 41:38:@36477.4]
  assign _T_75320 = select_61 == 6'h3d; // @[Switch.scala 41:52:@36479.4]
  assign output_61_61 = io_outValid_61 & _T_75320; // @[Switch.scala 41:38:@36480.4]
  assign _T_75323 = select_62 == 6'h3d; // @[Switch.scala 41:52:@36482.4]
  assign output_61_62 = io_outValid_62 & _T_75323; // @[Switch.scala 41:38:@36483.4]
  assign _T_75326 = select_63 == 6'h3d; // @[Switch.scala 41:52:@36485.4]
  assign output_61_63 = io_outValid_63 & _T_75326; // @[Switch.scala 41:38:@36486.4]
  assign _T_75334 = {output_61_7,output_61_6,output_61_5,output_61_4,output_61_3,output_61_2,output_61_1,output_61_0}; // @[Switch.scala 43:31:@36494.4]
  assign _T_75342 = {output_61_15,output_61_14,output_61_13,output_61_12,output_61_11,output_61_10,output_61_9,output_61_8,_T_75334}; // @[Switch.scala 43:31:@36502.4]
  assign _T_75349 = {output_61_23,output_61_22,output_61_21,output_61_20,output_61_19,output_61_18,output_61_17,output_61_16}; // @[Switch.scala 43:31:@36509.4]
  assign _T_75358 = {output_61_31,output_61_30,output_61_29,output_61_28,output_61_27,output_61_26,output_61_25,output_61_24,_T_75349,_T_75342}; // @[Switch.scala 43:31:@36518.4]
  assign _T_75365 = {output_61_39,output_61_38,output_61_37,output_61_36,output_61_35,output_61_34,output_61_33,output_61_32}; // @[Switch.scala 43:31:@36525.4]
  assign _T_75373 = {output_61_47,output_61_46,output_61_45,output_61_44,output_61_43,output_61_42,output_61_41,output_61_40,_T_75365}; // @[Switch.scala 43:31:@36533.4]
  assign _T_75380 = {output_61_55,output_61_54,output_61_53,output_61_52,output_61_51,output_61_50,output_61_49,output_61_48}; // @[Switch.scala 43:31:@36540.4]
  assign _T_75389 = {output_61_63,output_61_62,output_61_61,output_61_60,output_61_59,output_61_58,output_61_57,output_61_56,_T_75380,_T_75373}; // @[Switch.scala 43:31:@36549.4]
  assign _T_75390 = {_T_75389,_T_75358}; // @[Switch.scala 43:31:@36550.4]
  assign _T_75394 = select_0 == 6'h3e; // @[Switch.scala 41:52:@36553.4]
  assign output_62_0 = io_outValid_0 & _T_75394; // @[Switch.scala 41:38:@36554.4]
  assign _T_75397 = select_1 == 6'h3e; // @[Switch.scala 41:52:@36556.4]
  assign output_62_1 = io_outValid_1 & _T_75397; // @[Switch.scala 41:38:@36557.4]
  assign _T_75400 = select_2 == 6'h3e; // @[Switch.scala 41:52:@36559.4]
  assign output_62_2 = io_outValid_2 & _T_75400; // @[Switch.scala 41:38:@36560.4]
  assign _T_75403 = select_3 == 6'h3e; // @[Switch.scala 41:52:@36562.4]
  assign output_62_3 = io_outValid_3 & _T_75403; // @[Switch.scala 41:38:@36563.4]
  assign _T_75406 = select_4 == 6'h3e; // @[Switch.scala 41:52:@36565.4]
  assign output_62_4 = io_outValid_4 & _T_75406; // @[Switch.scala 41:38:@36566.4]
  assign _T_75409 = select_5 == 6'h3e; // @[Switch.scala 41:52:@36568.4]
  assign output_62_5 = io_outValid_5 & _T_75409; // @[Switch.scala 41:38:@36569.4]
  assign _T_75412 = select_6 == 6'h3e; // @[Switch.scala 41:52:@36571.4]
  assign output_62_6 = io_outValid_6 & _T_75412; // @[Switch.scala 41:38:@36572.4]
  assign _T_75415 = select_7 == 6'h3e; // @[Switch.scala 41:52:@36574.4]
  assign output_62_7 = io_outValid_7 & _T_75415; // @[Switch.scala 41:38:@36575.4]
  assign _T_75418 = select_8 == 6'h3e; // @[Switch.scala 41:52:@36577.4]
  assign output_62_8 = io_outValid_8 & _T_75418; // @[Switch.scala 41:38:@36578.4]
  assign _T_75421 = select_9 == 6'h3e; // @[Switch.scala 41:52:@36580.4]
  assign output_62_9 = io_outValid_9 & _T_75421; // @[Switch.scala 41:38:@36581.4]
  assign _T_75424 = select_10 == 6'h3e; // @[Switch.scala 41:52:@36583.4]
  assign output_62_10 = io_outValid_10 & _T_75424; // @[Switch.scala 41:38:@36584.4]
  assign _T_75427 = select_11 == 6'h3e; // @[Switch.scala 41:52:@36586.4]
  assign output_62_11 = io_outValid_11 & _T_75427; // @[Switch.scala 41:38:@36587.4]
  assign _T_75430 = select_12 == 6'h3e; // @[Switch.scala 41:52:@36589.4]
  assign output_62_12 = io_outValid_12 & _T_75430; // @[Switch.scala 41:38:@36590.4]
  assign _T_75433 = select_13 == 6'h3e; // @[Switch.scala 41:52:@36592.4]
  assign output_62_13 = io_outValid_13 & _T_75433; // @[Switch.scala 41:38:@36593.4]
  assign _T_75436 = select_14 == 6'h3e; // @[Switch.scala 41:52:@36595.4]
  assign output_62_14 = io_outValid_14 & _T_75436; // @[Switch.scala 41:38:@36596.4]
  assign _T_75439 = select_15 == 6'h3e; // @[Switch.scala 41:52:@36598.4]
  assign output_62_15 = io_outValid_15 & _T_75439; // @[Switch.scala 41:38:@36599.4]
  assign _T_75442 = select_16 == 6'h3e; // @[Switch.scala 41:52:@36601.4]
  assign output_62_16 = io_outValid_16 & _T_75442; // @[Switch.scala 41:38:@36602.4]
  assign _T_75445 = select_17 == 6'h3e; // @[Switch.scala 41:52:@36604.4]
  assign output_62_17 = io_outValid_17 & _T_75445; // @[Switch.scala 41:38:@36605.4]
  assign _T_75448 = select_18 == 6'h3e; // @[Switch.scala 41:52:@36607.4]
  assign output_62_18 = io_outValid_18 & _T_75448; // @[Switch.scala 41:38:@36608.4]
  assign _T_75451 = select_19 == 6'h3e; // @[Switch.scala 41:52:@36610.4]
  assign output_62_19 = io_outValid_19 & _T_75451; // @[Switch.scala 41:38:@36611.4]
  assign _T_75454 = select_20 == 6'h3e; // @[Switch.scala 41:52:@36613.4]
  assign output_62_20 = io_outValid_20 & _T_75454; // @[Switch.scala 41:38:@36614.4]
  assign _T_75457 = select_21 == 6'h3e; // @[Switch.scala 41:52:@36616.4]
  assign output_62_21 = io_outValid_21 & _T_75457; // @[Switch.scala 41:38:@36617.4]
  assign _T_75460 = select_22 == 6'h3e; // @[Switch.scala 41:52:@36619.4]
  assign output_62_22 = io_outValid_22 & _T_75460; // @[Switch.scala 41:38:@36620.4]
  assign _T_75463 = select_23 == 6'h3e; // @[Switch.scala 41:52:@36622.4]
  assign output_62_23 = io_outValid_23 & _T_75463; // @[Switch.scala 41:38:@36623.4]
  assign _T_75466 = select_24 == 6'h3e; // @[Switch.scala 41:52:@36625.4]
  assign output_62_24 = io_outValid_24 & _T_75466; // @[Switch.scala 41:38:@36626.4]
  assign _T_75469 = select_25 == 6'h3e; // @[Switch.scala 41:52:@36628.4]
  assign output_62_25 = io_outValid_25 & _T_75469; // @[Switch.scala 41:38:@36629.4]
  assign _T_75472 = select_26 == 6'h3e; // @[Switch.scala 41:52:@36631.4]
  assign output_62_26 = io_outValid_26 & _T_75472; // @[Switch.scala 41:38:@36632.4]
  assign _T_75475 = select_27 == 6'h3e; // @[Switch.scala 41:52:@36634.4]
  assign output_62_27 = io_outValid_27 & _T_75475; // @[Switch.scala 41:38:@36635.4]
  assign _T_75478 = select_28 == 6'h3e; // @[Switch.scala 41:52:@36637.4]
  assign output_62_28 = io_outValid_28 & _T_75478; // @[Switch.scala 41:38:@36638.4]
  assign _T_75481 = select_29 == 6'h3e; // @[Switch.scala 41:52:@36640.4]
  assign output_62_29 = io_outValid_29 & _T_75481; // @[Switch.scala 41:38:@36641.4]
  assign _T_75484 = select_30 == 6'h3e; // @[Switch.scala 41:52:@36643.4]
  assign output_62_30 = io_outValid_30 & _T_75484; // @[Switch.scala 41:38:@36644.4]
  assign _T_75487 = select_31 == 6'h3e; // @[Switch.scala 41:52:@36646.4]
  assign output_62_31 = io_outValid_31 & _T_75487; // @[Switch.scala 41:38:@36647.4]
  assign _T_75490 = select_32 == 6'h3e; // @[Switch.scala 41:52:@36649.4]
  assign output_62_32 = io_outValid_32 & _T_75490; // @[Switch.scala 41:38:@36650.4]
  assign _T_75493 = select_33 == 6'h3e; // @[Switch.scala 41:52:@36652.4]
  assign output_62_33 = io_outValid_33 & _T_75493; // @[Switch.scala 41:38:@36653.4]
  assign _T_75496 = select_34 == 6'h3e; // @[Switch.scala 41:52:@36655.4]
  assign output_62_34 = io_outValid_34 & _T_75496; // @[Switch.scala 41:38:@36656.4]
  assign _T_75499 = select_35 == 6'h3e; // @[Switch.scala 41:52:@36658.4]
  assign output_62_35 = io_outValid_35 & _T_75499; // @[Switch.scala 41:38:@36659.4]
  assign _T_75502 = select_36 == 6'h3e; // @[Switch.scala 41:52:@36661.4]
  assign output_62_36 = io_outValid_36 & _T_75502; // @[Switch.scala 41:38:@36662.4]
  assign _T_75505 = select_37 == 6'h3e; // @[Switch.scala 41:52:@36664.4]
  assign output_62_37 = io_outValid_37 & _T_75505; // @[Switch.scala 41:38:@36665.4]
  assign _T_75508 = select_38 == 6'h3e; // @[Switch.scala 41:52:@36667.4]
  assign output_62_38 = io_outValid_38 & _T_75508; // @[Switch.scala 41:38:@36668.4]
  assign _T_75511 = select_39 == 6'h3e; // @[Switch.scala 41:52:@36670.4]
  assign output_62_39 = io_outValid_39 & _T_75511; // @[Switch.scala 41:38:@36671.4]
  assign _T_75514 = select_40 == 6'h3e; // @[Switch.scala 41:52:@36673.4]
  assign output_62_40 = io_outValid_40 & _T_75514; // @[Switch.scala 41:38:@36674.4]
  assign _T_75517 = select_41 == 6'h3e; // @[Switch.scala 41:52:@36676.4]
  assign output_62_41 = io_outValid_41 & _T_75517; // @[Switch.scala 41:38:@36677.4]
  assign _T_75520 = select_42 == 6'h3e; // @[Switch.scala 41:52:@36679.4]
  assign output_62_42 = io_outValid_42 & _T_75520; // @[Switch.scala 41:38:@36680.4]
  assign _T_75523 = select_43 == 6'h3e; // @[Switch.scala 41:52:@36682.4]
  assign output_62_43 = io_outValid_43 & _T_75523; // @[Switch.scala 41:38:@36683.4]
  assign _T_75526 = select_44 == 6'h3e; // @[Switch.scala 41:52:@36685.4]
  assign output_62_44 = io_outValid_44 & _T_75526; // @[Switch.scala 41:38:@36686.4]
  assign _T_75529 = select_45 == 6'h3e; // @[Switch.scala 41:52:@36688.4]
  assign output_62_45 = io_outValid_45 & _T_75529; // @[Switch.scala 41:38:@36689.4]
  assign _T_75532 = select_46 == 6'h3e; // @[Switch.scala 41:52:@36691.4]
  assign output_62_46 = io_outValid_46 & _T_75532; // @[Switch.scala 41:38:@36692.4]
  assign _T_75535 = select_47 == 6'h3e; // @[Switch.scala 41:52:@36694.4]
  assign output_62_47 = io_outValid_47 & _T_75535; // @[Switch.scala 41:38:@36695.4]
  assign _T_75538 = select_48 == 6'h3e; // @[Switch.scala 41:52:@36697.4]
  assign output_62_48 = io_outValid_48 & _T_75538; // @[Switch.scala 41:38:@36698.4]
  assign _T_75541 = select_49 == 6'h3e; // @[Switch.scala 41:52:@36700.4]
  assign output_62_49 = io_outValid_49 & _T_75541; // @[Switch.scala 41:38:@36701.4]
  assign _T_75544 = select_50 == 6'h3e; // @[Switch.scala 41:52:@36703.4]
  assign output_62_50 = io_outValid_50 & _T_75544; // @[Switch.scala 41:38:@36704.4]
  assign _T_75547 = select_51 == 6'h3e; // @[Switch.scala 41:52:@36706.4]
  assign output_62_51 = io_outValid_51 & _T_75547; // @[Switch.scala 41:38:@36707.4]
  assign _T_75550 = select_52 == 6'h3e; // @[Switch.scala 41:52:@36709.4]
  assign output_62_52 = io_outValid_52 & _T_75550; // @[Switch.scala 41:38:@36710.4]
  assign _T_75553 = select_53 == 6'h3e; // @[Switch.scala 41:52:@36712.4]
  assign output_62_53 = io_outValid_53 & _T_75553; // @[Switch.scala 41:38:@36713.4]
  assign _T_75556 = select_54 == 6'h3e; // @[Switch.scala 41:52:@36715.4]
  assign output_62_54 = io_outValid_54 & _T_75556; // @[Switch.scala 41:38:@36716.4]
  assign _T_75559 = select_55 == 6'h3e; // @[Switch.scala 41:52:@36718.4]
  assign output_62_55 = io_outValid_55 & _T_75559; // @[Switch.scala 41:38:@36719.4]
  assign _T_75562 = select_56 == 6'h3e; // @[Switch.scala 41:52:@36721.4]
  assign output_62_56 = io_outValid_56 & _T_75562; // @[Switch.scala 41:38:@36722.4]
  assign _T_75565 = select_57 == 6'h3e; // @[Switch.scala 41:52:@36724.4]
  assign output_62_57 = io_outValid_57 & _T_75565; // @[Switch.scala 41:38:@36725.4]
  assign _T_75568 = select_58 == 6'h3e; // @[Switch.scala 41:52:@36727.4]
  assign output_62_58 = io_outValid_58 & _T_75568; // @[Switch.scala 41:38:@36728.4]
  assign _T_75571 = select_59 == 6'h3e; // @[Switch.scala 41:52:@36730.4]
  assign output_62_59 = io_outValid_59 & _T_75571; // @[Switch.scala 41:38:@36731.4]
  assign _T_75574 = select_60 == 6'h3e; // @[Switch.scala 41:52:@36733.4]
  assign output_62_60 = io_outValid_60 & _T_75574; // @[Switch.scala 41:38:@36734.4]
  assign _T_75577 = select_61 == 6'h3e; // @[Switch.scala 41:52:@36736.4]
  assign output_62_61 = io_outValid_61 & _T_75577; // @[Switch.scala 41:38:@36737.4]
  assign _T_75580 = select_62 == 6'h3e; // @[Switch.scala 41:52:@36739.4]
  assign output_62_62 = io_outValid_62 & _T_75580; // @[Switch.scala 41:38:@36740.4]
  assign _T_75583 = select_63 == 6'h3e; // @[Switch.scala 41:52:@36742.4]
  assign output_62_63 = io_outValid_63 & _T_75583; // @[Switch.scala 41:38:@36743.4]
  assign _T_75591 = {output_62_7,output_62_6,output_62_5,output_62_4,output_62_3,output_62_2,output_62_1,output_62_0}; // @[Switch.scala 43:31:@36751.4]
  assign _T_75599 = {output_62_15,output_62_14,output_62_13,output_62_12,output_62_11,output_62_10,output_62_9,output_62_8,_T_75591}; // @[Switch.scala 43:31:@36759.4]
  assign _T_75606 = {output_62_23,output_62_22,output_62_21,output_62_20,output_62_19,output_62_18,output_62_17,output_62_16}; // @[Switch.scala 43:31:@36766.4]
  assign _T_75615 = {output_62_31,output_62_30,output_62_29,output_62_28,output_62_27,output_62_26,output_62_25,output_62_24,_T_75606,_T_75599}; // @[Switch.scala 43:31:@36775.4]
  assign _T_75622 = {output_62_39,output_62_38,output_62_37,output_62_36,output_62_35,output_62_34,output_62_33,output_62_32}; // @[Switch.scala 43:31:@36782.4]
  assign _T_75630 = {output_62_47,output_62_46,output_62_45,output_62_44,output_62_43,output_62_42,output_62_41,output_62_40,_T_75622}; // @[Switch.scala 43:31:@36790.4]
  assign _T_75637 = {output_62_55,output_62_54,output_62_53,output_62_52,output_62_51,output_62_50,output_62_49,output_62_48}; // @[Switch.scala 43:31:@36797.4]
  assign _T_75646 = {output_62_63,output_62_62,output_62_61,output_62_60,output_62_59,output_62_58,output_62_57,output_62_56,_T_75637,_T_75630}; // @[Switch.scala 43:31:@36806.4]
  assign _T_75647 = {_T_75646,_T_75615}; // @[Switch.scala 43:31:@36807.4]
  assign _T_75651 = select_0 == 6'h3f; // @[Switch.scala 41:52:@36810.4]
  assign output_63_0 = io_outValid_0 & _T_75651; // @[Switch.scala 41:38:@36811.4]
  assign _T_75654 = select_1 == 6'h3f; // @[Switch.scala 41:52:@36813.4]
  assign output_63_1 = io_outValid_1 & _T_75654; // @[Switch.scala 41:38:@36814.4]
  assign _T_75657 = select_2 == 6'h3f; // @[Switch.scala 41:52:@36816.4]
  assign output_63_2 = io_outValid_2 & _T_75657; // @[Switch.scala 41:38:@36817.4]
  assign _T_75660 = select_3 == 6'h3f; // @[Switch.scala 41:52:@36819.4]
  assign output_63_3 = io_outValid_3 & _T_75660; // @[Switch.scala 41:38:@36820.4]
  assign _T_75663 = select_4 == 6'h3f; // @[Switch.scala 41:52:@36822.4]
  assign output_63_4 = io_outValid_4 & _T_75663; // @[Switch.scala 41:38:@36823.4]
  assign _T_75666 = select_5 == 6'h3f; // @[Switch.scala 41:52:@36825.4]
  assign output_63_5 = io_outValid_5 & _T_75666; // @[Switch.scala 41:38:@36826.4]
  assign _T_75669 = select_6 == 6'h3f; // @[Switch.scala 41:52:@36828.4]
  assign output_63_6 = io_outValid_6 & _T_75669; // @[Switch.scala 41:38:@36829.4]
  assign _T_75672 = select_7 == 6'h3f; // @[Switch.scala 41:52:@36831.4]
  assign output_63_7 = io_outValid_7 & _T_75672; // @[Switch.scala 41:38:@36832.4]
  assign _T_75675 = select_8 == 6'h3f; // @[Switch.scala 41:52:@36834.4]
  assign output_63_8 = io_outValid_8 & _T_75675; // @[Switch.scala 41:38:@36835.4]
  assign _T_75678 = select_9 == 6'h3f; // @[Switch.scala 41:52:@36837.4]
  assign output_63_9 = io_outValid_9 & _T_75678; // @[Switch.scala 41:38:@36838.4]
  assign _T_75681 = select_10 == 6'h3f; // @[Switch.scala 41:52:@36840.4]
  assign output_63_10 = io_outValid_10 & _T_75681; // @[Switch.scala 41:38:@36841.4]
  assign _T_75684 = select_11 == 6'h3f; // @[Switch.scala 41:52:@36843.4]
  assign output_63_11 = io_outValid_11 & _T_75684; // @[Switch.scala 41:38:@36844.4]
  assign _T_75687 = select_12 == 6'h3f; // @[Switch.scala 41:52:@36846.4]
  assign output_63_12 = io_outValid_12 & _T_75687; // @[Switch.scala 41:38:@36847.4]
  assign _T_75690 = select_13 == 6'h3f; // @[Switch.scala 41:52:@36849.4]
  assign output_63_13 = io_outValid_13 & _T_75690; // @[Switch.scala 41:38:@36850.4]
  assign _T_75693 = select_14 == 6'h3f; // @[Switch.scala 41:52:@36852.4]
  assign output_63_14 = io_outValid_14 & _T_75693; // @[Switch.scala 41:38:@36853.4]
  assign _T_75696 = select_15 == 6'h3f; // @[Switch.scala 41:52:@36855.4]
  assign output_63_15 = io_outValid_15 & _T_75696; // @[Switch.scala 41:38:@36856.4]
  assign _T_75699 = select_16 == 6'h3f; // @[Switch.scala 41:52:@36858.4]
  assign output_63_16 = io_outValid_16 & _T_75699; // @[Switch.scala 41:38:@36859.4]
  assign _T_75702 = select_17 == 6'h3f; // @[Switch.scala 41:52:@36861.4]
  assign output_63_17 = io_outValid_17 & _T_75702; // @[Switch.scala 41:38:@36862.4]
  assign _T_75705 = select_18 == 6'h3f; // @[Switch.scala 41:52:@36864.4]
  assign output_63_18 = io_outValid_18 & _T_75705; // @[Switch.scala 41:38:@36865.4]
  assign _T_75708 = select_19 == 6'h3f; // @[Switch.scala 41:52:@36867.4]
  assign output_63_19 = io_outValid_19 & _T_75708; // @[Switch.scala 41:38:@36868.4]
  assign _T_75711 = select_20 == 6'h3f; // @[Switch.scala 41:52:@36870.4]
  assign output_63_20 = io_outValid_20 & _T_75711; // @[Switch.scala 41:38:@36871.4]
  assign _T_75714 = select_21 == 6'h3f; // @[Switch.scala 41:52:@36873.4]
  assign output_63_21 = io_outValid_21 & _T_75714; // @[Switch.scala 41:38:@36874.4]
  assign _T_75717 = select_22 == 6'h3f; // @[Switch.scala 41:52:@36876.4]
  assign output_63_22 = io_outValid_22 & _T_75717; // @[Switch.scala 41:38:@36877.4]
  assign _T_75720 = select_23 == 6'h3f; // @[Switch.scala 41:52:@36879.4]
  assign output_63_23 = io_outValid_23 & _T_75720; // @[Switch.scala 41:38:@36880.4]
  assign _T_75723 = select_24 == 6'h3f; // @[Switch.scala 41:52:@36882.4]
  assign output_63_24 = io_outValid_24 & _T_75723; // @[Switch.scala 41:38:@36883.4]
  assign _T_75726 = select_25 == 6'h3f; // @[Switch.scala 41:52:@36885.4]
  assign output_63_25 = io_outValid_25 & _T_75726; // @[Switch.scala 41:38:@36886.4]
  assign _T_75729 = select_26 == 6'h3f; // @[Switch.scala 41:52:@36888.4]
  assign output_63_26 = io_outValid_26 & _T_75729; // @[Switch.scala 41:38:@36889.4]
  assign _T_75732 = select_27 == 6'h3f; // @[Switch.scala 41:52:@36891.4]
  assign output_63_27 = io_outValid_27 & _T_75732; // @[Switch.scala 41:38:@36892.4]
  assign _T_75735 = select_28 == 6'h3f; // @[Switch.scala 41:52:@36894.4]
  assign output_63_28 = io_outValid_28 & _T_75735; // @[Switch.scala 41:38:@36895.4]
  assign _T_75738 = select_29 == 6'h3f; // @[Switch.scala 41:52:@36897.4]
  assign output_63_29 = io_outValid_29 & _T_75738; // @[Switch.scala 41:38:@36898.4]
  assign _T_75741 = select_30 == 6'h3f; // @[Switch.scala 41:52:@36900.4]
  assign output_63_30 = io_outValid_30 & _T_75741; // @[Switch.scala 41:38:@36901.4]
  assign _T_75744 = select_31 == 6'h3f; // @[Switch.scala 41:52:@36903.4]
  assign output_63_31 = io_outValid_31 & _T_75744; // @[Switch.scala 41:38:@36904.4]
  assign _T_75747 = select_32 == 6'h3f; // @[Switch.scala 41:52:@36906.4]
  assign output_63_32 = io_outValid_32 & _T_75747; // @[Switch.scala 41:38:@36907.4]
  assign _T_75750 = select_33 == 6'h3f; // @[Switch.scala 41:52:@36909.4]
  assign output_63_33 = io_outValid_33 & _T_75750; // @[Switch.scala 41:38:@36910.4]
  assign _T_75753 = select_34 == 6'h3f; // @[Switch.scala 41:52:@36912.4]
  assign output_63_34 = io_outValid_34 & _T_75753; // @[Switch.scala 41:38:@36913.4]
  assign _T_75756 = select_35 == 6'h3f; // @[Switch.scala 41:52:@36915.4]
  assign output_63_35 = io_outValid_35 & _T_75756; // @[Switch.scala 41:38:@36916.4]
  assign _T_75759 = select_36 == 6'h3f; // @[Switch.scala 41:52:@36918.4]
  assign output_63_36 = io_outValid_36 & _T_75759; // @[Switch.scala 41:38:@36919.4]
  assign _T_75762 = select_37 == 6'h3f; // @[Switch.scala 41:52:@36921.4]
  assign output_63_37 = io_outValid_37 & _T_75762; // @[Switch.scala 41:38:@36922.4]
  assign _T_75765 = select_38 == 6'h3f; // @[Switch.scala 41:52:@36924.4]
  assign output_63_38 = io_outValid_38 & _T_75765; // @[Switch.scala 41:38:@36925.4]
  assign _T_75768 = select_39 == 6'h3f; // @[Switch.scala 41:52:@36927.4]
  assign output_63_39 = io_outValid_39 & _T_75768; // @[Switch.scala 41:38:@36928.4]
  assign _T_75771 = select_40 == 6'h3f; // @[Switch.scala 41:52:@36930.4]
  assign output_63_40 = io_outValid_40 & _T_75771; // @[Switch.scala 41:38:@36931.4]
  assign _T_75774 = select_41 == 6'h3f; // @[Switch.scala 41:52:@36933.4]
  assign output_63_41 = io_outValid_41 & _T_75774; // @[Switch.scala 41:38:@36934.4]
  assign _T_75777 = select_42 == 6'h3f; // @[Switch.scala 41:52:@36936.4]
  assign output_63_42 = io_outValid_42 & _T_75777; // @[Switch.scala 41:38:@36937.4]
  assign _T_75780 = select_43 == 6'h3f; // @[Switch.scala 41:52:@36939.4]
  assign output_63_43 = io_outValid_43 & _T_75780; // @[Switch.scala 41:38:@36940.4]
  assign _T_75783 = select_44 == 6'h3f; // @[Switch.scala 41:52:@36942.4]
  assign output_63_44 = io_outValid_44 & _T_75783; // @[Switch.scala 41:38:@36943.4]
  assign _T_75786 = select_45 == 6'h3f; // @[Switch.scala 41:52:@36945.4]
  assign output_63_45 = io_outValid_45 & _T_75786; // @[Switch.scala 41:38:@36946.4]
  assign _T_75789 = select_46 == 6'h3f; // @[Switch.scala 41:52:@36948.4]
  assign output_63_46 = io_outValid_46 & _T_75789; // @[Switch.scala 41:38:@36949.4]
  assign _T_75792 = select_47 == 6'h3f; // @[Switch.scala 41:52:@36951.4]
  assign output_63_47 = io_outValid_47 & _T_75792; // @[Switch.scala 41:38:@36952.4]
  assign _T_75795 = select_48 == 6'h3f; // @[Switch.scala 41:52:@36954.4]
  assign output_63_48 = io_outValid_48 & _T_75795; // @[Switch.scala 41:38:@36955.4]
  assign _T_75798 = select_49 == 6'h3f; // @[Switch.scala 41:52:@36957.4]
  assign output_63_49 = io_outValid_49 & _T_75798; // @[Switch.scala 41:38:@36958.4]
  assign _T_75801 = select_50 == 6'h3f; // @[Switch.scala 41:52:@36960.4]
  assign output_63_50 = io_outValid_50 & _T_75801; // @[Switch.scala 41:38:@36961.4]
  assign _T_75804 = select_51 == 6'h3f; // @[Switch.scala 41:52:@36963.4]
  assign output_63_51 = io_outValid_51 & _T_75804; // @[Switch.scala 41:38:@36964.4]
  assign _T_75807 = select_52 == 6'h3f; // @[Switch.scala 41:52:@36966.4]
  assign output_63_52 = io_outValid_52 & _T_75807; // @[Switch.scala 41:38:@36967.4]
  assign _T_75810 = select_53 == 6'h3f; // @[Switch.scala 41:52:@36969.4]
  assign output_63_53 = io_outValid_53 & _T_75810; // @[Switch.scala 41:38:@36970.4]
  assign _T_75813 = select_54 == 6'h3f; // @[Switch.scala 41:52:@36972.4]
  assign output_63_54 = io_outValid_54 & _T_75813; // @[Switch.scala 41:38:@36973.4]
  assign _T_75816 = select_55 == 6'h3f; // @[Switch.scala 41:52:@36975.4]
  assign output_63_55 = io_outValid_55 & _T_75816; // @[Switch.scala 41:38:@36976.4]
  assign _T_75819 = select_56 == 6'h3f; // @[Switch.scala 41:52:@36978.4]
  assign output_63_56 = io_outValid_56 & _T_75819; // @[Switch.scala 41:38:@36979.4]
  assign _T_75822 = select_57 == 6'h3f; // @[Switch.scala 41:52:@36981.4]
  assign output_63_57 = io_outValid_57 & _T_75822; // @[Switch.scala 41:38:@36982.4]
  assign _T_75825 = select_58 == 6'h3f; // @[Switch.scala 41:52:@36984.4]
  assign output_63_58 = io_outValid_58 & _T_75825; // @[Switch.scala 41:38:@36985.4]
  assign _T_75828 = select_59 == 6'h3f; // @[Switch.scala 41:52:@36987.4]
  assign output_63_59 = io_outValid_59 & _T_75828; // @[Switch.scala 41:38:@36988.4]
  assign _T_75831 = select_60 == 6'h3f; // @[Switch.scala 41:52:@36990.4]
  assign output_63_60 = io_outValid_60 & _T_75831; // @[Switch.scala 41:38:@36991.4]
  assign _T_75834 = select_61 == 6'h3f; // @[Switch.scala 41:52:@36993.4]
  assign output_63_61 = io_outValid_61 & _T_75834; // @[Switch.scala 41:38:@36994.4]
  assign _T_75837 = select_62 == 6'h3f; // @[Switch.scala 41:52:@36996.4]
  assign output_63_62 = io_outValid_62 & _T_75837; // @[Switch.scala 41:38:@36997.4]
  assign _T_75840 = select_63 == 6'h3f; // @[Switch.scala 41:52:@36999.4]
  assign output_63_63 = io_outValid_63 & _T_75840; // @[Switch.scala 41:38:@37000.4]
  assign _T_75848 = {output_63_7,output_63_6,output_63_5,output_63_4,output_63_3,output_63_2,output_63_1,output_63_0}; // @[Switch.scala 43:31:@37008.4]
  assign _T_75856 = {output_63_15,output_63_14,output_63_13,output_63_12,output_63_11,output_63_10,output_63_9,output_63_8,_T_75848}; // @[Switch.scala 43:31:@37016.4]
  assign _T_75863 = {output_63_23,output_63_22,output_63_21,output_63_20,output_63_19,output_63_18,output_63_17,output_63_16}; // @[Switch.scala 43:31:@37023.4]
  assign _T_75872 = {output_63_31,output_63_30,output_63_29,output_63_28,output_63_27,output_63_26,output_63_25,output_63_24,_T_75863,_T_75856}; // @[Switch.scala 43:31:@37032.4]
  assign _T_75879 = {output_63_39,output_63_38,output_63_37,output_63_36,output_63_35,output_63_34,output_63_33,output_63_32}; // @[Switch.scala 43:31:@37039.4]
  assign _T_75887 = {output_63_47,output_63_46,output_63_45,output_63_44,output_63_43,output_63_42,output_63_41,output_63_40,_T_75879}; // @[Switch.scala 43:31:@37047.4]
  assign _T_75894 = {output_63_55,output_63_54,output_63_53,output_63_52,output_63_51,output_63_50,output_63_49,output_63_48}; // @[Switch.scala 43:31:@37054.4]
  assign _T_75903 = {output_63_63,output_63_62,output_63_61,output_63_60,output_63_59,output_63_58,output_63_57,output_63_56,_T_75894,_T_75887}; // @[Switch.scala 43:31:@37063.4]
  assign _T_75904 = {_T_75903,_T_75872}; // @[Switch.scala 43:31:@37064.4]
  assign io_outAck_0 = _T_59713 != 64'h0; // @[Switch.scala 43:18:@20875.4]
  assign io_outAck_1 = _T_59970 != 64'h0; // @[Switch.scala 43:18:@21132.4]
  assign io_outAck_2 = _T_60227 != 64'h0; // @[Switch.scala 43:18:@21389.4]
  assign io_outAck_3 = _T_60484 != 64'h0; // @[Switch.scala 43:18:@21646.4]
  assign io_outAck_4 = _T_60741 != 64'h0; // @[Switch.scala 43:18:@21903.4]
  assign io_outAck_5 = _T_60998 != 64'h0; // @[Switch.scala 43:18:@22160.4]
  assign io_outAck_6 = _T_61255 != 64'h0; // @[Switch.scala 43:18:@22417.4]
  assign io_outAck_7 = _T_61512 != 64'h0; // @[Switch.scala 43:18:@22674.4]
  assign io_outAck_8 = _T_61769 != 64'h0; // @[Switch.scala 43:18:@22931.4]
  assign io_outAck_9 = _T_62026 != 64'h0; // @[Switch.scala 43:18:@23188.4]
  assign io_outAck_10 = _T_62283 != 64'h0; // @[Switch.scala 43:18:@23445.4]
  assign io_outAck_11 = _T_62540 != 64'h0; // @[Switch.scala 43:18:@23702.4]
  assign io_outAck_12 = _T_62797 != 64'h0; // @[Switch.scala 43:18:@23959.4]
  assign io_outAck_13 = _T_63054 != 64'h0; // @[Switch.scala 43:18:@24216.4]
  assign io_outAck_14 = _T_63311 != 64'h0; // @[Switch.scala 43:18:@24473.4]
  assign io_outAck_15 = _T_63568 != 64'h0; // @[Switch.scala 43:18:@24730.4]
  assign io_outAck_16 = _T_63825 != 64'h0; // @[Switch.scala 43:18:@24987.4]
  assign io_outAck_17 = _T_64082 != 64'h0; // @[Switch.scala 43:18:@25244.4]
  assign io_outAck_18 = _T_64339 != 64'h0; // @[Switch.scala 43:18:@25501.4]
  assign io_outAck_19 = _T_64596 != 64'h0; // @[Switch.scala 43:18:@25758.4]
  assign io_outAck_20 = _T_64853 != 64'h0; // @[Switch.scala 43:18:@26015.4]
  assign io_outAck_21 = _T_65110 != 64'h0; // @[Switch.scala 43:18:@26272.4]
  assign io_outAck_22 = _T_65367 != 64'h0; // @[Switch.scala 43:18:@26529.4]
  assign io_outAck_23 = _T_65624 != 64'h0; // @[Switch.scala 43:18:@26786.4]
  assign io_outAck_24 = _T_65881 != 64'h0; // @[Switch.scala 43:18:@27043.4]
  assign io_outAck_25 = _T_66138 != 64'h0; // @[Switch.scala 43:18:@27300.4]
  assign io_outAck_26 = _T_66395 != 64'h0; // @[Switch.scala 43:18:@27557.4]
  assign io_outAck_27 = _T_66652 != 64'h0; // @[Switch.scala 43:18:@27814.4]
  assign io_outAck_28 = _T_66909 != 64'h0; // @[Switch.scala 43:18:@28071.4]
  assign io_outAck_29 = _T_67166 != 64'h0; // @[Switch.scala 43:18:@28328.4]
  assign io_outAck_30 = _T_67423 != 64'h0; // @[Switch.scala 43:18:@28585.4]
  assign io_outAck_31 = _T_67680 != 64'h0; // @[Switch.scala 43:18:@28842.4]
  assign io_outAck_32 = _T_67937 != 64'h0; // @[Switch.scala 43:18:@29099.4]
  assign io_outAck_33 = _T_68194 != 64'h0; // @[Switch.scala 43:18:@29356.4]
  assign io_outAck_34 = _T_68451 != 64'h0; // @[Switch.scala 43:18:@29613.4]
  assign io_outAck_35 = _T_68708 != 64'h0; // @[Switch.scala 43:18:@29870.4]
  assign io_outAck_36 = _T_68965 != 64'h0; // @[Switch.scala 43:18:@30127.4]
  assign io_outAck_37 = _T_69222 != 64'h0; // @[Switch.scala 43:18:@30384.4]
  assign io_outAck_38 = _T_69479 != 64'h0; // @[Switch.scala 43:18:@30641.4]
  assign io_outAck_39 = _T_69736 != 64'h0; // @[Switch.scala 43:18:@30898.4]
  assign io_outAck_40 = _T_69993 != 64'h0; // @[Switch.scala 43:18:@31155.4]
  assign io_outAck_41 = _T_70250 != 64'h0; // @[Switch.scala 43:18:@31412.4]
  assign io_outAck_42 = _T_70507 != 64'h0; // @[Switch.scala 43:18:@31669.4]
  assign io_outAck_43 = _T_70764 != 64'h0; // @[Switch.scala 43:18:@31926.4]
  assign io_outAck_44 = _T_71021 != 64'h0; // @[Switch.scala 43:18:@32183.4]
  assign io_outAck_45 = _T_71278 != 64'h0; // @[Switch.scala 43:18:@32440.4]
  assign io_outAck_46 = _T_71535 != 64'h0; // @[Switch.scala 43:18:@32697.4]
  assign io_outAck_47 = _T_71792 != 64'h0; // @[Switch.scala 43:18:@32954.4]
  assign io_outAck_48 = _T_72049 != 64'h0; // @[Switch.scala 43:18:@33211.4]
  assign io_outAck_49 = _T_72306 != 64'h0; // @[Switch.scala 43:18:@33468.4]
  assign io_outAck_50 = _T_72563 != 64'h0; // @[Switch.scala 43:18:@33725.4]
  assign io_outAck_51 = _T_72820 != 64'h0; // @[Switch.scala 43:18:@33982.4]
  assign io_outAck_52 = _T_73077 != 64'h0; // @[Switch.scala 43:18:@34239.4]
  assign io_outAck_53 = _T_73334 != 64'h0; // @[Switch.scala 43:18:@34496.4]
  assign io_outAck_54 = _T_73591 != 64'h0; // @[Switch.scala 43:18:@34753.4]
  assign io_outAck_55 = _T_73848 != 64'h0; // @[Switch.scala 43:18:@35010.4]
  assign io_outAck_56 = _T_74105 != 64'h0; // @[Switch.scala 43:18:@35267.4]
  assign io_outAck_57 = _T_74362 != 64'h0; // @[Switch.scala 43:18:@35524.4]
  assign io_outAck_58 = _T_74619 != 64'h0; // @[Switch.scala 43:18:@35781.4]
  assign io_outAck_59 = _T_74876 != 64'h0; // @[Switch.scala 43:18:@36038.4]
  assign io_outAck_60 = _T_75133 != 64'h0; // @[Switch.scala 43:18:@36295.4]
  assign io_outAck_61 = _T_75390 != 64'h0; // @[Switch.scala 43:18:@36552.4]
  assign io_outAck_62 = _T_75647 != 64'h0; // @[Switch.scala 43:18:@36809.4]
  assign io_outAck_63 = _T_75904 != 64'h0; // @[Switch.scala 43:18:@37066.4]
  assign io_outData_0 = 6'h3f == select_0 ? io_inData_63 : _GEN_62; // @[Switch.scala 33:19:@266.4]
  assign io_outData_1 = 6'h3f == select_1 ? io_inData_63 : _GEN_126; // @[Switch.scala 33:19:@588.4]
  assign io_outData_2 = 6'h3f == select_2 ? io_inData_63 : _GEN_190; // @[Switch.scala 33:19:@910.4]
  assign io_outData_3 = 6'h3f == select_3 ? io_inData_63 : _GEN_254; // @[Switch.scala 33:19:@1232.4]
  assign io_outData_4 = 6'h3f == select_4 ? io_inData_63 : _GEN_318; // @[Switch.scala 33:19:@1554.4]
  assign io_outData_5 = 6'h3f == select_5 ? io_inData_63 : _GEN_382; // @[Switch.scala 33:19:@1876.4]
  assign io_outData_6 = 6'h3f == select_6 ? io_inData_63 : _GEN_446; // @[Switch.scala 33:19:@2198.4]
  assign io_outData_7 = 6'h3f == select_7 ? io_inData_63 : _GEN_510; // @[Switch.scala 33:19:@2520.4]
  assign io_outData_8 = 6'h3f == select_8 ? io_inData_63 : _GEN_574; // @[Switch.scala 33:19:@2842.4]
  assign io_outData_9 = 6'h3f == select_9 ? io_inData_63 : _GEN_638; // @[Switch.scala 33:19:@3164.4]
  assign io_outData_10 = 6'h3f == select_10 ? io_inData_63 : _GEN_702; // @[Switch.scala 33:19:@3486.4]
  assign io_outData_11 = 6'h3f == select_11 ? io_inData_63 : _GEN_766; // @[Switch.scala 33:19:@3808.4]
  assign io_outData_12 = 6'h3f == select_12 ? io_inData_63 : _GEN_830; // @[Switch.scala 33:19:@4130.4]
  assign io_outData_13 = 6'h3f == select_13 ? io_inData_63 : _GEN_894; // @[Switch.scala 33:19:@4452.4]
  assign io_outData_14 = 6'h3f == select_14 ? io_inData_63 : _GEN_958; // @[Switch.scala 33:19:@4774.4]
  assign io_outData_15 = 6'h3f == select_15 ? io_inData_63 : _GEN_1022; // @[Switch.scala 33:19:@5096.4]
  assign io_outData_16 = 6'h3f == select_16 ? io_inData_63 : _GEN_1086; // @[Switch.scala 33:19:@5418.4]
  assign io_outData_17 = 6'h3f == select_17 ? io_inData_63 : _GEN_1150; // @[Switch.scala 33:19:@5740.4]
  assign io_outData_18 = 6'h3f == select_18 ? io_inData_63 : _GEN_1214; // @[Switch.scala 33:19:@6062.4]
  assign io_outData_19 = 6'h3f == select_19 ? io_inData_63 : _GEN_1278; // @[Switch.scala 33:19:@6384.4]
  assign io_outData_20 = 6'h3f == select_20 ? io_inData_63 : _GEN_1342; // @[Switch.scala 33:19:@6706.4]
  assign io_outData_21 = 6'h3f == select_21 ? io_inData_63 : _GEN_1406; // @[Switch.scala 33:19:@7028.4]
  assign io_outData_22 = 6'h3f == select_22 ? io_inData_63 : _GEN_1470; // @[Switch.scala 33:19:@7350.4]
  assign io_outData_23 = 6'h3f == select_23 ? io_inData_63 : _GEN_1534; // @[Switch.scala 33:19:@7672.4]
  assign io_outData_24 = 6'h3f == select_24 ? io_inData_63 : _GEN_1598; // @[Switch.scala 33:19:@7994.4]
  assign io_outData_25 = 6'h3f == select_25 ? io_inData_63 : _GEN_1662; // @[Switch.scala 33:19:@8316.4]
  assign io_outData_26 = 6'h3f == select_26 ? io_inData_63 : _GEN_1726; // @[Switch.scala 33:19:@8638.4]
  assign io_outData_27 = 6'h3f == select_27 ? io_inData_63 : _GEN_1790; // @[Switch.scala 33:19:@8960.4]
  assign io_outData_28 = 6'h3f == select_28 ? io_inData_63 : _GEN_1854; // @[Switch.scala 33:19:@9282.4]
  assign io_outData_29 = 6'h3f == select_29 ? io_inData_63 : _GEN_1918; // @[Switch.scala 33:19:@9604.4]
  assign io_outData_30 = 6'h3f == select_30 ? io_inData_63 : _GEN_1982; // @[Switch.scala 33:19:@9926.4]
  assign io_outData_31 = 6'h3f == select_31 ? io_inData_63 : _GEN_2046; // @[Switch.scala 33:19:@10248.4]
  assign io_outData_32 = 6'h3f == select_32 ? io_inData_63 : _GEN_2110; // @[Switch.scala 33:19:@10570.4]
  assign io_outData_33 = 6'h3f == select_33 ? io_inData_63 : _GEN_2174; // @[Switch.scala 33:19:@10892.4]
  assign io_outData_34 = 6'h3f == select_34 ? io_inData_63 : _GEN_2238; // @[Switch.scala 33:19:@11214.4]
  assign io_outData_35 = 6'h3f == select_35 ? io_inData_63 : _GEN_2302; // @[Switch.scala 33:19:@11536.4]
  assign io_outData_36 = 6'h3f == select_36 ? io_inData_63 : _GEN_2366; // @[Switch.scala 33:19:@11858.4]
  assign io_outData_37 = 6'h3f == select_37 ? io_inData_63 : _GEN_2430; // @[Switch.scala 33:19:@12180.4]
  assign io_outData_38 = 6'h3f == select_38 ? io_inData_63 : _GEN_2494; // @[Switch.scala 33:19:@12502.4]
  assign io_outData_39 = 6'h3f == select_39 ? io_inData_63 : _GEN_2558; // @[Switch.scala 33:19:@12824.4]
  assign io_outData_40 = 6'h3f == select_40 ? io_inData_63 : _GEN_2622; // @[Switch.scala 33:19:@13146.4]
  assign io_outData_41 = 6'h3f == select_41 ? io_inData_63 : _GEN_2686; // @[Switch.scala 33:19:@13468.4]
  assign io_outData_42 = 6'h3f == select_42 ? io_inData_63 : _GEN_2750; // @[Switch.scala 33:19:@13790.4]
  assign io_outData_43 = 6'h3f == select_43 ? io_inData_63 : _GEN_2814; // @[Switch.scala 33:19:@14112.4]
  assign io_outData_44 = 6'h3f == select_44 ? io_inData_63 : _GEN_2878; // @[Switch.scala 33:19:@14434.4]
  assign io_outData_45 = 6'h3f == select_45 ? io_inData_63 : _GEN_2942; // @[Switch.scala 33:19:@14756.4]
  assign io_outData_46 = 6'h3f == select_46 ? io_inData_63 : _GEN_3006; // @[Switch.scala 33:19:@15078.4]
  assign io_outData_47 = 6'h3f == select_47 ? io_inData_63 : _GEN_3070; // @[Switch.scala 33:19:@15400.4]
  assign io_outData_48 = 6'h3f == select_48 ? io_inData_63 : _GEN_3134; // @[Switch.scala 33:19:@15722.4]
  assign io_outData_49 = 6'h3f == select_49 ? io_inData_63 : _GEN_3198; // @[Switch.scala 33:19:@16044.4]
  assign io_outData_50 = 6'h3f == select_50 ? io_inData_63 : _GEN_3262; // @[Switch.scala 33:19:@16366.4]
  assign io_outData_51 = 6'h3f == select_51 ? io_inData_63 : _GEN_3326; // @[Switch.scala 33:19:@16688.4]
  assign io_outData_52 = 6'h3f == select_52 ? io_inData_63 : _GEN_3390; // @[Switch.scala 33:19:@17010.4]
  assign io_outData_53 = 6'h3f == select_53 ? io_inData_63 : _GEN_3454; // @[Switch.scala 33:19:@17332.4]
  assign io_outData_54 = 6'h3f == select_54 ? io_inData_63 : _GEN_3518; // @[Switch.scala 33:19:@17654.4]
  assign io_outData_55 = 6'h3f == select_55 ? io_inData_63 : _GEN_3582; // @[Switch.scala 33:19:@17976.4]
  assign io_outData_56 = 6'h3f == select_56 ? io_inData_63 : _GEN_3646; // @[Switch.scala 33:19:@18298.4]
  assign io_outData_57 = 6'h3f == select_57 ? io_inData_63 : _GEN_3710; // @[Switch.scala 33:19:@18620.4]
  assign io_outData_58 = 6'h3f == select_58 ? io_inData_63 : _GEN_3774; // @[Switch.scala 33:19:@18942.4]
  assign io_outData_59 = 6'h3f == select_59 ? io_inData_63 : _GEN_3838; // @[Switch.scala 33:19:@19264.4]
  assign io_outData_60 = 6'h3f == select_60 ? io_inData_63 : _GEN_3902; // @[Switch.scala 33:19:@19586.4]
  assign io_outData_61 = 6'h3f == select_61 ? io_inData_63 : _GEN_3966; // @[Switch.scala 33:19:@19908.4]
  assign io_outData_62 = 6'h3f == select_62 ? io_inData_63 : _GEN_4030; // @[Switch.scala 33:19:@20230.4]
  assign io_outData_63 = 6'h3f == select_63 ? io_inData_63 : _GEN_4094; // @[Switch.scala 33:19:@20552.4]
  assign io_outValid_0 = _T_18035 != 64'h0; // @[Switch.scala 34:20:@331.4]
  assign io_outValid_1 = _T_18420 != 64'h0; // @[Switch.scala 34:20:@653.4]
  assign io_outValid_2 = _T_18805 != 64'h0; // @[Switch.scala 34:20:@975.4]
  assign io_outValid_3 = _T_19190 != 64'h0; // @[Switch.scala 34:20:@1297.4]
  assign io_outValid_4 = _T_19575 != 64'h0; // @[Switch.scala 34:20:@1619.4]
  assign io_outValid_5 = _T_19960 != 64'h0; // @[Switch.scala 34:20:@1941.4]
  assign io_outValid_6 = _T_20345 != 64'h0; // @[Switch.scala 34:20:@2263.4]
  assign io_outValid_7 = _T_20730 != 64'h0; // @[Switch.scala 34:20:@2585.4]
  assign io_outValid_8 = _T_21115 != 64'h0; // @[Switch.scala 34:20:@2907.4]
  assign io_outValid_9 = _T_21500 != 64'h0; // @[Switch.scala 34:20:@3229.4]
  assign io_outValid_10 = _T_21885 != 64'h0; // @[Switch.scala 34:20:@3551.4]
  assign io_outValid_11 = _T_22270 != 64'h0; // @[Switch.scala 34:20:@3873.4]
  assign io_outValid_12 = _T_22655 != 64'h0; // @[Switch.scala 34:20:@4195.4]
  assign io_outValid_13 = _T_23040 != 64'h0; // @[Switch.scala 34:20:@4517.4]
  assign io_outValid_14 = _T_23425 != 64'h0; // @[Switch.scala 34:20:@4839.4]
  assign io_outValid_15 = _T_23810 != 64'h0; // @[Switch.scala 34:20:@5161.4]
  assign io_outValid_16 = _T_24195 != 64'h0; // @[Switch.scala 34:20:@5483.4]
  assign io_outValid_17 = _T_24580 != 64'h0; // @[Switch.scala 34:20:@5805.4]
  assign io_outValid_18 = _T_24965 != 64'h0; // @[Switch.scala 34:20:@6127.4]
  assign io_outValid_19 = _T_25350 != 64'h0; // @[Switch.scala 34:20:@6449.4]
  assign io_outValid_20 = _T_25735 != 64'h0; // @[Switch.scala 34:20:@6771.4]
  assign io_outValid_21 = _T_26120 != 64'h0; // @[Switch.scala 34:20:@7093.4]
  assign io_outValid_22 = _T_26505 != 64'h0; // @[Switch.scala 34:20:@7415.4]
  assign io_outValid_23 = _T_26890 != 64'h0; // @[Switch.scala 34:20:@7737.4]
  assign io_outValid_24 = _T_27275 != 64'h0; // @[Switch.scala 34:20:@8059.4]
  assign io_outValid_25 = _T_27660 != 64'h0; // @[Switch.scala 34:20:@8381.4]
  assign io_outValid_26 = _T_28045 != 64'h0; // @[Switch.scala 34:20:@8703.4]
  assign io_outValid_27 = _T_28430 != 64'h0; // @[Switch.scala 34:20:@9025.4]
  assign io_outValid_28 = _T_28815 != 64'h0; // @[Switch.scala 34:20:@9347.4]
  assign io_outValid_29 = _T_29200 != 64'h0; // @[Switch.scala 34:20:@9669.4]
  assign io_outValid_30 = _T_29585 != 64'h0; // @[Switch.scala 34:20:@9991.4]
  assign io_outValid_31 = _T_29970 != 64'h0; // @[Switch.scala 34:20:@10313.4]
  assign io_outValid_32 = _T_30355 != 64'h0; // @[Switch.scala 34:20:@10635.4]
  assign io_outValid_33 = _T_30740 != 64'h0; // @[Switch.scala 34:20:@10957.4]
  assign io_outValid_34 = _T_31125 != 64'h0; // @[Switch.scala 34:20:@11279.4]
  assign io_outValid_35 = _T_31510 != 64'h0; // @[Switch.scala 34:20:@11601.4]
  assign io_outValid_36 = _T_31895 != 64'h0; // @[Switch.scala 34:20:@11923.4]
  assign io_outValid_37 = _T_32280 != 64'h0; // @[Switch.scala 34:20:@12245.4]
  assign io_outValid_38 = _T_32665 != 64'h0; // @[Switch.scala 34:20:@12567.4]
  assign io_outValid_39 = _T_33050 != 64'h0; // @[Switch.scala 34:20:@12889.4]
  assign io_outValid_40 = _T_33435 != 64'h0; // @[Switch.scala 34:20:@13211.4]
  assign io_outValid_41 = _T_33820 != 64'h0; // @[Switch.scala 34:20:@13533.4]
  assign io_outValid_42 = _T_34205 != 64'h0; // @[Switch.scala 34:20:@13855.4]
  assign io_outValid_43 = _T_34590 != 64'h0; // @[Switch.scala 34:20:@14177.4]
  assign io_outValid_44 = _T_34975 != 64'h0; // @[Switch.scala 34:20:@14499.4]
  assign io_outValid_45 = _T_35360 != 64'h0; // @[Switch.scala 34:20:@14821.4]
  assign io_outValid_46 = _T_35745 != 64'h0; // @[Switch.scala 34:20:@15143.4]
  assign io_outValid_47 = _T_36130 != 64'h0; // @[Switch.scala 34:20:@15465.4]
  assign io_outValid_48 = _T_36515 != 64'h0; // @[Switch.scala 34:20:@15787.4]
  assign io_outValid_49 = _T_36900 != 64'h0; // @[Switch.scala 34:20:@16109.4]
  assign io_outValid_50 = _T_37285 != 64'h0; // @[Switch.scala 34:20:@16431.4]
  assign io_outValid_51 = _T_37670 != 64'h0; // @[Switch.scala 34:20:@16753.4]
  assign io_outValid_52 = _T_38055 != 64'h0; // @[Switch.scala 34:20:@17075.4]
  assign io_outValid_53 = _T_38440 != 64'h0; // @[Switch.scala 34:20:@17397.4]
  assign io_outValid_54 = _T_38825 != 64'h0; // @[Switch.scala 34:20:@17719.4]
  assign io_outValid_55 = _T_39210 != 64'h0; // @[Switch.scala 34:20:@18041.4]
  assign io_outValid_56 = _T_39595 != 64'h0; // @[Switch.scala 34:20:@18363.4]
  assign io_outValid_57 = _T_39980 != 64'h0; // @[Switch.scala 34:20:@18685.4]
  assign io_outValid_58 = _T_40365 != 64'h0; // @[Switch.scala 34:20:@19007.4]
  assign io_outValid_59 = _T_40750 != 64'h0; // @[Switch.scala 34:20:@19329.4]
  assign io_outValid_60 = _T_41135 != 64'h0; // @[Switch.scala 34:20:@19651.4]
  assign io_outValid_61 = _T_41520 != 64'h0; // @[Switch.scala 34:20:@19973.4]
  assign io_outValid_62 = _T_41905 != 64'h0; // @[Switch.scala 34:20:@20295.4]
  assign io_outValid_63 = _T_42290 != 64'h0; // @[Switch.scala 34:20:@20617.4]
endmodule
module SwitchWrapper( // @[:@37068.2]
  input         clock, // @[:@37069.4]
  input         reset, // @[:@37070.4]
  input  [5:0]  io_inAddr_0, // @[:@37071.4]
  input  [5:0]  io_inAddr_1, // @[:@37071.4]
  input  [5:0]  io_inAddr_2, // @[:@37071.4]
  input  [5:0]  io_inAddr_3, // @[:@37071.4]
  input  [5:0]  io_inAddr_4, // @[:@37071.4]
  input  [5:0]  io_inAddr_5, // @[:@37071.4]
  input  [5:0]  io_inAddr_6, // @[:@37071.4]
  input  [5:0]  io_inAddr_7, // @[:@37071.4]
  input  [5:0]  io_inAddr_8, // @[:@37071.4]
  input  [5:0]  io_inAddr_9, // @[:@37071.4]
  input  [5:0]  io_inAddr_10, // @[:@37071.4]
  input  [5:0]  io_inAddr_11, // @[:@37071.4]
  input  [5:0]  io_inAddr_12, // @[:@37071.4]
  input  [5:0]  io_inAddr_13, // @[:@37071.4]
  input  [5:0]  io_inAddr_14, // @[:@37071.4]
  input  [5:0]  io_inAddr_15, // @[:@37071.4]
  input  [5:0]  io_inAddr_16, // @[:@37071.4]
  input  [5:0]  io_inAddr_17, // @[:@37071.4]
  input  [5:0]  io_inAddr_18, // @[:@37071.4]
  input  [5:0]  io_inAddr_19, // @[:@37071.4]
  input  [5:0]  io_inAddr_20, // @[:@37071.4]
  input  [5:0]  io_inAddr_21, // @[:@37071.4]
  input  [5:0]  io_inAddr_22, // @[:@37071.4]
  input  [5:0]  io_inAddr_23, // @[:@37071.4]
  input  [5:0]  io_inAddr_24, // @[:@37071.4]
  input  [5:0]  io_inAddr_25, // @[:@37071.4]
  input  [5:0]  io_inAddr_26, // @[:@37071.4]
  input  [5:0]  io_inAddr_27, // @[:@37071.4]
  input  [5:0]  io_inAddr_28, // @[:@37071.4]
  input  [5:0]  io_inAddr_29, // @[:@37071.4]
  input  [5:0]  io_inAddr_30, // @[:@37071.4]
  input  [5:0]  io_inAddr_31, // @[:@37071.4]
  input  [5:0]  io_inAddr_32, // @[:@37071.4]
  input  [5:0]  io_inAddr_33, // @[:@37071.4]
  input  [5:0]  io_inAddr_34, // @[:@37071.4]
  input  [5:0]  io_inAddr_35, // @[:@37071.4]
  input  [5:0]  io_inAddr_36, // @[:@37071.4]
  input  [5:0]  io_inAddr_37, // @[:@37071.4]
  input  [5:0]  io_inAddr_38, // @[:@37071.4]
  input  [5:0]  io_inAddr_39, // @[:@37071.4]
  input  [5:0]  io_inAddr_40, // @[:@37071.4]
  input  [5:0]  io_inAddr_41, // @[:@37071.4]
  input  [5:0]  io_inAddr_42, // @[:@37071.4]
  input  [5:0]  io_inAddr_43, // @[:@37071.4]
  input  [5:0]  io_inAddr_44, // @[:@37071.4]
  input  [5:0]  io_inAddr_45, // @[:@37071.4]
  input  [5:0]  io_inAddr_46, // @[:@37071.4]
  input  [5:0]  io_inAddr_47, // @[:@37071.4]
  input  [5:0]  io_inAddr_48, // @[:@37071.4]
  input  [5:0]  io_inAddr_49, // @[:@37071.4]
  input  [5:0]  io_inAddr_50, // @[:@37071.4]
  input  [5:0]  io_inAddr_51, // @[:@37071.4]
  input  [5:0]  io_inAddr_52, // @[:@37071.4]
  input  [5:0]  io_inAddr_53, // @[:@37071.4]
  input  [5:0]  io_inAddr_54, // @[:@37071.4]
  input  [5:0]  io_inAddr_55, // @[:@37071.4]
  input  [5:0]  io_inAddr_56, // @[:@37071.4]
  input  [5:0]  io_inAddr_57, // @[:@37071.4]
  input  [5:0]  io_inAddr_58, // @[:@37071.4]
  input  [5:0]  io_inAddr_59, // @[:@37071.4]
  input  [5:0]  io_inAddr_60, // @[:@37071.4]
  input  [5:0]  io_inAddr_61, // @[:@37071.4]
  input  [5:0]  io_inAddr_62, // @[:@37071.4]
  input  [5:0]  io_inAddr_63, // @[:@37071.4]
  input  [47:0] io_inData_0, // @[:@37071.4]
  input  [47:0] io_inData_1, // @[:@37071.4]
  input  [47:0] io_inData_2, // @[:@37071.4]
  input  [47:0] io_inData_3, // @[:@37071.4]
  input  [47:0] io_inData_4, // @[:@37071.4]
  input  [47:0] io_inData_5, // @[:@37071.4]
  input  [47:0] io_inData_6, // @[:@37071.4]
  input  [47:0] io_inData_7, // @[:@37071.4]
  input  [47:0] io_inData_8, // @[:@37071.4]
  input  [47:0] io_inData_9, // @[:@37071.4]
  input  [47:0] io_inData_10, // @[:@37071.4]
  input  [47:0] io_inData_11, // @[:@37071.4]
  input  [47:0] io_inData_12, // @[:@37071.4]
  input  [47:0] io_inData_13, // @[:@37071.4]
  input  [47:0] io_inData_14, // @[:@37071.4]
  input  [47:0] io_inData_15, // @[:@37071.4]
  input  [47:0] io_inData_16, // @[:@37071.4]
  input  [47:0] io_inData_17, // @[:@37071.4]
  input  [47:0] io_inData_18, // @[:@37071.4]
  input  [47:0] io_inData_19, // @[:@37071.4]
  input  [47:0] io_inData_20, // @[:@37071.4]
  input  [47:0] io_inData_21, // @[:@37071.4]
  input  [47:0] io_inData_22, // @[:@37071.4]
  input  [47:0] io_inData_23, // @[:@37071.4]
  input  [47:0] io_inData_24, // @[:@37071.4]
  input  [47:0] io_inData_25, // @[:@37071.4]
  input  [47:0] io_inData_26, // @[:@37071.4]
  input  [47:0] io_inData_27, // @[:@37071.4]
  input  [47:0] io_inData_28, // @[:@37071.4]
  input  [47:0] io_inData_29, // @[:@37071.4]
  input  [47:0] io_inData_30, // @[:@37071.4]
  input  [47:0] io_inData_31, // @[:@37071.4]
  input  [47:0] io_inData_32, // @[:@37071.4]
  input  [47:0] io_inData_33, // @[:@37071.4]
  input  [47:0] io_inData_34, // @[:@37071.4]
  input  [47:0] io_inData_35, // @[:@37071.4]
  input  [47:0] io_inData_36, // @[:@37071.4]
  input  [47:0] io_inData_37, // @[:@37071.4]
  input  [47:0] io_inData_38, // @[:@37071.4]
  input  [47:0] io_inData_39, // @[:@37071.4]
  input  [47:0] io_inData_40, // @[:@37071.4]
  input  [47:0] io_inData_41, // @[:@37071.4]
  input  [47:0] io_inData_42, // @[:@37071.4]
  input  [47:0] io_inData_43, // @[:@37071.4]
  input  [47:0] io_inData_44, // @[:@37071.4]
  input  [47:0] io_inData_45, // @[:@37071.4]
  input  [47:0] io_inData_46, // @[:@37071.4]
  input  [47:0] io_inData_47, // @[:@37071.4]
  input  [47:0] io_inData_48, // @[:@37071.4]
  input  [47:0] io_inData_49, // @[:@37071.4]
  input  [47:0] io_inData_50, // @[:@37071.4]
  input  [47:0] io_inData_51, // @[:@37071.4]
  input  [47:0] io_inData_52, // @[:@37071.4]
  input  [47:0] io_inData_53, // @[:@37071.4]
  input  [47:0] io_inData_54, // @[:@37071.4]
  input  [47:0] io_inData_55, // @[:@37071.4]
  input  [47:0] io_inData_56, // @[:@37071.4]
  input  [47:0] io_inData_57, // @[:@37071.4]
  input  [47:0] io_inData_58, // @[:@37071.4]
  input  [47:0] io_inData_59, // @[:@37071.4]
  input  [47:0] io_inData_60, // @[:@37071.4]
  input  [47:0] io_inData_61, // @[:@37071.4]
  input  [47:0] io_inData_62, // @[:@37071.4]
  input  [47:0] io_inData_63, // @[:@37071.4]
  input         io_inValid_0, // @[:@37071.4]
  input         io_inValid_1, // @[:@37071.4]
  input         io_inValid_2, // @[:@37071.4]
  input         io_inValid_3, // @[:@37071.4]
  input         io_inValid_4, // @[:@37071.4]
  input         io_inValid_5, // @[:@37071.4]
  input         io_inValid_6, // @[:@37071.4]
  input         io_inValid_7, // @[:@37071.4]
  input         io_inValid_8, // @[:@37071.4]
  input         io_inValid_9, // @[:@37071.4]
  input         io_inValid_10, // @[:@37071.4]
  input         io_inValid_11, // @[:@37071.4]
  input         io_inValid_12, // @[:@37071.4]
  input         io_inValid_13, // @[:@37071.4]
  input         io_inValid_14, // @[:@37071.4]
  input         io_inValid_15, // @[:@37071.4]
  input         io_inValid_16, // @[:@37071.4]
  input         io_inValid_17, // @[:@37071.4]
  input         io_inValid_18, // @[:@37071.4]
  input         io_inValid_19, // @[:@37071.4]
  input         io_inValid_20, // @[:@37071.4]
  input         io_inValid_21, // @[:@37071.4]
  input         io_inValid_22, // @[:@37071.4]
  input         io_inValid_23, // @[:@37071.4]
  input         io_inValid_24, // @[:@37071.4]
  input         io_inValid_25, // @[:@37071.4]
  input         io_inValid_26, // @[:@37071.4]
  input         io_inValid_27, // @[:@37071.4]
  input         io_inValid_28, // @[:@37071.4]
  input         io_inValid_29, // @[:@37071.4]
  input         io_inValid_30, // @[:@37071.4]
  input         io_inValid_31, // @[:@37071.4]
  input         io_inValid_32, // @[:@37071.4]
  input         io_inValid_33, // @[:@37071.4]
  input         io_inValid_34, // @[:@37071.4]
  input         io_inValid_35, // @[:@37071.4]
  input         io_inValid_36, // @[:@37071.4]
  input         io_inValid_37, // @[:@37071.4]
  input         io_inValid_38, // @[:@37071.4]
  input         io_inValid_39, // @[:@37071.4]
  input         io_inValid_40, // @[:@37071.4]
  input         io_inValid_41, // @[:@37071.4]
  input         io_inValid_42, // @[:@37071.4]
  input         io_inValid_43, // @[:@37071.4]
  input         io_inValid_44, // @[:@37071.4]
  input         io_inValid_45, // @[:@37071.4]
  input         io_inValid_46, // @[:@37071.4]
  input         io_inValid_47, // @[:@37071.4]
  input         io_inValid_48, // @[:@37071.4]
  input         io_inValid_49, // @[:@37071.4]
  input         io_inValid_50, // @[:@37071.4]
  input         io_inValid_51, // @[:@37071.4]
  input         io_inValid_52, // @[:@37071.4]
  input         io_inValid_53, // @[:@37071.4]
  input         io_inValid_54, // @[:@37071.4]
  input         io_inValid_55, // @[:@37071.4]
  input         io_inValid_56, // @[:@37071.4]
  input         io_inValid_57, // @[:@37071.4]
  input         io_inValid_58, // @[:@37071.4]
  input         io_inValid_59, // @[:@37071.4]
  input         io_inValid_60, // @[:@37071.4]
  input         io_inValid_61, // @[:@37071.4]
  input         io_inValid_62, // @[:@37071.4]
  input         io_inValid_63, // @[:@37071.4]
  output        io_outAck_0, // @[:@37071.4]
  output        io_outAck_1, // @[:@37071.4]
  output        io_outAck_2, // @[:@37071.4]
  output        io_outAck_3, // @[:@37071.4]
  output        io_outAck_4, // @[:@37071.4]
  output        io_outAck_5, // @[:@37071.4]
  output        io_outAck_6, // @[:@37071.4]
  output        io_outAck_7, // @[:@37071.4]
  output        io_outAck_8, // @[:@37071.4]
  output        io_outAck_9, // @[:@37071.4]
  output        io_outAck_10, // @[:@37071.4]
  output        io_outAck_11, // @[:@37071.4]
  output        io_outAck_12, // @[:@37071.4]
  output        io_outAck_13, // @[:@37071.4]
  output        io_outAck_14, // @[:@37071.4]
  output        io_outAck_15, // @[:@37071.4]
  output        io_outAck_16, // @[:@37071.4]
  output        io_outAck_17, // @[:@37071.4]
  output        io_outAck_18, // @[:@37071.4]
  output        io_outAck_19, // @[:@37071.4]
  output        io_outAck_20, // @[:@37071.4]
  output        io_outAck_21, // @[:@37071.4]
  output        io_outAck_22, // @[:@37071.4]
  output        io_outAck_23, // @[:@37071.4]
  output        io_outAck_24, // @[:@37071.4]
  output        io_outAck_25, // @[:@37071.4]
  output        io_outAck_26, // @[:@37071.4]
  output        io_outAck_27, // @[:@37071.4]
  output        io_outAck_28, // @[:@37071.4]
  output        io_outAck_29, // @[:@37071.4]
  output        io_outAck_30, // @[:@37071.4]
  output        io_outAck_31, // @[:@37071.4]
  output        io_outAck_32, // @[:@37071.4]
  output        io_outAck_33, // @[:@37071.4]
  output        io_outAck_34, // @[:@37071.4]
  output        io_outAck_35, // @[:@37071.4]
  output        io_outAck_36, // @[:@37071.4]
  output        io_outAck_37, // @[:@37071.4]
  output        io_outAck_38, // @[:@37071.4]
  output        io_outAck_39, // @[:@37071.4]
  output        io_outAck_40, // @[:@37071.4]
  output        io_outAck_41, // @[:@37071.4]
  output        io_outAck_42, // @[:@37071.4]
  output        io_outAck_43, // @[:@37071.4]
  output        io_outAck_44, // @[:@37071.4]
  output        io_outAck_45, // @[:@37071.4]
  output        io_outAck_46, // @[:@37071.4]
  output        io_outAck_47, // @[:@37071.4]
  output        io_outAck_48, // @[:@37071.4]
  output        io_outAck_49, // @[:@37071.4]
  output        io_outAck_50, // @[:@37071.4]
  output        io_outAck_51, // @[:@37071.4]
  output        io_outAck_52, // @[:@37071.4]
  output        io_outAck_53, // @[:@37071.4]
  output        io_outAck_54, // @[:@37071.4]
  output        io_outAck_55, // @[:@37071.4]
  output        io_outAck_56, // @[:@37071.4]
  output        io_outAck_57, // @[:@37071.4]
  output        io_outAck_58, // @[:@37071.4]
  output        io_outAck_59, // @[:@37071.4]
  output        io_outAck_60, // @[:@37071.4]
  output        io_outAck_61, // @[:@37071.4]
  output        io_outAck_62, // @[:@37071.4]
  output        io_outAck_63, // @[:@37071.4]
  output [47:0] io_outData_0, // @[:@37071.4]
  output [47:0] io_outData_1, // @[:@37071.4]
  output [47:0] io_outData_2, // @[:@37071.4]
  output [47:0] io_outData_3, // @[:@37071.4]
  output [47:0] io_outData_4, // @[:@37071.4]
  output [47:0] io_outData_5, // @[:@37071.4]
  output [47:0] io_outData_6, // @[:@37071.4]
  output [47:0] io_outData_7, // @[:@37071.4]
  output [47:0] io_outData_8, // @[:@37071.4]
  output [47:0] io_outData_9, // @[:@37071.4]
  output [47:0] io_outData_10, // @[:@37071.4]
  output [47:0] io_outData_11, // @[:@37071.4]
  output [47:0] io_outData_12, // @[:@37071.4]
  output [47:0] io_outData_13, // @[:@37071.4]
  output [47:0] io_outData_14, // @[:@37071.4]
  output [47:0] io_outData_15, // @[:@37071.4]
  output [47:0] io_outData_16, // @[:@37071.4]
  output [47:0] io_outData_17, // @[:@37071.4]
  output [47:0] io_outData_18, // @[:@37071.4]
  output [47:0] io_outData_19, // @[:@37071.4]
  output [47:0] io_outData_20, // @[:@37071.4]
  output [47:0] io_outData_21, // @[:@37071.4]
  output [47:0] io_outData_22, // @[:@37071.4]
  output [47:0] io_outData_23, // @[:@37071.4]
  output [47:0] io_outData_24, // @[:@37071.4]
  output [47:0] io_outData_25, // @[:@37071.4]
  output [47:0] io_outData_26, // @[:@37071.4]
  output [47:0] io_outData_27, // @[:@37071.4]
  output [47:0] io_outData_28, // @[:@37071.4]
  output [47:0] io_outData_29, // @[:@37071.4]
  output [47:0] io_outData_30, // @[:@37071.4]
  output [47:0] io_outData_31, // @[:@37071.4]
  output [47:0] io_outData_32, // @[:@37071.4]
  output [47:0] io_outData_33, // @[:@37071.4]
  output [47:0] io_outData_34, // @[:@37071.4]
  output [47:0] io_outData_35, // @[:@37071.4]
  output [47:0] io_outData_36, // @[:@37071.4]
  output [47:0] io_outData_37, // @[:@37071.4]
  output [47:0] io_outData_38, // @[:@37071.4]
  output [47:0] io_outData_39, // @[:@37071.4]
  output [47:0] io_outData_40, // @[:@37071.4]
  output [47:0] io_outData_41, // @[:@37071.4]
  output [47:0] io_outData_42, // @[:@37071.4]
  output [47:0] io_outData_43, // @[:@37071.4]
  output [47:0] io_outData_44, // @[:@37071.4]
  output [47:0] io_outData_45, // @[:@37071.4]
  output [47:0] io_outData_46, // @[:@37071.4]
  output [47:0] io_outData_47, // @[:@37071.4]
  output [47:0] io_outData_48, // @[:@37071.4]
  output [47:0] io_outData_49, // @[:@37071.4]
  output [47:0] io_outData_50, // @[:@37071.4]
  output [47:0] io_outData_51, // @[:@37071.4]
  output [47:0] io_outData_52, // @[:@37071.4]
  output [47:0] io_outData_53, // @[:@37071.4]
  output [47:0] io_outData_54, // @[:@37071.4]
  output [47:0] io_outData_55, // @[:@37071.4]
  output [47:0] io_outData_56, // @[:@37071.4]
  output [47:0] io_outData_57, // @[:@37071.4]
  output [47:0] io_outData_58, // @[:@37071.4]
  output [47:0] io_outData_59, // @[:@37071.4]
  output [47:0] io_outData_60, // @[:@37071.4]
  output [47:0] io_outData_61, // @[:@37071.4]
  output [47:0] io_outData_62, // @[:@37071.4]
  output [47:0] io_outData_63, // @[:@37071.4]
  output        io_outValid_0, // @[:@37071.4]
  output        io_outValid_1, // @[:@37071.4]
  output        io_outValid_2, // @[:@37071.4]
  output        io_outValid_3, // @[:@37071.4]
  output        io_outValid_4, // @[:@37071.4]
  output        io_outValid_5, // @[:@37071.4]
  output        io_outValid_6, // @[:@37071.4]
  output        io_outValid_7, // @[:@37071.4]
  output        io_outValid_8, // @[:@37071.4]
  output        io_outValid_9, // @[:@37071.4]
  output        io_outValid_10, // @[:@37071.4]
  output        io_outValid_11, // @[:@37071.4]
  output        io_outValid_12, // @[:@37071.4]
  output        io_outValid_13, // @[:@37071.4]
  output        io_outValid_14, // @[:@37071.4]
  output        io_outValid_15, // @[:@37071.4]
  output        io_outValid_16, // @[:@37071.4]
  output        io_outValid_17, // @[:@37071.4]
  output        io_outValid_18, // @[:@37071.4]
  output        io_outValid_19, // @[:@37071.4]
  output        io_outValid_20, // @[:@37071.4]
  output        io_outValid_21, // @[:@37071.4]
  output        io_outValid_22, // @[:@37071.4]
  output        io_outValid_23, // @[:@37071.4]
  output        io_outValid_24, // @[:@37071.4]
  output        io_outValid_25, // @[:@37071.4]
  output        io_outValid_26, // @[:@37071.4]
  output        io_outValid_27, // @[:@37071.4]
  output        io_outValid_28, // @[:@37071.4]
  output        io_outValid_29, // @[:@37071.4]
  output        io_outValid_30, // @[:@37071.4]
  output        io_outValid_31, // @[:@37071.4]
  output        io_outValid_32, // @[:@37071.4]
  output        io_outValid_33, // @[:@37071.4]
  output        io_outValid_34, // @[:@37071.4]
  output        io_outValid_35, // @[:@37071.4]
  output        io_outValid_36, // @[:@37071.4]
  output        io_outValid_37, // @[:@37071.4]
  output        io_outValid_38, // @[:@37071.4]
  output        io_outValid_39, // @[:@37071.4]
  output        io_outValid_40, // @[:@37071.4]
  output        io_outValid_41, // @[:@37071.4]
  output        io_outValid_42, // @[:@37071.4]
  output        io_outValid_43, // @[:@37071.4]
  output        io_outValid_44, // @[:@37071.4]
  output        io_outValid_45, // @[:@37071.4]
  output        io_outValid_46, // @[:@37071.4]
  output        io_outValid_47, // @[:@37071.4]
  output        io_outValid_48, // @[:@37071.4]
  output        io_outValid_49, // @[:@37071.4]
  output        io_outValid_50, // @[:@37071.4]
  output        io_outValid_51, // @[:@37071.4]
  output        io_outValid_52, // @[:@37071.4]
  output        io_outValid_53, // @[:@37071.4]
  output        io_outValid_54, // @[:@37071.4]
  output        io_outValid_55, // @[:@37071.4]
  output        io_outValid_56, // @[:@37071.4]
  output        io_outValid_57, // @[:@37071.4]
  output        io_outValid_58, // @[:@37071.4]
  output        io_outValid_59, // @[:@37071.4]
  output        io_outValid_60, // @[:@37071.4]
  output        io_outValid_61, // @[:@37071.4]
  output        io_outValid_62, // @[:@37071.4]
  output        io_outValid_63 // @[:@37071.4]
);
  wire [5:0] switch_io_inAddr_0; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_1; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_2; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_3; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_4; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_5; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_6; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_7; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_8; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_9; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_10; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_11; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_12; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_13; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_14; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_15; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_16; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_17; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_18; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_19; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_20; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_21; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_22; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_23; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_24; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_25; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_26; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_27; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_28; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_29; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_30; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_31; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_32; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_33; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_34; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_35; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_36; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_37; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_38; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_39; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_40; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_41; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_42; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_43; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_44; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_45; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_46; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_47; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_48; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_49; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_50; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_51; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_52; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_53; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_54; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_55; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_56; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_57; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_58; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_59; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_60; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_61; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_62; // @[Switch.scala 50:22:@37073.4]
  wire [5:0] switch_io_inAddr_63; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_0; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_1; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_2; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_3; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_4; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_5; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_6; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_7; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_8; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_9; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_10; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_11; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_12; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_13; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_14; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_15; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_16; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_17; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_18; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_19; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_20; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_21; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_22; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_23; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_24; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_25; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_26; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_27; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_28; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_29; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_30; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_31; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_32; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_33; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_34; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_35; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_36; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_37; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_38; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_39; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_40; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_41; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_42; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_43; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_44; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_45; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_46; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_47; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_48; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_49; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_50; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_51; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_52; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_53; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_54; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_55; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_56; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_57; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_58; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_59; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_60; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_61; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_62; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_inData_63; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_0; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_1; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_2; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_3; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_4; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_5; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_6; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_7; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_8; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_9; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_10; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_11; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_12; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_13; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_14; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_15; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_16; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_17; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_18; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_19; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_20; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_21; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_22; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_23; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_24; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_25; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_26; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_27; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_28; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_29; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_30; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_31; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_32; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_33; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_34; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_35; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_36; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_37; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_38; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_39; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_40; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_41; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_42; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_43; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_44; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_45; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_46; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_47; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_48; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_49; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_50; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_51; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_52; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_53; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_54; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_55; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_56; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_57; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_58; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_59; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_60; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_61; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_62; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_inValid_63; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_0; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_1; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_2; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_3; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_4; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_5; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_6; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_7; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_8; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_9; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_10; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_11; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_12; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_13; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_14; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_15; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_16; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_17; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_18; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_19; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_20; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_21; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_22; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_23; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_24; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_25; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_26; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_27; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_28; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_29; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_30; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_31; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_32; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_33; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_34; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_35; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_36; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_37; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_38; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_39; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_40; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_41; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_42; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_43; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_44; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_45; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_46; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_47; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_48; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_49; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_50; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_51; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_52; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_53; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_54; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_55; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_56; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_57; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_58; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_59; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_60; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_61; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_62; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outAck_63; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_0; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_1; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_2; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_3; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_4; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_5; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_6; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_7; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_8; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_9; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_10; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_11; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_12; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_13; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_14; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_15; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_16; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_17; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_18; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_19; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_20; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_21; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_22; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_23; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_24; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_25; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_26; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_27; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_28; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_29; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_30; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_31; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_32; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_33; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_34; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_35; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_36; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_37; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_38; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_39; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_40; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_41; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_42; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_43; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_44; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_45; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_46; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_47; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_48; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_49; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_50; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_51; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_52; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_53; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_54; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_55; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_56; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_57; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_58; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_59; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_60; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_61; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_62; // @[Switch.scala 50:22:@37073.4]
  wire [47:0] switch_io_outData_63; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_0; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_1; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_2; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_3; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_4; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_5; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_6; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_7; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_8; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_9; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_10; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_11; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_12; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_13; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_14; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_15; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_16; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_17; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_18; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_19; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_20; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_21; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_22; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_23; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_24; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_25; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_26; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_27; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_28; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_29; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_30; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_31; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_32; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_33; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_34; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_35; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_36; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_37; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_38; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_39; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_40; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_41; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_42; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_43; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_44; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_45; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_46; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_47; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_48; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_49; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_50; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_51; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_52; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_53; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_54; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_55; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_56; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_57; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_58; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_59; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_60; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_61; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_62; // @[Switch.scala 50:22:@37073.4]
  wire  switch_io_outValid_63; // @[Switch.scala 50:22:@37073.4]
  reg [5:0] _T_550_0; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_0;
  reg [5:0] _T_550_1; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_1;
  reg [5:0] _T_550_2; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_2;
  reg [5:0] _T_550_3; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_3;
  reg [5:0] _T_550_4; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_4;
  reg [5:0] _T_550_5; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_5;
  reg [5:0] _T_550_6; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_6;
  reg [5:0] _T_550_7; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_7;
  reg [5:0] _T_550_8; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_8;
  reg [5:0] _T_550_9; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_9;
  reg [5:0] _T_550_10; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_10;
  reg [5:0] _T_550_11; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_11;
  reg [5:0] _T_550_12; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_12;
  reg [5:0] _T_550_13; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_13;
  reg [5:0] _T_550_14; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_14;
  reg [5:0] _T_550_15; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_15;
  reg [5:0] _T_550_16; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_16;
  reg [5:0] _T_550_17; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_17;
  reg [5:0] _T_550_18; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_18;
  reg [5:0] _T_550_19; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_19;
  reg [5:0] _T_550_20; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_20;
  reg [5:0] _T_550_21; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_21;
  reg [5:0] _T_550_22; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_22;
  reg [5:0] _T_550_23; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_23;
  reg [5:0] _T_550_24; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_24;
  reg [5:0] _T_550_25; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_25;
  reg [5:0] _T_550_26; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_26;
  reg [5:0] _T_550_27; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_27;
  reg [5:0] _T_550_28; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_28;
  reg [5:0] _T_550_29; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_29;
  reg [5:0] _T_550_30; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_30;
  reg [5:0] _T_550_31; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_31;
  reg [5:0] _T_550_32; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_32;
  reg [5:0] _T_550_33; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_33;
  reg [5:0] _T_550_34; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_34;
  reg [5:0] _T_550_35; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_35;
  reg [5:0] _T_550_36; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_36;
  reg [5:0] _T_550_37; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_37;
  reg [5:0] _T_550_38; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_38;
  reg [5:0] _T_550_39; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_39;
  reg [5:0] _T_550_40; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_40;
  reg [5:0] _T_550_41; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_41;
  reg [5:0] _T_550_42; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_42;
  reg [5:0] _T_550_43; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_43;
  reg [5:0] _T_550_44; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_44;
  reg [5:0] _T_550_45; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_45;
  reg [5:0] _T_550_46; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_46;
  reg [5:0] _T_550_47; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_47;
  reg [5:0] _T_550_48; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_48;
  reg [5:0] _T_550_49; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_49;
  reg [5:0] _T_550_50; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_50;
  reg [5:0] _T_550_51; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_51;
  reg [5:0] _T_550_52; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_52;
  reg [5:0] _T_550_53; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_53;
  reg [5:0] _T_550_54; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_54;
  reg [5:0] _T_550_55; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_55;
  reg [5:0] _T_550_56; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_56;
  reg [5:0] _T_550_57; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_57;
  reg [5:0] _T_550_58; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_58;
  reg [5:0] _T_550_59; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_59;
  reg [5:0] _T_550_60; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_60;
  reg [5:0] _T_550_61; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_61;
  reg [5:0] _T_550_62; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_62;
  reg [5:0] _T_550_63; // @[Switch.scala 51:30:@37076.4]
  reg [31:0] _RAND_63;
  reg [47:0] _T_879_0; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_64;
  reg [47:0] _T_879_1; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_65;
  reg [47:0] _T_879_2; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_66;
  reg [47:0] _T_879_3; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_67;
  reg [47:0] _T_879_4; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_68;
  reg [47:0] _T_879_5; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_69;
  reg [47:0] _T_879_6; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_70;
  reg [47:0] _T_879_7; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_71;
  reg [47:0] _T_879_8; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_72;
  reg [47:0] _T_879_9; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_73;
  reg [47:0] _T_879_10; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_74;
  reg [47:0] _T_879_11; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_75;
  reg [47:0] _T_879_12; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_76;
  reg [47:0] _T_879_13; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_77;
  reg [47:0] _T_879_14; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_78;
  reg [47:0] _T_879_15; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_79;
  reg [47:0] _T_879_16; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_80;
  reg [47:0] _T_879_17; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_81;
  reg [47:0] _T_879_18; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_82;
  reg [47:0] _T_879_19; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_83;
  reg [47:0] _T_879_20; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_84;
  reg [47:0] _T_879_21; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_85;
  reg [47:0] _T_879_22; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_86;
  reg [47:0] _T_879_23; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_87;
  reg [47:0] _T_879_24; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_88;
  reg [47:0] _T_879_25; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_89;
  reg [47:0] _T_879_26; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_90;
  reg [47:0] _T_879_27; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_91;
  reg [47:0] _T_879_28; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_92;
  reg [47:0] _T_879_29; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_93;
  reg [47:0] _T_879_30; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_94;
  reg [47:0] _T_879_31; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_95;
  reg [47:0] _T_879_32; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_96;
  reg [47:0] _T_879_33; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_97;
  reg [47:0] _T_879_34; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_98;
  reg [47:0] _T_879_35; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_99;
  reg [47:0] _T_879_36; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_100;
  reg [47:0] _T_879_37; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_101;
  reg [47:0] _T_879_38; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_102;
  reg [47:0] _T_879_39; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_103;
  reg [47:0] _T_879_40; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_104;
  reg [47:0] _T_879_41; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_105;
  reg [47:0] _T_879_42; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_106;
  reg [47:0] _T_879_43; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_107;
  reg [47:0] _T_879_44; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_108;
  reg [47:0] _T_879_45; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_109;
  reg [47:0] _T_879_46; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_110;
  reg [47:0] _T_879_47; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_111;
  reg [47:0] _T_879_48; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_112;
  reg [47:0] _T_879_49; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_113;
  reg [47:0] _T_879_50; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_114;
  reg [47:0] _T_879_51; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_115;
  reg [47:0] _T_879_52; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_116;
  reg [47:0] _T_879_53; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_117;
  reg [47:0] _T_879_54; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_118;
  reg [47:0] _T_879_55; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_119;
  reg [47:0] _T_879_56; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_120;
  reg [47:0] _T_879_57; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_121;
  reg [47:0] _T_879_58; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_122;
  reg [47:0] _T_879_59; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_123;
  reg [47:0] _T_879_60; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_124;
  reg [47:0] _T_879_61; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_125;
  reg [47:0] _T_879_62; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_126;
  reg [47:0] _T_879_63; // @[Switch.scala 52:30:@37205.4]
  reg [63:0] _RAND_127;
  reg  _T_1208_0; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_128;
  reg  _T_1208_1; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_129;
  reg  _T_1208_2; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_130;
  reg  _T_1208_3; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_131;
  reg  _T_1208_4; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_132;
  reg  _T_1208_5; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_133;
  reg  _T_1208_6; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_134;
  reg  _T_1208_7; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_135;
  reg  _T_1208_8; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_136;
  reg  _T_1208_9; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_137;
  reg  _T_1208_10; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_138;
  reg  _T_1208_11; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_139;
  reg  _T_1208_12; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_140;
  reg  _T_1208_13; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_141;
  reg  _T_1208_14; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_142;
  reg  _T_1208_15; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_143;
  reg  _T_1208_16; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_144;
  reg  _T_1208_17; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_145;
  reg  _T_1208_18; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_146;
  reg  _T_1208_19; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_147;
  reg  _T_1208_20; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_148;
  reg  _T_1208_21; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_149;
  reg  _T_1208_22; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_150;
  reg  _T_1208_23; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_151;
  reg  _T_1208_24; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_152;
  reg  _T_1208_25; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_153;
  reg  _T_1208_26; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_154;
  reg  _T_1208_27; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_155;
  reg  _T_1208_28; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_156;
  reg  _T_1208_29; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_157;
  reg  _T_1208_30; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_158;
  reg  _T_1208_31; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_159;
  reg  _T_1208_32; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_160;
  reg  _T_1208_33; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_161;
  reg  _T_1208_34; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_162;
  reg  _T_1208_35; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_163;
  reg  _T_1208_36; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_164;
  reg  _T_1208_37; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_165;
  reg  _T_1208_38; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_166;
  reg  _T_1208_39; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_167;
  reg  _T_1208_40; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_168;
  reg  _T_1208_41; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_169;
  reg  _T_1208_42; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_170;
  reg  _T_1208_43; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_171;
  reg  _T_1208_44; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_172;
  reg  _T_1208_45; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_173;
  reg  _T_1208_46; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_174;
  reg  _T_1208_47; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_175;
  reg  _T_1208_48; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_176;
  reg  _T_1208_49; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_177;
  reg  _T_1208_50; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_178;
  reg  _T_1208_51; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_179;
  reg  _T_1208_52; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_180;
  reg  _T_1208_53; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_181;
  reg  _T_1208_54; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_182;
  reg  _T_1208_55; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_183;
  reg  _T_1208_56; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_184;
  reg  _T_1208_57; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_185;
  reg  _T_1208_58; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_186;
  reg  _T_1208_59; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_187;
  reg  _T_1208_60; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_188;
  reg  _T_1208_61; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_189;
  reg  _T_1208_62; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_190;
  reg  _T_1208_63; // @[Switch.scala 53:31:@37334.4]
  reg [31:0] _RAND_191;
  reg  _T_1537_0; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_192;
  reg  _T_1537_1; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_193;
  reg  _T_1537_2; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_194;
  reg  _T_1537_3; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_195;
  reg  _T_1537_4; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_196;
  reg  _T_1537_5; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_197;
  reg  _T_1537_6; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_198;
  reg  _T_1537_7; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_199;
  reg  _T_1537_8; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_200;
  reg  _T_1537_9; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_201;
  reg  _T_1537_10; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_202;
  reg  _T_1537_11; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_203;
  reg  _T_1537_12; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_204;
  reg  _T_1537_13; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_205;
  reg  _T_1537_14; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_206;
  reg  _T_1537_15; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_207;
  reg  _T_1537_16; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_208;
  reg  _T_1537_17; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_209;
  reg  _T_1537_18; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_210;
  reg  _T_1537_19; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_211;
  reg  _T_1537_20; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_212;
  reg  _T_1537_21; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_213;
  reg  _T_1537_22; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_214;
  reg  _T_1537_23; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_215;
  reg  _T_1537_24; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_216;
  reg  _T_1537_25; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_217;
  reg  _T_1537_26; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_218;
  reg  _T_1537_27; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_219;
  reg  _T_1537_28; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_220;
  reg  _T_1537_29; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_221;
  reg  _T_1537_30; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_222;
  reg  _T_1537_31; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_223;
  reg  _T_1537_32; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_224;
  reg  _T_1537_33; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_225;
  reg  _T_1537_34; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_226;
  reg  _T_1537_35; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_227;
  reg  _T_1537_36; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_228;
  reg  _T_1537_37; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_229;
  reg  _T_1537_38; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_230;
  reg  _T_1537_39; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_231;
  reg  _T_1537_40; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_232;
  reg  _T_1537_41; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_233;
  reg  _T_1537_42; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_234;
  reg  _T_1537_43; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_235;
  reg  _T_1537_44; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_236;
  reg  _T_1537_45; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_237;
  reg  _T_1537_46; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_238;
  reg  _T_1537_47; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_239;
  reg  _T_1537_48; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_240;
  reg  _T_1537_49; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_241;
  reg  _T_1537_50; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_242;
  reg  _T_1537_51; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_243;
  reg  _T_1537_52; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_244;
  reg  _T_1537_53; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_245;
  reg  _T_1537_54; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_246;
  reg  _T_1537_55; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_247;
  reg  _T_1537_56; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_248;
  reg  _T_1537_57; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_249;
  reg  _T_1537_58; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_250;
  reg  _T_1537_59; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_251;
  reg  _T_1537_60; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_252;
  reg  _T_1537_61; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_253;
  reg  _T_1537_62; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_254;
  reg  _T_1537_63; // @[Switch.scala 54:23:@37463.4]
  reg [31:0] _RAND_255;
  reg [47:0] _T_1866_0; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_256;
  reg [47:0] _T_1866_1; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_257;
  reg [47:0] _T_1866_2; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_258;
  reg [47:0] _T_1866_3; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_259;
  reg [47:0] _T_1866_4; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_260;
  reg [47:0] _T_1866_5; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_261;
  reg [47:0] _T_1866_6; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_262;
  reg [47:0] _T_1866_7; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_263;
  reg [47:0] _T_1866_8; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_264;
  reg [47:0] _T_1866_9; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_265;
  reg [47:0] _T_1866_10; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_266;
  reg [47:0] _T_1866_11; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_267;
  reg [47:0] _T_1866_12; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_268;
  reg [47:0] _T_1866_13; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_269;
  reg [47:0] _T_1866_14; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_270;
  reg [47:0] _T_1866_15; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_271;
  reg [47:0] _T_1866_16; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_272;
  reg [47:0] _T_1866_17; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_273;
  reg [47:0] _T_1866_18; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_274;
  reg [47:0] _T_1866_19; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_275;
  reg [47:0] _T_1866_20; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_276;
  reg [47:0] _T_1866_21; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_277;
  reg [47:0] _T_1866_22; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_278;
  reg [47:0] _T_1866_23; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_279;
  reg [47:0] _T_1866_24; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_280;
  reg [47:0] _T_1866_25; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_281;
  reg [47:0] _T_1866_26; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_282;
  reg [47:0] _T_1866_27; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_283;
  reg [47:0] _T_1866_28; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_284;
  reg [47:0] _T_1866_29; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_285;
  reg [47:0] _T_1866_30; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_286;
  reg [47:0] _T_1866_31; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_287;
  reg [47:0] _T_1866_32; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_288;
  reg [47:0] _T_1866_33; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_289;
  reg [47:0] _T_1866_34; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_290;
  reg [47:0] _T_1866_35; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_291;
  reg [47:0] _T_1866_36; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_292;
  reg [47:0] _T_1866_37; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_293;
  reg [47:0] _T_1866_38; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_294;
  reg [47:0] _T_1866_39; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_295;
  reg [47:0] _T_1866_40; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_296;
  reg [47:0] _T_1866_41; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_297;
  reg [47:0] _T_1866_42; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_298;
  reg [47:0] _T_1866_43; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_299;
  reg [47:0] _T_1866_44; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_300;
  reg [47:0] _T_1866_45; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_301;
  reg [47:0] _T_1866_46; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_302;
  reg [47:0] _T_1866_47; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_303;
  reg [47:0] _T_1866_48; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_304;
  reg [47:0] _T_1866_49; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_305;
  reg [47:0] _T_1866_50; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_306;
  reg [47:0] _T_1866_51; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_307;
  reg [47:0] _T_1866_52; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_308;
  reg [47:0] _T_1866_53; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_309;
  reg [47:0] _T_1866_54; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_310;
  reg [47:0] _T_1866_55; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_311;
  reg [47:0] _T_1866_56; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_312;
  reg [47:0] _T_1866_57; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_313;
  reg [47:0] _T_1866_58; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_314;
  reg [47:0] _T_1866_59; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_315;
  reg [47:0] _T_1866_60; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_316;
  reg [47:0] _T_1866_61; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_317;
  reg [47:0] _T_1866_62; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_318;
  reg [47:0] _T_1866_63; // @[Switch.scala 55:24:@37592.4]
  reg [63:0] _RAND_319;
  reg  _T_2195_0; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_320;
  reg  _T_2195_1; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_321;
  reg  _T_2195_2; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_322;
  reg  _T_2195_3; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_323;
  reg  _T_2195_4; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_324;
  reg  _T_2195_5; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_325;
  reg  _T_2195_6; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_326;
  reg  _T_2195_7; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_327;
  reg  _T_2195_8; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_328;
  reg  _T_2195_9; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_329;
  reg  _T_2195_10; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_330;
  reg  _T_2195_11; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_331;
  reg  _T_2195_12; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_332;
  reg  _T_2195_13; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_333;
  reg  _T_2195_14; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_334;
  reg  _T_2195_15; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_335;
  reg  _T_2195_16; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_336;
  reg  _T_2195_17; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_337;
  reg  _T_2195_18; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_338;
  reg  _T_2195_19; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_339;
  reg  _T_2195_20; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_340;
  reg  _T_2195_21; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_341;
  reg  _T_2195_22; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_342;
  reg  _T_2195_23; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_343;
  reg  _T_2195_24; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_344;
  reg  _T_2195_25; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_345;
  reg  _T_2195_26; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_346;
  reg  _T_2195_27; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_347;
  reg  _T_2195_28; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_348;
  reg  _T_2195_29; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_349;
  reg  _T_2195_30; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_350;
  reg  _T_2195_31; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_351;
  reg  _T_2195_32; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_352;
  reg  _T_2195_33; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_353;
  reg  _T_2195_34; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_354;
  reg  _T_2195_35; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_355;
  reg  _T_2195_36; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_356;
  reg  _T_2195_37; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_357;
  reg  _T_2195_38; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_358;
  reg  _T_2195_39; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_359;
  reg  _T_2195_40; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_360;
  reg  _T_2195_41; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_361;
  reg  _T_2195_42; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_362;
  reg  _T_2195_43; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_363;
  reg  _T_2195_44; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_364;
  reg  _T_2195_45; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_365;
  reg  _T_2195_46; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_366;
  reg  _T_2195_47; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_367;
  reg  _T_2195_48; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_368;
  reg  _T_2195_49; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_369;
  reg  _T_2195_50; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_370;
  reg  _T_2195_51; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_371;
  reg  _T_2195_52; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_372;
  reg  _T_2195_53; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_373;
  reg  _T_2195_54; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_374;
  reg  _T_2195_55; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_375;
  reg  _T_2195_56; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_376;
  reg  _T_2195_57; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_377;
  reg  _T_2195_58; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_378;
  reg  _T_2195_59; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_379;
  reg  _T_2195_60; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_380;
  reg  _T_2195_61; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_381;
  reg  _T_2195_62; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_382;
  reg  _T_2195_63; // @[Switch.scala 56:25:@37721.4]
  reg [31:0] _RAND_383;
  Switch switch ( // @[Switch.scala 50:22:@37073.4]
    .io_inAddr_0(switch_io_inAddr_0),
    .io_inAddr_1(switch_io_inAddr_1),
    .io_inAddr_2(switch_io_inAddr_2),
    .io_inAddr_3(switch_io_inAddr_3),
    .io_inAddr_4(switch_io_inAddr_4),
    .io_inAddr_5(switch_io_inAddr_5),
    .io_inAddr_6(switch_io_inAddr_6),
    .io_inAddr_7(switch_io_inAddr_7),
    .io_inAddr_8(switch_io_inAddr_8),
    .io_inAddr_9(switch_io_inAddr_9),
    .io_inAddr_10(switch_io_inAddr_10),
    .io_inAddr_11(switch_io_inAddr_11),
    .io_inAddr_12(switch_io_inAddr_12),
    .io_inAddr_13(switch_io_inAddr_13),
    .io_inAddr_14(switch_io_inAddr_14),
    .io_inAddr_15(switch_io_inAddr_15),
    .io_inAddr_16(switch_io_inAddr_16),
    .io_inAddr_17(switch_io_inAddr_17),
    .io_inAddr_18(switch_io_inAddr_18),
    .io_inAddr_19(switch_io_inAddr_19),
    .io_inAddr_20(switch_io_inAddr_20),
    .io_inAddr_21(switch_io_inAddr_21),
    .io_inAddr_22(switch_io_inAddr_22),
    .io_inAddr_23(switch_io_inAddr_23),
    .io_inAddr_24(switch_io_inAddr_24),
    .io_inAddr_25(switch_io_inAddr_25),
    .io_inAddr_26(switch_io_inAddr_26),
    .io_inAddr_27(switch_io_inAddr_27),
    .io_inAddr_28(switch_io_inAddr_28),
    .io_inAddr_29(switch_io_inAddr_29),
    .io_inAddr_30(switch_io_inAddr_30),
    .io_inAddr_31(switch_io_inAddr_31),
    .io_inAddr_32(switch_io_inAddr_32),
    .io_inAddr_33(switch_io_inAddr_33),
    .io_inAddr_34(switch_io_inAddr_34),
    .io_inAddr_35(switch_io_inAddr_35),
    .io_inAddr_36(switch_io_inAddr_36),
    .io_inAddr_37(switch_io_inAddr_37),
    .io_inAddr_38(switch_io_inAddr_38),
    .io_inAddr_39(switch_io_inAddr_39),
    .io_inAddr_40(switch_io_inAddr_40),
    .io_inAddr_41(switch_io_inAddr_41),
    .io_inAddr_42(switch_io_inAddr_42),
    .io_inAddr_43(switch_io_inAddr_43),
    .io_inAddr_44(switch_io_inAddr_44),
    .io_inAddr_45(switch_io_inAddr_45),
    .io_inAddr_46(switch_io_inAddr_46),
    .io_inAddr_47(switch_io_inAddr_47),
    .io_inAddr_48(switch_io_inAddr_48),
    .io_inAddr_49(switch_io_inAddr_49),
    .io_inAddr_50(switch_io_inAddr_50),
    .io_inAddr_51(switch_io_inAddr_51),
    .io_inAddr_52(switch_io_inAddr_52),
    .io_inAddr_53(switch_io_inAddr_53),
    .io_inAddr_54(switch_io_inAddr_54),
    .io_inAddr_55(switch_io_inAddr_55),
    .io_inAddr_56(switch_io_inAddr_56),
    .io_inAddr_57(switch_io_inAddr_57),
    .io_inAddr_58(switch_io_inAddr_58),
    .io_inAddr_59(switch_io_inAddr_59),
    .io_inAddr_60(switch_io_inAddr_60),
    .io_inAddr_61(switch_io_inAddr_61),
    .io_inAddr_62(switch_io_inAddr_62),
    .io_inAddr_63(switch_io_inAddr_63),
    .io_inData_0(switch_io_inData_0),
    .io_inData_1(switch_io_inData_1),
    .io_inData_2(switch_io_inData_2),
    .io_inData_3(switch_io_inData_3),
    .io_inData_4(switch_io_inData_4),
    .io_inData_5(switch_io_inData_5),
    .io_inData_6(switch_io_inData_6),
    .io_inData_7(switch_io_inData_7),
    .io_inData_8(switch_io_inData_8),
    .io_inData_9(switch_io_inData_9),
    .io_inData_10(switch_io_inData_10),
    .io_inData_11(switch_io_inData_11),
    .io_inData_12(switch_io_inData_12),
    .io_inData_13(switch_io_inData_13),
    .io_inData_14(switch_io_inData_14),
    .io_inData_15(switch_io_inData_15),
    .io_inData_16(switch_io_inData_16),
    .io_inData_17(switch_io_inData_17),
    .io_inData_18(switch_io_inData_18),
    .io_inData_19(switch_io_inData_19),
    .io_inData_20(switch_io_inData_20),
    .io_inData_21(switch_io_inData_21),
    .io_inData_22(switch_io_inData_22),
    .io_inData_23(switch_io_inData_23),
    .io_inData_24(switch_io_inData_24),
    .io_inData_25(switch_io_inData_25),
    .io_inData_26(switch_io_inData_26),
    .io_inData_27(switch_io_inData_27),
    .io_inData_28(switch_io_inData_28),
    .io_inData_29(switch_io_inData_29),
    .io_inData_30(switch_io_inData_30),
    .io_inData_31(switch_io_inData_31),
    .io_inData_32(switch_io_inData_32),
    .io_inData_33(switch_io_inData_33),
    .io_inData_34(switch_io_inData_34),
    .io_inData_35(switch_io_inData_35),
    .io_inData_36(switch_io_inData_36),
    .io_inData_37(switch_io_inData_37),
    .io_inData_38(switch_io_inData_38),
    .io_inData_39(switch_io_inData_39),
    .io_inData_40(switch_io_inData_40),
    .io_inData_41(switch_io_inData_41),
    .io_inData_42(switch_io_inData_42),
    .io_inData_43(switch_io_inData_43),
    .io_inData_44(switch_io_inData_44),
    .io_inData_45(switch_io_inData_45),
    .io_inData_46(switch_io_inData_46),
    .io_inData_47(switch_io_inData_47),
    .io_inData_48(switch_io_inData_48),
    .io_inData_49(switch_io_inData_49),
    .io_inData_50(switch_io_inData_50),
    .io_inData_51(switch_io_inData_51),
    .io_inData_52(switch_io_inData_52),
    .io_inData_53(switch_io_inData_53),
    .io_inData_54(switch_io_inData_54),
    .io_inData_55(switch_io_inData_55),
    .io_inData_56(switch_io_inData_56),
    .io_inData_57(switch_io_inData_57),
    .io_inData_58(switch_io_inData_58),
    .io_inData_59(switch_io_inData_59),
    .io_inData_60(switch_io_inData_60),
    .io_inData_61(switch_io_inData_61),
    .io_inData_62(switch_io_inData_62),
    .io_inData_63(switch_io_inData_63),
    .io_inValid_0(switch_io_inValid_0),
    .io_inValid_1(switch_io_inValid_1),
    .io_inValid_2(switch_io_inValid_2),
    .io_inValid_3(switch_io_inValid_3),
    .io_inValid_4(switch_io_inValid_4),
    .io_inValid_5(switch_io_inValid_5),
    .io_inValid_6(switch_io_inValid_6),
    .io_inValid_7(switch_io_inValid_7),
    .io_inValid_8(switch_io_inValid_8),
    .io_inValid_9(switch_io_inValid_9),
    .io_inValid_10(switch_io_inValid_10),
    .io_inValid_11(switch_io_inValid_11),
    .io_inValid_12(switch_io_inValid_12),
    .io_inValid_13(switch_io_inValid_13),
    .io_inValid_14(switch_io_inValid_14),
    .io_inValid_15(switch_io_inValid_15),
    .io_inValid_16(switch_io_inValid_16),
    .io_inValid_17(switch_io_inValid_17),
    .io_inValid_18(switch_io_inValid_18),
    .io_inValid_19(switch_io_inValid_19),
    .io_inValid_20(switch_io_inValid_20),
    .io_inValid_21(switch_io_inValid_21),
    .io_inValid_22(switch_io_inValid_22),
    .io_inValid_23(switch_io_inValid_23),
    .io_inValid_24(switch_io_inValid_24),
    .io_inValid_25(switch_io_inValid_25),
    .io_inValid_26(switch_io_inValid_26),
    .io_inValid_27(switch_io_inValid_27),
    .io_inValid_28(switch_io_inValid_28),
    .io_inValid_29(switch_io_inValid_29),
    .io_inValid_30(switch_io_inValid_30),
    .io_inValid_31(switch_io_inValid_31),
    .io_inValid_32(switch_io_inValid_32),
    .io_inValid_33(switch_io_inValid_33),
    .io_inValid_34(switch_io_inValid_34),
    .io_inValid_35(switch_io_inValid_35),
    .io_inValid_36(switch_io_inValid_36),
    .io_inValid_37(switch_io_inValid_37),
    .io_inValid_38(switch_io_inValid_38),
    .io_inValid_39(switch_io_inValid_39),
    .io_inValid_40(switch_io_inValid_40),
    .io_inValid_41(switch_io_inValid_41),
    .io_inValid_42(switch_io_inValid_42),
    .io_inValid_43(switch_io_inValid_43),
    .io_inValid_44(switch_io_inValid_44),
    .io_inValid_45(switch_io_inValid_45),
    .io_inValid_46(switch_io_inValid_46),
    .io_inValid_47(switch_io_inValid_47),
    .io_inValid_48(switch_io_inValid_48),
    .io_inValid_49(switch_io_inValid_49),
    .io_inValid_50(switch_io_inValid_50),
    .io_inValid_51(switch_io_inValid_51),
    .io_inValid_52(switch_io_inValid_52),
    .io_inValid_53(switch_io_inValid_53),
    .io_inValid_54(switch_io_inValid_54),
    .io_inValid_55(switch_io_inValid_55),
    .io_inValid_56(switch_io_inValid_56),
    .io_inValid_57(switch_io_inValid_57),
    .io_inValid_58(switch_io_inValid_58),
    .io_inValid_59(switch_io_inValid_59),
    .io_inValid_60(switch_io_inValid_60),
    .io_inValid_61(switch_io_inValid_61),
    .io_inValid_62(switch_io_inValid_62),
    .io_inValid_63(switch_io_inValid_63),
    .io_outAck_0(switch_io_outAck_0),
    .io_outAck_1(switch_io_outAck_1),
    .io_outAck_2(switch_io_outAck_2),
    .io_outAck_3(switch_io_outAck_3),
    .io_outAck_4(switch_io_outAck_4),
    .io_outAck_5(switch_io_outAck_5),
    .io_outAck_6(switch_io_outAck_6),
    .io_outAck_7(switch_io_outAck_7),
    .io_outAck_8(switch_io_outAck_8),
    .io_outAck_9(switch_io_outAck_9),
    .io_outAck_10(switch_io_outAck_10),
    .io_outAck_11(switch_io_outAck_11),
    .io_outAck_12(switch_io_outAck_12),
    .io_outAck_13(switch_io_outAck_13),
    .io_outAck_14(switch_io_outAck_14),
    .io_outAck_15(switch_io_outAck_15),
    .io_outAck_16(switch_io_outAck_16),
    .io_outAck_17(switch_io_outAck_17),
    .io_outAck_18(switch_io_outAck_18),
    .io_outAck_19(switch_io_outAck_19),
    .io_outAck_20(switch_io_outAck_20),
    .io_outAck_21(switch_io_outAck_21),
    .io_outAck_22(switch_io_outAck_22),
    .io_outAck_23(switch_io_outAck_23),
    .io_outAck_24(switch_io_outAck_24),
    .io_outAck_25(switch_io_outAck_25),
    .io_outAck_26(switch_io_outAck_26),
    .io_outAck_27(switch_io_outAck_27),
    .io_outAck_28(switch_io_outAck_28),
    .io_outAck_29(switch_io_outAck_29),
    .io_outAck_30(switch_io_outAck_30),
    .io_outAck_31(switch_io_outAck_31),
    .io_outAck_32(switch_io_outAck_32),
    .io_outAck_33(switch_io_outAck_33),
    .io_outAck_34(switch_io_outAck_34),
    .io_outAck_35(switch_io_outAck_35),
    .io_outAck_36(switch_io_outAck_36),
    .io_outAck_37(switch_io_outAck_37),
    .io_outAck_38(switch_io_outAck_38),
    .io_outAck_39(switch_io_outAck_39),
    .io_outAck_40(switch_io_outAck_40),
    .io_outAck_41(switch_io_outAck_41),
    .io_outAck_42(switch_io_outAck_42),
    .io_outAck_43(switch_io_outAck_43),
    .io_outAck_44(switch_io_outAck_44),
    .io_outAck_45(switch_io_outAck_45),
    .io_outAck_46(switch_io_outAck_46),
    .io_outAck_47(switch_io_outAck_47),
    .io_outAck_48(switch_io_outAck_48),
    .io_outAck_49(switch_io_outAck_49),
    .io_outAck_50(switch_io_outAck_50),
    .io_outAck_51(switch_io_outAck_51),
    .io_outAck_52(switch_io_outAck_52),
    .io_outAck_53(switch_io_outAck_53),
    .io_outAck_54(switch_io_outAck_54),
    .io_outAck_55(switch_io_outAck_55),
    .io_outAck_56(switch_io_outAck_56),
    .io_outAck_57(switch_io_outAck_57),
    .io_outAck_58(switch_io_outAck_58),
    .io_outAck_59(switch_io_outAck_59),
    .io_outAck_60(switch_io_outAck_60),
    .io_outAck_61(switch_io_outAck_61),
    .io_outAck_62(switch_io_outAck_62),
    .io_outAck_63(switch_io_outAck_63),
    .io_outData_0(switch_io_outData_0),
    .io_outData_1(switch_io_outData_1),
    .io_outData_2(switch_io_outData_2),
    .io_outData_3(switch_io_outData_3),
    .io_outData_4(switch_io_outData_4),
    .io_outData_5(switch_io_outData_5),
    .io_outData_6(switch_io_outData_6),
    .io_outData_7(switch_io_outData_7),
    .io_outData_8(switch_io_outData_8),
    .io_outData_9(switch_io_outData_9),
    .io_outData_10(switch_io_outData_10),
    .io_outData_11(switch_io_outData_11),
    .io_outData_12(switch_io_outData_12),
    .io_outData_13(switch_io_outData_13),
    .io_outData_14(switch_io_outData_14),
    .io_outData_15(switch_io_outData_15),
    .io_outData_16(switch_io_outData_16),
    .io_outData_17(switch_io_outData_17),
    .io_outData_18(switch_io_outData_18),
    .io_outData_19(switch_io_outData_19),
    .io_outData_20(switch_io_outData_20),
    .io_outData_21(switch_io_outData_21),
    .io_outData_22(switch_io_outData_22),
    .io_outData_23(switch_io_outData_23),
    .io_outData_24(switch_io_outData_24),
    .io_outData_25(switch_io_outData_25),
    .io_outData_26(switch_io_outData_26),
    .io_outData_27(switch_io_outData_27),
    .io_outData_28(switch_io_outData_28),
    .io_outData_29(switch_io_outData_29),
    .io_outData_30(switch_io_outData_30),
    .io_outData_31(switch_io_outData_31),
    .io_outData_32(switch_io_outData_32),
    .io_outData_33(switch_io_outData_33),
    .io_outData_34(switch_io_outData_34),
    .io_outData_35(switch_io_outData_35),
    .io_outData_36(switch_io_outData_36),
    .io_outData_37(switch_io_outData_37),
    .io_outData_38(switch_io_outData_38),
    .io_outData_39(switch_io_outData_39),
    .io_outData_40(switch_io_outData_40),
    .io_outData_41(switch_io_outData_41),
    .io_outData_42(switch_io_outData_42),
    .io_outData_43(switch_io_outData_43),
    .io_outData_44(switch_io_outData_44),
    .io_outData_45(switch_io_outData_45),
    .io_outData_46(switch_io_outData_46),
    .io_outData_47(switch_io_outData_47),
    .io_outData_48(switch_io_outData_48),
    .io_outData_49(switch_io_outData_49),
    .io_outData_50(switch_io_outData_50),
    .io_outData_51(switch_io_outData_51),
    .io_outData_52(switch_io_outData_52),
    .io_outData_53(switch_io_outData_53),
    .io_outData_54(switch_io_outData_54),
    .io_outData_55(switch_io_outData_55),
    .io_outData_56(switch_io_outData_56),
    .io_outData_57(switch_io_outData_57),
    .io_outData_58(switch_io_outData_58),
    .io_outData_59(switch_io_outData_59),
    .io_outData_60(switch_io_outData_60),
    .io_outData_61(switch_io_outData_61),
    .io_outData_62(switch_io_outData_62),
    .io_outData_63(switch_io_outData_63),
    .io_outValid_0(switch_io_outValid_0),
    .io_outValid_1(switch_io_outValid_1),
    .io_outValid_2(switch_io_outValid_2),
    .io_outValid_3(switch_io_outValid_3),
    .io_outValid_4(switch_io_outValid_4),
    .io_outValid_5(switch_io_outValid_5),
    .io_outValid_6(switch_io_outValid_6),
    .io_outValid_7(switch_io_outValid_7),
    .io_outValid_8(switch_io_outValid_8),
    .io_outValid_9(switch_io_outValid_9),
    .io_outValid_10(switch_io_outValid_10),
    .io_outValid_11(switch_io_outValid_11),
    .io_outValid_12(switch_io_outValid_12),
    .io_outValid_13(switch_io_outValid_13),
    .io_outValid_14(switch_io_outValid_14),
    .io_outValid_15(switch_io_outValid_15),
    .io_outValid_16(switch_io_outValid_16),
    .io_outValid_17(switch_io_outValid_17),
    .io_outValid_18(switch_io_outValid_18),
    .io_outValid_19(switch_io_outValid_19),
    .io_outValid_20(switch_io_outValid_20),
    .io_outValid_21(switch_io_outValid_21),
    .io_outValid_22(switch_io_outValid_22),
    .io_outValid_23(switch_io_outValid_23),
    .io_outValid_24(switch_io_outValid_24),
    .io_outValid_25(switch_io_outValid_25),
    .io_outValid_26(switch_io_outValid_26),
    .io_outValid_27(switch_io_outValid_27),
    .io_outValid_28(switch_io_outValid_28),
    .io_outValid_29(switch_io_outValid_29),
    .io_outValid_30(switch_io_outValid_30),
    .io_outValid_31(switch_io_outValid_31),
    .io_outValid_32(switch_io_outValid_32),
    .io_outValid_33(switch_io_outValid_33),
    .io_outValid_34(switch_io_outValid_34),
    .io_outValid_35(switch_io_outValid_35),
    .io_outValid_36(switch_io_outValid_36),
    .io_outValid_37(switch_io_outValid_37),
    .io_outValid_38(switch_io_outValid_38),
    .io_outValid_39(switch_io_outValid_39),
    .io_outValid_40(switch_io_outValid_40),
    .io_outValid_41(switch_io_outValid_41),
    .io_outValid_42(switch_io_outValid_42),
    .io_outValid_43(switch_io_outValid_43),
    .io_outValid_44(switch_io_outValid_44),
    .io_outValid_45(switch_io_outValid_45),
    .io_outValid_46(switch_io_outValid_46),
    .io_outValid_47(switch_io_outValid_47),
    .io_outValid_48(switch_io_outValid_48),
    .io_outValid_49(switch_io_outValid_49),
    .io_outValid_50(switch_io_outValid_50),
    .io_outValid_51(switch_io_outValid_51),
    .io_outValid_52(switch_io_outValid_52),
    .io_outValid_53(switch_io_outValid_53),
    .io_outValid_54(switch_io_outValid_54),
    .io_outValid_55(switch_io_outValid_55),
    .io_outValid_56(switch_io_outValid_56),
    .io_outValid_57(switch_io_outValid_57),
    .io_outValid_58(switch_io_outValid_58),
    .io_outValid_59(switch_io_outValid_59),
    .io_outValid_60(switch_io_outValid_60),
    .io_outValid_61(switch_io_outValid_61),
    .io_outValid_62(switch_io_outValid_62),
    .io_outValid_63(switch_io_outValid_63)
  );
  assign io_outAck_0 = _T_1537_0; // @[Switch.scala 54:13:@37528.4]
  assign io_outAck_1 = _T_1537_1; // @[Switch.scala 54:13:@37529.4]
  assign io_outAck_2 = _T_1537_2; // @[Switch.scala 54:13:@37530.4]
  assign io_outAck_3 = _T_1537_3; // @[Switch.scala 54:13:@37531.4]
  assign io_outAck_4 = _T_1537_4; // @[Switch.scala 54:13:@37532.4]
  assign io_outAck_5 = _T_1537_5; // @[Switch.scala 54:13:@37533.4]
  assign io_outAck_6 = _T_1537_6; // @[Switch.scala 54:13:@37534.4]
  assign io_outAck_7 = _T_1537_7; // @[Switch.scala 54:13:@37535.4]
  assign io_outAck_8 = _T_1537_8; // @[Switch.scala 54:13:@37536.4]
  assign io_outAck_9 = _T_1537_9; // @[Switch.scala 54:13:@37537.4]
  assign io_outAck_10 = _T_1537_10; // @[Switch.scala 54:13:@37538.4]
  assign io_outAck_11 = _T_1537_11; // @[Switch.scala 54:13:@37539.4]
  assign io_outAck_12 = _T_1537_12; // @[Switch.scala 54:13:@37540.4]
  assign io_outAck_13 = _T_1537_13; // @[Switch.scala 54:13:@37541.4]
  assign io_outAck_14 = _T_1537_14; // @[Switch.scala 54:13:@37542.4]
  assign io_outAck_15 = _T_1537_15; // @[Switch.scala 54:13:@37543.4]
  assign io_outAck_16 = _T_1537_16; // @[Switch.scala 54:13:@37544.4]
  assign io_outAck_17 = _T_1537_17; // @[Switch.scala 54:13:@37545.4]
  assign io_outAck_18 = _T_1537_18; // @[Switch.scala 54:13:@37546.4]
  assign io_outAck_19 = _T_1537_19; // @[Switch.scala 54:13:@37547.4]
  assign io_outAck_20 = _T_1537_20; // @[Switch.scala 54:13:@37548.4]
  assign io_outAck_21 = _T_1537_21; // @[Switch.scala 54:13:@37549.4]
  assign io_outAck_22 = _T_1537_22; // @[Switch.scala 54:13:@37550.4]
  assign io_outAck_23 = _T_1537_23; // @[Switch.scala 54:13:@37551.4]
  assign io_outAck_24 = _T_1537_24; // @[Switch.scala 54:13:@37552.4]
  assign io_outAck_25 = _T_1537_25; // @[Switch.scala 54:13:@37553.4]
  assign io_outAck_26 = _T_1537_26; // @[Switch.scala 54:13:@37554.4]
  assign io_outAck_27 = _T_1537_27; // @[Switch.scala 54:13:@37555.4]
  assign io_outAck_28 = _T_1537_28; // @[Switch.scala 54:13:@37556.4]
  assign io_outAck_29 = _T_1537_29; // @[Switch.scala 54:13:@37557.4]
  assign io_outAck_30 = _T_1537_30; // @[Switch.scala 54:13:@37558.4]
  assign io_outAck_31 = _T_1537_31; // @[Switch.scala 54:13:@37559.4]
  assign io_outAck_32 = _T_1537_32; // @[Switch.scala 54:13:@37560.4]
  assign io_outAck_33 = _T_1537_33; // @[Switch.scala 54:13:@37561.4]
  assign io_outAck_34 = _T_1537_34; // @[Switch.scala 54:13:@37562.4]
  assign io_outAck_35 = _T_1537_35; // @[Switch.scala 54:13:@37563.4]
  assign io_outAck_36 = _T_1537_36; // @[Switch.scala 54:13:@37564.4]
  assign io_outAck_37 = _T_1537_37; // @[Switch.scala 54:13:@37565.4]
  assign io_outAck_38 = _T_1537_38; // @[Switch.scala 54:13:@37566.4]
  assign io_outAck_39 = _T_1537_39; // @[Switch.scala 54:13:@37567.4]
  assign io_outAck_40 = _T_1537_40; // @[Switch.scala 54:13:@37568.4]
  assign io_outAck_41 = _T_1537_41; // @[Switch.scala 54:13:@37569.4]
  assign io_outAck_42 = _T_1537_42; // @[Switch.scala 54:13:@37570.4]
  assign io_outAck_43 = _T_1537_43; // @[Switch.scala 54:13:@37571.4]
  assign io_outAck_44 = _T_1537_44; // @[Switch.scala 54:13:@37572.4]
  assign io_outAck_45 = _T_1537_45; // @[Switch.scala 54:13:@37573.4]
  assign io_outAck_46 = _T_1537_46; // @[Switch.scala 54:13:@37574.4]
  assign io_outAck_47 = _T_1537_47; // @[Switch.scala 54:13:@37575.4]
  assign io_outAck_48 = _T_1537_48; // @[Switch.scala 54:13:@37576.4]
  assign io_outAck_49 = _T_1537_49; // @[Switch.scala 54:13:@37577.4]
  assign io_outAck_50 = _T_1537_50; // @[Switch.scala 54:13:@37578.4]
  assign io_outAck_51 = _T_1537_51; // @[Switch.scala 54:13:@37579.4]
  assign io_outAck_52 = _T_1537_52; // @[Switch.scala 54:13:@37580.4]
  assign io_outAck_53 = _T_1537_53; // @[Switch.scala 54:13:@37581.4]
  assign io_outAck_54 = _T_1537_54; // @[Switch.scala 54:13:@37582.4]
  assign io_outAck_55 = _T_1537_55; // @[Switch.scala 54:13:@37583.4]
  assign io_outAck_56 = _T_1537_56; // @[Switch.scala 54:13:@37584.4]
  assign io_outAck_57 = _T_1537_57; // @[Switch.scala 54:13:@37585.4]
  assign io_outAck_58 = _T_1537_58; // @[Switch.scala 54:13:@37586.4]
  assign io_outAck_59 = _T_1537_59; // @[Switch.scala 54:13:@37587.4]
  assign io_outAck_60 = _T_1537_60; // @[Switch.scala 54:13:@37588.4]
  assign io_outAck_61 = _T_1537_61; // @[Switch.scala 54:13:@37589.4]
  assign io_outAck_62 = _T_1537_62; // @[Switch.scala 54:13:@37590.4]
  assign io_outAck_63 = _T_1537_63; // @[Switch.scala 54:13:@37591.4]
  assign io_outData_0 = _T_1866_0; // @[Switch.scala 55:14:@37657.4]
  assign io_outData_1 = _T_1866_1; // @[Switch.scala 55:14:@37658.4]
  assign io_outData_2 = _T_1866_2; // @[Switch.scala 55:14:@37659.4]
  assign io_outData_3 = _T_1866_3; // @[Switch.scala 55:14:@37660.4]
  assign io_outData_4 = _T_1866_4; // @[Switch.scala 55:14:@37661.4]
  assign io_outData_5 = _T_1866_5; // @[Switch.scala 55:14:@37662.4]
  assign io_outData_6 = _T_1866_6; // @[Switch.scala 55:14:@37663.4]
  assign io_outData_7 = _T_1866_7; // @[Switch.scala 55:14:@37664.4]
  assign io_outData_8 = _T_1866_8; // @[Switch.scala 55:14:@37665.4]
  assign io_outData_9 = _T_1866_9; // @[Switch.scala 55:14:@37666.4]
  assign io_outData_10 = _T_1866_10; // @[Switch.scala 55:14:@37667.4]
  assign io_outData_11 = _T_1866_11; // @[Switch.scala 55:14:@37668.4]
  assign io_outData_12 = _T_1866_12; // @[Switch.scala 55:14:@37669.4]
  assign io_outData_13 = _T_1866_13; // @[Switch.scala 55:14:@37670.4]
  assign io_outData_14 = _T_1866_14; // @[Switch.scala 55:14:@37671.4]
  assign io_outData_15 = _T_1866_15; // @[Switch.scala 55:14:@37672.4]
  assign io_outData_16 = _T_1866_16; // @[Switch.scala 55:14:@37673.4]
  assign io_outData_17 = _T_1866_17; // @[Switch.scala 55:14:@37674.4]
  assign io_outData_18 = _T_1866_18; // @[Switch.scala 55:14:@37675.4]
  assign io_outData_19 = _T_1866_19; // @[Switch.scala 55:14:@37676.4]
  assign io_outData_20 = _T_1866_20; // @[Switch.scala 55:14:@37677.4]
  assign io_outData_21 = _T_1866_21; // @[Switch.scala 55:14:@37678.4]
  assign io_outData_22 = _T_1866_22; // @[Switch.scala 55:14:@37679.4]
  assign io_outData_23 = _T_1866_23; // @[Switch.scala 55:14:@37680.4]
  assign io_outData_24 = _T_1866_24; // @[Switch.scala 55:14:@37681.4]
  assign io_outData_25 = _T_1866_25; // @[Switch.scala 55:14:@37682.4]
  assign io_outData_26 = _T_1866_26; // @[Switch.scala 55:14:@37683.4]
  assign io_outData_27 = _T_1866_27; // @[Switch.scala 55:14:@37684.4]
  assign io_outData_28 = _T_1866_28; // @[Switch.scala 55:14:@37685.4]
  assign io_outData_29 = _T_1866_29; // @[Switch.scala 55:14:@37686.4]
  assign io_outData_30 = _T_1866_30; // @[Switch.scala 55:14:@37687.4]
  assign io_outData_31 = _T_1866_31; // @[Switch.scala 55:14:@37688.4]
  assign io_outData_32 = _T_1866_32; // @[Switch.scala 55:14:@37689.4]
  assign io_outData_33 = _T_1866_33; // @[Switch.scala 55:14:@37690.4]
  assign io_outData_34 = _T_1866_34; // @[Switch.scala 55:14:@37691.4]
  assign io_outData_35 = _T_1866_35; // @[Switch.scala 55:14:@37692.4]
  assign io_outData_36 = _T_1866_36; // @[Switch.scala 55:14:@37693.4]
  assign io_outData_37 = _T_1866_37; // @[Switch.scala 55:14:@37694.4]
  assign io_outData_38 = _T_1866_38; // @[Switch.scala 55:14:@37695.4]
  assign io_outData_39 = _T_1866_39; // @[Switch.scala 55:14:@37696.4]
  assign io_outData_40 = _T_1866_40; // @[Switch.scala 55:14:@37697.4]
  assign io_outData_41 = _T_1866_41; // @[Switch.scala 55:14:@37698.4]
  assign io_outData_42 = _T_1866_42; // @[Switch.scala 55:14:@37699.4]
  assign io_outData_43 = _T_1866_43; // @[Switch.scala 55:14:@37700.4]
  assign io_outData_44 = _T_1866_44; // @[Switch.scala 55:14:@37701.4]
  assign io_outData_45 = _T_1866_45; // @[Switch.scala 55:14:@37702.4]
  assign io_outData_46 = _T_1866_46; // @[Switch.scala 55:14:@37703.4]
  assign io_outData_47 = _T_1866_47; // @[Switch.scala 55:14:@37704.4]
  assign io_outData_48 = _T_1866_48; // @[Switch.scala 55:14:@37705.4]
  assign io_outData_49 = _T_1866_49; // @[Switch.scala 55:14:@37706.4]
  assign io_outData_50 = _T_1866_50; // @[Switch.scala 55:14:@37707.4]
  assign io_outData_51 = _T_1866_51; // @[Switch.scala 55:14:@37708.4]
  assign io_outData_52 = _T_1866_52; // @[Switch.scala 55:14:@37709.4]
  assign io_outData_53 = _T_1866_53; // @[Switch.scala 55:14:@37710.4]
  assign io_outData_54 = _T_1866_54; // @[Switch.scala 55:14:@37711.4]
  assign io_outData_55 = _T_1866_55; // @[Switch.scala 55:14:@37712.4]
  assign io_outData_56 = _T_1866_56; // @[Switch.scala 55:14:@37713.4]
  assign io_outData_57 = _T_1866_57; // @[Switch.scala 55:14:@37714.4]
  assign io_outData_58 = _T_1866_58; // @[Switch.scala 55:14:@37715.4]
  assign io_outData_59 = _T_1866_59; // @[Switch.scala 55:14:@37716.4]
  assign io_outData_60 = _T_1866_60; // @[Switch.scala 55:14:@37717.4]
  assign io_outData_61 = _T_1866_61; // @[Switch.scala 55:14:@37718.4]
  assign io_outData_62 = _T_1866_62; // @[Switch.scala 55:14:@37719.4]
  assign io_outData_63 = _T_1866_63; // @[Switch.scala 55:14:@37720.4]
  assign io_outValid_0 = _T_2195_0; // @[Switch.scala 56:15:@37786.4]
  assign io_outValid_1 = _T_2195_1; // @[Switch.scala 56:15:@37787.4]
  assign io_outValid_2 = _T_2195_2; // @[Switch.scala 56:15:@37788.4]
  assign io_outValid_3 = _T_2195_3; // @[Switch.scala 56:15:@37789.4]
  assign io_outValid_4 = _T_2195_4; // @[Switch.scala 56:15:@37790.4]
  assign io_outValid_5 = _T_2195_5; // @[Switch.scala 56:15:@37791.4]
  assign io_outValid_6 = _T_2195_6; // @[Switch.scala 56:15:@37792.4]
  assign io_outValid_7 = _T_2195_7; // @[Switch.scala 56:15:@37793.4]
  assign io_outValid_8 = _T_2195_8; // @[Switch.scala 56:15:@37794.4]
  assign io_outValid_9 = _T_2195_9; // @[Switch.scala 56:15:@37795.4]
  assign io_outValid_10 = _T_2195_10; // @[Switch.scala 56:15:@37796.4]
  assign io_outValid_11 = _T_2195_11; // @[Switch.scala 56:15:@37797.4]
  assign io_outValid_12 = _T_2195_12; // @[Switch.scala 56:15:@37798.4]
  assign io_outValid_13 = _T_2195_13; // @[Switch.scala 56:15:@37799.4]
  assign io_outValid_14 = _T_2195_14; // @[Switch.scala 56:15:@37800.4]
  assign io_outValid_15 = _T_2195_15; // @[Switch.scala 56:15:@37801.4]
  assign io_outValid_16 = _T_2195_16; // @[Switch.scala 56:15:@37802.4]
  assign io_outValid_17 = _T_2195_17; // @[Switch.scala 56:15:@37803.4]
  assign io_outValid_18 = _T_2195_18; // @[Switch.scala 56:15:@37804.4]
  assign io_outValid_19 = _T_2195_19; // @[Switch.scala 56:15:@37805.4]
  assign io_outValid_20 = _T_2195_20; // @[Switch.scala 56:15:@37806.4]
  assign io_outValid_21 = _T_2195_21; // @[Switch.scala 56:15:@37807.4]
  assign io_outValid_22 = _T_2195_22; // @[Switch.scala 56:15:@37808.4]
  assign io_outValid_23 = _T_2195_23; // @[Switch.scala 56:15:@37809.4]
  assign io_outValid_24 = _T_2195_24; // @[Switch.scala 56:15:@37810.4]
  assign io_outValid_25 = _T_2195_25; // @[Switch.scala 56:15:@37811.4]
  assign io_outValid_26 = _T_2195_26; // @[Switch.scala 56:15:@37812.4]
  assign io_outValid_27 = _T_2195_27; // @[Switch.scala 56:15:@37813.4]
  assign io_outValid_28 = _T_2195_28; // @[Switch.scala 56:15:@37814.4]
  assign io_outValid_29 = _T_2195_29; // @[Switch.scala 56:15:@37815.4]
  assign io_outValid_30 = _T_2195_30; // @[Switch.scala 56:15:@37816.4]
  assign io_outValid_31 = _T_2195_31; // @[Switch.scala 56:15:@37817.4]
  assign io_outValid_32 = _T_2195_32; // @[Switch.scala 56:15:@37818.4]
  assign io_outValid_33 = _T_2195_33; // @[Switch.scala 56:15:@37819.4]
  assign io_outValid_34 = _T_2195_34; // @[Switch.scala 56:15:@37820.4]
  assign io_outValid_35 = _T_2195_35; // @[Switch.scala 56:15:@37821.4]
  assign io_outValid_36 = _T_2195_36; // @[Switch.scala 56:15:@37822.4]
  assign io_outValid_37 = _T_2195_37; // @[Switch.scala 56:15:@37823.4]
  assign io_outValid_38 = _T_2195_38; // @[Switch.scala 56:15:@37824.4]
  assign io_outValid_39 = _T_2195_39; // @[Switch.scala 56:15:@37825.4]
  assign io_outValid_40 = _T_2195_40; // @[Switch.scala 56:15:@37826.4]
  assign io_outValid_41 = _T_2195_41; // @[Switch.scala 56:15:@37827.4]
  assign io_outValid_42 = _T_2195_42; // @[Switch.scala 56:15:@37828.4]
  assign io_outValid_43 = _T_2195_43; // @[Switch.scala 56:15:@37829.4]
  assign io_outValid_44 = _T_2195_44; // @[Switch.scala 56:15:@37830.4]
  assign io_outValid_45 = _T_2195_45; // @[Switch.scala 56:15:@37831.4]
  assign io_outValid_46 = _T_2195_46; // @[Switch.scala 56:15:@37832.4]
  assign io_outValid_47 = _T_2195_47; // @[Switch.scala 56:15:@37833.4]
  assign io_outValid_48 = _T_2195_48; // @[Switch.scala 56:15:@37834.4]
  assign io_outValid_49 = _T_2195_49; // @[Switch.scala 56:15:@37835.4]
  assign io_outValid_50 = _T_2195_50; // @[Switch.scala 56:15:@37836.4]
  assign io_outValid_51 = _T_2195_51; // @[Switch.scala 56:15:@37837.4]
  assign io_outValid_52 = _T_2195_52; // @[Switch.scala 56:15:@37838.4]
  assign io_outValid_53 = _T_2195_53; // @[Switch.scala 56:15:@37839.4]
  assign io_outValid_54 = _T_2195_54; // @[Switch.scala 56:15:@37840.4]
  assign io_outValid_55 = _T_2195_55; // @[Switch.scala 56:15:@37841.4]
  assign io_outValid_56 = _T_2195_56; // @[Switch.scala 56:15:@37842.4]
  assign io_outValid_57 = _T_2195_57; // @[Switch.scala 56:15:@37843.4]
  assign io_outValid_58 = _T_2195_58; // @[Switch.scala 56:15:@37844.4]
  assign io_outValid_59 = _T_2195_59; // @[Switch.scala 56:15:@37845.4]
  assign io_outValid_60 = _T_2195_60; // @[Switch.scala 56:15:@37846.4]
  assign io_outValid_61 = _T_2195_61; // @[Switch.scala 56:15:@37847.4]
  assign io_outValid_62 = _T_2195_62; // @[Switch.scala 56:15:@37848.4]
  assign io_outValid_63 = _T_2195_63; // @[Switch.scala 56:15:@37849.4]
  assign switch_io_inAddr_0 = _T_550_0; // @[Switch.scala 51:20:@37141.4]
  assign switch_io_inAddr_1 = _T_550_1; // @[Switch.scala 51:20:@37142.4]
  assign switch_io_inAddr_2 = _T_550_2; // @[Switch.scala 51:20:@37143.4]
  assign switch_io_inAddr_3 = _T_550_3; // @[Switch.scala 51:20:@37144.4]
  assign switch_io_inAddr_4 = _T_550_4; // @[Switch.scala 51:20:@37145.4]
  assign switch_io_inAddr_5 = _T_550_5; // @[Switch.scala 51:20:@37146.4]
  assign switch_io_inAddr_6 = _T_550_6; // @[Switch.scala 51:20:@37147.4]
  assign switch_io_inAddr_7 = _T_550_7; // @[Switch.scala 51:20:@37148.4]
  assign switch_io_inAddr_8 = _T_550_8; // @[Switch.scala 51:20:@37149.4]
  assign switch_io_inAddr_9 = _T_550_9; // @[Switch.scala 51:20:@37150.4]
  assign switch_io_inAddr_10 = _T_550_10; // @[Switch.scala 51:20:@37151.4]
  assign switch_io_inAddr_11 = _T_550_11; // @[Switch.scala 51:20:@37152.4]
  assign switch_io_inAddr_12 = _T_550_12; // @[Switch.scala 51:20:@37153.4]
  assign switch_io_inAddr_13 = _T_550_13; // @[Switch.scala 51:20:@37154.4]
  assign switch_io_inAddr_14 = _T_550_14; // @[Switch.scala 51:20:@37155.4]
  assign switch_io_inAddr_15 = _T_550_15; // @[Switch.scala 51:20:@37156.4]
  assign switch_io_inAddr_16 = _T_550_16; // @[Switch.scala 51:20:@37157.4]
  assign switch_io_inAddr_17 = _T_550_17; // @[Switch.scala 51:20:@37158.4]
  assign switch_io_inAddr_18 = _T_550_18; // @[Switch.scala 51:20:@37159.4]
  assign switch_io_inAddr_19 = _T_550_19; // @[Switch.scala 51:20:@37160.4]
  assign switch_io_inAddr_20 = _T_550_20; // @[Switch.scala 51:20:@37161.4]
  assign switch_io_inAddr_21 = _T_550_21; // @[Switch.scala 51:20:@37162.4]
  assign switch_io_inAddr_22 = _T_550_22; // @[Switch.scala 51:20:@37163.4]
  assign switch_io_inAddr_23 = _T_550_23; // @[Switch.scala 51:20:@37164.4]
  assign switch_io_inAddr_24 = _T_550_24; // @[Switch.scala 51:20:@37165.4]
  assign switch_io_inAddr_25 = _T_550_25; // @[Switch.scala 51:20:@37166.4]
  assign switch_io_inAddr_26 = _T_550_26; // @[Switch.scala 51:20:@37167.4]
  assign switch_io_inAddr_27 = _T_550_27; // @[Switch.scala 51:20:@37168.4]
  assign switch_io_inAddr_28 = _T_550_28; // @[Switch.scala 51:20:@37169.4]
  assign switch_io_inAddr_29 = _T_550_29; // @[Switch.scala 51:20:@37170.4]
  assign switch_io_inAddr_30 = _T_550_30; // @[Switch.scala 51:20:@37171.4]
  assign switch_io_inAddr_31 = _T_550_31; // @[Switch.scala 51:20:@37172.4]
  assign switch_io_inAddr_32 = _T_550_32; // @[Switch.scala 51:20:@37173.4]
  assign switch_io_inAddr_33 = _T_550_33; // @[Switch.scala 51:20:@37174.4]
  assign switch_io_inAddr_34 = _T_550_34; // @[Switch.scala 51:20:@37175.4]
  assign switch_io_inAddr_35 = _T_550_35; // @[Switch.scala 51:20:@37176.4]
  assign switch_io_inAddr_36 = _T_550_36; // @[Switch.scala 51:20:@37177.4]
  assign switch_io_inAddr_37 = _T_550_37; // @[Switch.scala 51:20:@37178.4]
  assign switch_io_inAddr_38 = _T_550_38; // @[Switch.scala 51:20:@37179.4]
  assign switch_io_inAddr_39 = _T_550_39; // @[Switch.scala 51:20:@37180.4]
  assign switch_io_inAddr_40 = _T_550_40; // @[Switch.scala 51:20:@37181.4]
  assign switch_io_inAddr_41 = _T_550_41; // @[Switch.scala 51:20:@37182.4]
  assign switch_io_inAddr_42 = _T_550_42; // @[Switch.scala 51:20:@37183.4]
  assign switch_io_inAddr_43 = _T_550_43; // @[Switch.scala 51:20:@37184.4]
  assign switch_io_inAddr_44 = _T_550_44; // @[Switch.scala 51:20:@37185.4]
  assign switch_io_inAddr_45 = _T_550_45; // @[Switch.scala 51:20:@37186.4]
  assign switch_io_inAddr_46 = _T_550_46; // @[Switch.scala 51:20:@37187.4]
  assign switch_io_inAddr_47 = _T_550_47; // @[Switch.scala 51:20:@37188.4]
  assign switch_io_inAddr_48 = _T_550_48; // @[Switch.scala 51:20:@37189.4]
  assign switch_io_inAddr_49 = _T_550_49; // @[Switch.scala 51:20:@37190.4]
  assign switch_io_inAddr_50 = _T_550_50; // @[Switch.scala 51:20:@37191.4]
  assign switch_io_inAddr_51 = _T_550_51; // @[Switch.scala 51:20:@37192.4]
  assign switch_io_inAddr_52 = _T_550_52; // @[Switch.scala 51:20:@37193.4]
  assign switch_io_inAddr_53 = _T_550_53; // @[Switch.scala 51:20:@37194.4]
  assign switch_io_inAddr_54 = _T_550_54; // @[Switch.scala 51:20:@37195.4]
  assign switch_io_inAddr_55 = _T_550_55; // @[Switch.scala 51:20:@37196.4]
  assign switch_io_inAddr_56 = _T_550_56; // @[Switch.scala 51:20:@37197.4]
  assign switch_io_inAddr_57 = _T_550_57; // @[Switch.scala 51:20:@37198.4]
  assign switch_io_inAddr_58 = _T_550_58; // @[Switch.scala 51:20:@37199.4]
  assign switch_io_inAddr_59 = _T_550_59; // @[Switch.scala 51:20:@37200.4]
  assign switch_io_inAddr_60 = _T_550_60; // @[Switch.scala 51:20:@37201.4]
  assign switch_io_inAddr_61 = _T_550_61; // @[Switch.scala 51:20:@37202.4]
  assign switch_io_inAddr_62 = _T_550_62; // @[Switch.scala 51:20:@37203.4]
  assign switch_io_inAddr_63 = _T_550_63; // @[Switch.scala 51:20:@37204.4]
  assign switch_io_inData_0 = _T_879_0; // @[Switch.scala 52:20:@37270.4]
  assign switch_io_inData_1 = _T_879_1; // @[Switch.scala 52:20:@37271.4]
  assign switch_io_inData_2 = _T_879_2; // @[Switch.scala 52:20:@37272.4]
  assign switch_io_inData_3 = _T_879_3; // @[Switch.scala 52:20:@37273.4]
  assign switch_io_inData_4 = _T_879_4; // @[Switch.scala 52:20:@37274.4]
  assign switch_io_inData_5 = _T_879_5; // @[Switch.scala 52:20:@37275.4]
  assign switch_io_inData_6 = _T_879_6; // @[Switch.scala 52:20:@37276.4]
  assign switch_io_inData_7 = _T_879_7; // @[Switch.scala 52:20:@37277.4]
  assign switch_io_inData_8 = _T_879_8; // @[Switch.scala 52:20:@37278.4]
  assign switch_io_inData_9 = _T_879_9; // @[Switch.scala 52:20:@37279.4]
  assign switch_io_inData_10 = _T_879_10; // @[Switch.scala 52:20:@37280.4]
  assign switch_io_inData_11 = _T_879_11; // @[Switch.scala 52:20:@37281.4]
  assign switch_io_inData_12 = _T_879_12; // @[Switch.scala 52:20:@37282.4]
  assign switch_io_inData_13 = _T_879_13; // @[Switch.scala 52:20:@37283.4]
  assign switch_io_inData_14 = _T_879_14; // @[Switch.scala 52:20:@37284.4]
  assign switch_io_inData_15 = _T_879_15; // @[Switch.scala 52:20:@37285.4]
  assign switch_io_inData_16 = _T_879_16; // @[Switch.scala 52:20:@37286.4]
  assign switch_io_inData_17 = _T_879_17; // @[Switch.scala 52:20:@37287.4]
  assign switch_io_inData_18 = _T_879_18; // @[Switch.scala 52:20:@37288.4]
  assign switch_io_inData_19 = _T_879_19; // @[Switch.scala 52:20:@37289.4]
  assign switch_io_inData_20 = _T_879_20; // @[Switch.scala 52:20:@37290.4]
  assign switch_io_inData_21 = _T_879_21; // @[Switch.scala 52:20:@37291.4]
  assign switch_io_inData_22 = _T_879_22; // @[Switch.scala 52:20:@37292.4]
  assign switch_io_inData_23 = _T_879_23; // @[Switch.scala 52:20:@37293.4]
  assign switch_io_inData_24 = _T_879_24; // @[Switch.scala 52:20:@37294.4]
  assign switch_io_inData_25 = _T_879_25; // @[Switch.scala 52:20:@37295.4]
  assign switch_io_inData_26 = _T_879_26; // @[Switch.scala 52:20:@37296.4]
  assign switch_io_inData_27 = _T_879_27; // @[Switch.scala 52:20:@37297.4]
  assign switch_io_inData_28 = _T_879_28; // @[Switch.scala 52:20:@37298.4]
  assign switch_io_inData_29 = _T_879_29; // @[Switch.scala 52:20:@37299.4]
  assign switch_io_inData_30 = _T_879_30; // @[Switch.scala 52:20:@37300.4]
  assign switch_io_inData_31 = _T_879_31; // @[Switch.scala 52:20:@37301.4]
  assign switch_io_inData_32 = _T_879_32; // @[Switch.scala 52:20:@37302.4]
  assign switch_io_inData_33 = _T_879_33; // @[Switch.scala 52:20:@37303.4]
  assign switch_io_inData_34 = _T_879_34; // @[Switch.scala 52:20:@37304.4]
  assign switch_io_inData_35 = _T_879_35; // @[Switch.scala 52:20:@37305.4]
  assign switch_io_inData_36 = _T_879_36; // @[Switch.scala 52:20:@37306.4]
  assign switch_io_inData_37 = _T_879_37; // @[Switch.scala 52:20:@37307.4]
  assign switch_io_inData_38 = _T_879_38; // @[Switch.scala 52:20:@37308.4]
  assign switch_io_inData_39 = _T_879_39; // @[Switch.scala 52:20:@37309.4]
  assign switch_io_inData_40 = _T_879_40; // @[Switch.scala 52:20:@37310.4]
  assign switch_io_inData_41 = _T_879_41; // @[Switch.scala 52:20:@37311.4]
  assign switch_io_inData_42 = _T_879_42; // @[Switch.scala 52:20:@37312.4]
  assign switch_io_inData_43 = _T_879_43; // @[Switch.scala 52:20:@37313.4]
  assign switch_io_inData_44 = _T_879_44; // @[Switch.scala 52:20:@37314.4]
  assign switch_io_inData_45 = _T_879_45; // @[Switch.scala 52:20:@37315.4]
  assign switch_io_inData_46 = _T_879_46; // @[Switch.scala 52:20:@37316.4]
  assign switch_io_inData_47 = _T_879_47; // @[Switch.scala 52:20:@37317.4]
  assign switch_io_inData_48 = _T_879_48; // @[Switch.scala 52:20:@37318.4]
  assign switch_io_inData_49 = _T_879_49; // @[Switch.scala 52:20:@37319.4]
  assign switch_io_inData_50 = _T_879_50; // @[Switch.scala 52:20:@37320.4]
  assign switch_io_inData_51 = _T_879_51; // @[Switch.scala 52:20:@37321.4]
  assign switch_io_inData_52 = _T_879_52; // @[Switch.scala 52:20:@37322.4]
  assign switch_io_inData_53 = _T_879_53; // @[Switch.scala 52:20:@37323.4]
  assign switch_io_inData_54 = _T_879_54; // @[Switch.scala 52:20:@37324.4]
  assign switch_io_inData_55 = _T_879_55; // @[Switch.scala 52:20:@37325.4]
  assign switch_io_inData_56 = _T_879_56; // @[Switch.scala 52:20:@37326.4]
  assign switch_io_inData_57 = _T_879_57; // @[Switch.scala 52:20:@37327.4]
  assign switch_io_inData_58 = _T_879_58; // @[Switch.scala 52:20:@37328.4]
  assign switch_io_inData_59 = _T_879_59; // @[Switch.scala 52:20:@37329.4]
  assign switch_io_inData_60 = _T_879_60; // @[Switch.scala 52:20:@37330.4]
  assign switch_io_inData_61 = _T_879_61; // @[Switch.scala 52:20:@37331.4]
  assign switch_io_inData_62 = _T_879_62; // @[Switch.scala 52:20:@37332.4]
  assign switch_io_inData_63 = _T_879_63; // @[Switch.scala 52:20:@37333.4]
  assign switch_io_inValid_0 = _T_1208_0; // @[Switch.scala 53:21:@37399.4]
  assign switch_io_inValid_1 = _T_1208_1; // @[Switch.scala 53:21:@37400.4]
  assign switch_io_inValid_2 = _T_1208_2; // @[Switch.scala 53:21:@37401.4]
  assign switch_io_inValid_3 = _T_1208_3; // @[Switch.scala 53:21:@37402.4]
  assign switch_io_inValid_4 = _T_1208_4; // @[Switch.scala 53:21:@37403.4]
  assign switch_io_inValid_5 = _T_1208_5; // @[Switch.scala 53:21:@37404.4]
  assign switch_io_inValid_6 = _T_1208_6; // @[Switch.scala 53:21:@37405.4]
  assign switch_io_inValid_7 = _T_1208_7; // @[Switch.scala 53:21:@37406.4]
  assign switch_io_inValid_8 = _T_1208_8; // @[Switch.scala 53:21:@37407.4]
  assign switch_io_inValid_9 = _T_1208_9; // @[Switch.scala 53:21:@37408.4]
  assign switch_io_inValid_10 = _T_1208_10; // @[Switch.scala 53:21:@37409.4]
  assign switch_io_inValid_11 = _T_1208_11; // @[Switch.scala 53:21:@37410.4]
  assign switch_io_inValid_12 = _T_1208_12; // @[Switch.scala 53:21:@37411.4]
  assign switch_io_inValid_13 = _T_1208_13; // @[Switch.scala 53:21:@37412.4]
  assign switch_io_inValid_14 = _T_1208_14; // @[Switch.scala 53:21:@37413.4]
  assign switch_io_inValid_15 = _T_1208_15; // @[Switch.scala 53:21:@37414.4]
  assign switch_io_inValid_16 = _T_1208_16; // @[Switch.scala 53:21:@37415.4]
  assign switch_io_inValid_17 = _T_1208_17; // @[Switch.scala 53:21:@37416.4]
  assign switch_io_inValid_18 = _T_1208_18; // @[Switch.scala 53:21:@37417.4]
  assign switch_io_inValid_19 = _T_1208_19; // @[Switch.scala 53:21:@37418.4]
  assign switch_io_inValid_20 = _T_1208_20; // @[Switch.scala 53:21:@37419.4]
  assign switch_io_inValid_21 = _T_1208_21; // @[Switch.scala 53:21:@37420.4]
  assign switch_io_inValid_22 = _T_1208_22; // @[Switch.scala 53:21:@37421.4]
  assign switch_io_inValid_23 = _T_1208_23; // @[Switch.scala 53:21:@37422.4]
  assign switch_io_inValid_24 = _T_1208_24; // @[Switch.scala 53:21:@37423.4]
  assign switch_io_inValid_25 = _T_1208_25; // @[Switch.scala 53:21:@37424.4]
  assign switch_io_inValid_26 = _T_1208_26; // @[Switch.scala 53:21:@37425.4]
  assign switch_io_inValid_27 = _T_1208_27; // @[Switch.scala 53:21:@37426.4]
  assign switch_io_inValid_28 = _T_1208_28; // @[Switch.scala 53:21:@37427.4]
  assign switch_io_inValid_29 = _T_1208_29; // @[Switch.scala 53:21:@37428.4]
  assign switch_io_inValid_30 = _T_1208_30; // @[Switch.scala 53:21:@37429.4]
  assign switch_io_inValid_31 = _T_1208_31; // @[Switch.scala 53:21:@37430.4]
  assign switch_io_inValid_32 = _T_1208_32; // @[Switch.scala 53:21:@37431.4]
  assign switch_io_inValid_33 = _T_1208_33; // @[Switch.scala 53:21:@37432.4]
  assign switch_io_inValid_34 = _T_1208_34; // @[Switch.scala 53:21:@37433.4]
  assign switch_io_inValid_35 = _T_1208_35; // @[Switch.scala 53:21:@37434.4]
  assign switch_io_inValid_36 = _T_1208_36; // @[Switch.scala 53:21:@37435.4]
  assign switch_io_inValid_37 = _T_1208_37; // @[Switch.scala 53:21:@37436.4]
  assign switch_io_inValid_38 = _T_1208_38; // @[Switch.scala 53:21:@37437.4]
  assign switch_io_inValid_39 = _T_1208_39; // @[Switch.scala 53:21:@37438.4]
  assign switch_io_inValid_40 = _T_1208_40; // @[Switch.scala 53:21:@37439.4]
  assign switch_io_inValid_41 = _T_1208_41; // @[Switch.scala 53:21:@37440.4]
  assign switch_io_inValid_42 = _T_1208_42; // @[Switch.scala 53:21:@37441.4]
  assign switch_io_inValid_43 = _T_1208_43; // @[Switch.scala 53:21:@37442.4]
  assign switch_io_inValid_44 = _T_1208_44; // @[Switch.scala 53:21:@37443.4]
  assign switch_io_inValid_45 = _T_1208_45; // @[Switch.scala 53:21:@37444.4]
  assign switch_io_inValid_46 = _T_1208_46; // @[Switch.scala 53:21:@37445.4]
  assign switch_io_inValid_47 = _T_1208_47; // @[Switch.scala 53:21:@37446.4]
  assign switch_io_inValid_48 = _T_1208_48; // @[Switch.scala 53:21:@37447.4]
  assign switch_io_inValid_49 = _T_1208_49; // @[Switch.scala 53:21:@37448.4]
  assign switch_io_inValid_50 = _T_1208_50; // @[Switch.scala 53:21:@37449.4]
  assign switch_io_inValid_51 = _T_1208_51; // @[Switch.scala 53:21:@37450.4]
  assign switch_io_inValid_52 = _T_1208_52; // @[Switch.scala 53:21:@37451.4]
  assign switch_io_inValid_53 = _T_1208_53; // @[Switch.scala 53:21:@37452.4]
  assign switch_io_inValid_54 = _T_1208_54; // @[Switch.scala 53:21:@37453.4]
  assign switch_io_inValid_55 = _T_1208_55; // @[Switch.scala 53:21:@37454.4]
  assign switch_io_inValid_56 = _T_1208_56; // @[Switch.scala 53:21:@37455.4]
  assign switch_io_inValid_57 = _T_1208_57; // @[Switch.scala 53:21:@37456.4]
  assign switch_io_inValid_58 = _T_1208_58; // @[Switch.scala 53:21:@37457.4]
  assign switch_io_inValid_59 = _T_1208_59; // @[Switch.scala 53:21:@37458.4]
  assign switch_io_inValid_60 = _T_1208_60; // @[Switch.scala 53:21:@37459.4]
  assign switch_io_inValid_61 = _T_1208_61; // @[Switch.scala 53:21:@37460.4]
  assign switch_io_inValid_62 = _T_1208_62; // @[Switch.scala 53:21:@37461.4]
  assign switch_io_inValid_63 = _T_1208_63; // @[Switch.scala 53:21:@37462.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_550_0 = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_550_1 = _RAND_1[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_550_2 = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_550_3 = _RAND_3[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_550_4 = _RAND_4[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_550_5 = _RAND_5[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_550_6 = _RAND_6[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_550_7 = _RAND_7[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_550_8 = _RAND_8[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_550_9 = _RAND_9[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_550_10 = _RAND_10[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_550_11 = _RAND_11[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_550_12 = _RAND_12[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_550_13 = _RAND_13[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_550_14 = _RAND_14[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_550_15 = _RAND_15[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_550_16 = _RAND_16[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_550_17 = _RAND_17[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_550_18 = _RAND_18[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_550_19 = _RAND_19[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_550_20 = _RAND_20[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_550_21 = _RAND_21[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_550_22 = _RAND_22[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_550_23 = _RAND_23[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_550_24 = _RAND_24[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_550_25 = _RAND_25[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_550_26 = _RAND_26[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_550_27 = _RAND_27[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_550_28 = _RAND_28[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_550_29 = _RAND_29[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_550_30 = _RAND_30[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_550_31 = _RAND_31[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_550_32 = _RAND_32[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_550_33 = _RAND_33[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_550_34 = _RAND_34[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_550_35 = _RAND_35[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_550_36 = _RAND_36[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_550_37 = _RAND_37[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_550_38 = _RAND_38[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_550_39 = _RAND_39[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_550_40 = _RAND_40[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_550_41 = _RAND_41[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_550_42 = _RAND_42[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_550_43 = _RAND_43[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_550_44 = _RAND_44[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_550_45 = _RAND_45[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_550_46 = _RAND_46[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_550_47 = _RAND_47[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_550_48 = _RAND_48[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_550_49 = _RAND_49[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_550_50 = _RAND_50[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_550_51 = _RAND_51[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_550_52 = _RAND_52[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_550_53 = _RAND_53[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_550_54 = _RAND_54[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_550_55 = _RAND_55[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_550_56 = _RAND_56[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_550_57 = _RAND_57[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_550_58 = _RAND_58[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_550_59 = _RAND_59[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_550_60 = _RAND_60[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_550_61 = _RAND_61[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_550_62 = _RAND_62[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_550_63 = _RAND_63[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {2{`RANDOM}};
  _T_879_0 = _RAND_64[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {2{`RANDOM}};
  _T_879_1 = _RAND_65[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {2{`RANDOM}};
  _T_879_2 = _RAND_66[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {2{`RANDOM}};
  _T_879_3 = _RAND_67[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {2{`RANDOM}};
  _T_879_4 = _RAND_68[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {2{`RANDOM}};
  _T_879_5 = _RAND_69[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {2{`RANDOM}};
  _T_879_6 = _RAND_70[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {2{`RANDOM}};
  _T_879_7 = _RAND_71[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {2{`RANDOM}};
  _T_879_8 = _RAND_72[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {2{`RANDOM}};
  _T_879_9 = _RAND_73[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {2{`RANDOM}};
  _T_879_10 = _RAND_74[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {2{`RANDOM}};
  _T_879_11 = _RAND_75[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {2{`RANDOM}};
  _T_879_12 = _RAND_76[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {2{`RANDOM}};
  _T_879_13 = _RAND_77[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {2{`RANDOM}};
  _T_879_14 = _RAND_78[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {2{`RANDOM}};
  _T_879_15 = _RAND_79[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {2{`RANDOM}};
  _T_879_16 = _RAND_80[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {2{`RANDOM}};
  _T_879_17 = _RAND_81[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {2{`RANDOM}};
  _T_879_18 = _RAND_82[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {2{`RANDOM}};
  _T_879_19 = _RAND_83[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {2{`RANDOM}};
  _T_879_20 = _RAND_84[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {2{`RANDOM}};
  _T_879_21 = _RAND_85[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {2{`RANDOM}};
  _T_879_22 = _RAND_86[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {2{`RANDOM}};
  _T_879_23 = _RAND_87[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {2{`RANDOM}};
  _T_879_24 = _RAND_88[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {2{`RANDOM}};
  _T_879_25 = _RAND_89[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {2{`RANDOM}};
  _T_879_26 = _RAND_90[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {2{`RANDOM}};
  _T_879_27 = _RAND_91[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {2{`RANDOM}};
  _T_879_28 = _RAND_92[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {2{`RANDOM}};
  _T_879_29 = _RAND_93[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {2{`RANDOM}};
  _T_879_30 = _RAND_94[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {2{`RANDOM}};
  _T_879_31 = _RAND_95[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {2{`RANDOM}};
  _T_879_32 = _RAND_96[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {2{`RANDOM}};
  _T_879_33 = _RAND_97[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {2{`RANDOM}};
  _T_879_34 = _RAND_98[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {2{`RANDOM}};
  _T_879_35 = _RAND_99[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {2{`RANDOM}};
  _T_879_36 = _RAND_100[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {2{`RANDOM}};
  _T_879_37 = _RAND_101[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {2{`RANDOM}};
  _T_879_38 = _RAND_102[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {2{`RANDOM}};
  _T_879_39 = _RAND_103[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {2{`RANDOM}};
  _T_879_40 = _RAND_104[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {2{`RANDOM}};
  _T_879_41 = _RAND_105[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {2{`RANDOM}};
  _T_879_42 = _RAND_106[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {2{`RANDOM}};
  _T_879_43 = _RAND_107[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {2{`RANDOM}};
  _T_879_44 = _RAND_108[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {2{`RANDOM}};
  _T_879_45 = _RAND_109[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {2{`RANDOM}};
  _T_879_46 = _RAND_110[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {2{`RANDOM}};
  _T_879_47 = _RAND_111[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {2{`RANDOM}};
  _T_879_48 = _RAND_112[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {2{`RANDOM}};
  _T_879_49 = _RAND_113[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {2{`RANDOM}};
  _T_879_50 = _RAND_114[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {2{`RANDOM}};
  _T_879_51 = _RAND_115[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {2{`RANDOM}};
  _T_879_52 = _RAND_116[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {2{`RANDOM}};
  _T_879_53 = _RAND_117[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {2{`RANDOM}};
  _T_879_54 = _RAND_118[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {2{`RANDOM}};
  _T_879_55 = _RAND_119[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {2{`RANDOM}};
  _T_879_56 = _RAND_120[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {2{`RANDOM}};
  _T_879_57 = _RAND_121[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {2{`RANDOM}};
  _T_879_58 = _RAND_122[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {2{`RANDOM}};
  _T_879_59 = _RAND_123[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {2{`RANDOM}};
  _T_879_60 = _RAND_124[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {2{`RANDOM}};
  _T_879_61 = _RAND_125[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {2{`RANDOM}};
  _T_879_62 = _RAND_126[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {2{`RANDOM}};
  _T_879_63 = _RAND_127[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_1208_0 = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T_1208_1 = _RAND_129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _T_1208_2 = _RAND_130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _T_1208_3 = _RAND_131[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _T_1208_4 = _RAND_132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _T_1208_5 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _T_1208_6 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _T_1208_7 = _RAND_135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _T_1208_8 = _RAND_136[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _T_1208_9 = _RAND_137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _T_1208_10 = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _T_1208_11 = _RAND_139[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _T_1208_12 = _RAND_140[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _T_1208_13 = _RAND_141[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _T_1208_14 = _RAND_142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _T_1208_15 = _RAND_143[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _T_1208_16 = _RAND_144[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _T_1208_17 = _RAND_145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _T_1208_18 = _RAND_146[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  _T_1208_19 = _RAND_147[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  _T_1208_20 = _RAND_148[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  _T_1208_21 = _RAND_149[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _T_1208_22 = _RAND_150[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _T_1208_23 = _RAND_151[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  _T_1208_24 = _RAND_152[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _T_1208_25 = _RAND_153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _T_1208_26 = _RAND_154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _T_1208_27 = _RAND_155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _T_1208_28 = _RAND_156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _T_1208_29 = _RAND_157[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _T_1208_30 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _T_1208_31 = _RAND_159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _T_1208_32 = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _T_1208_33 = _RAND_161[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _T_1208_34 = _RAND_162[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _T_1208_35 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _T_1208_36 = _RAND_164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _T_1208_37 = _RAND_165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _T_1208_38 = _RAND_166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _T_1208_39 = _RAND_167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _T_1208_40 = _RAND_168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _T_1208_41 = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _T_1208_42 = _RAND_170[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _T_1208_43 = _RAND_171[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _T_1208_44 = _RAND_172[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _T_1208_45 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _T_1208_46 = _RAND_174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _T_1208_47 = _RAND_175[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _T_1208_48 = _RAND_176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _T_1208_49 = _RAND_177[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _T_1208_50 = _RAND_178[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _T_1208_51 = _RAND_179[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  _T_1208_52 = _RAND_180[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _T_1208_53 = _RAND_181[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _T_1208_54 = _RAND_182[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _T_1208_55 = _RAND_183[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _T_1208_56 = _RAND_184[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _T_1208_57 = _RAND_185[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _T_1208_58 = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _T_1208_59 = _RAND_187[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _T_1208_60 = _RAND_188[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _T_1208_61 = _RAND_189[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _T_1208_62 = _RAND_190[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  _T_1208_63 = _RAND_191[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  _T_1537_0 = _RAND_192[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  _T_1537_1 = _RAND_193[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _T_1537_2 = _RAND_194[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _T_1537_3 = _RAND_195[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _T_1537_4 = _RAND_196[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  _T_1537_5 = _RAND_197[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  _T_1537_6 = _RAND_198[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  _T_1537_7 = _RAND_199[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _T_1537_8 = _RAND_200[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  _T_1537_9 = _RAND_201[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  _T_1537_10 = _RAND_202[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  _T_1537_11 = _RAND_203[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  _T_1537_12 = _RAND_204[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  _T_1537_13 = _RAND_205[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  _T_1537_14 = _RAND_206[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  _T_1537_15 = _RAND_207[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  _T_1537_16 = _RAND_208[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  _T_1537_17 = _RAND_209[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  _T_1537_18 = _RAND_210[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  _T_1537_19 = _RAND_211[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  _T_1537_20 = _RAND_212[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  _T_1537_21 = _RAND_213[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  _T_1537_22 = _RAND_214[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  _T_1537_23 = _RAND_215[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  _T_1537_24 = _RAND_216[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  _T_1537_25 = _RAND_217[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  _T_1537_26 = _RAND_218[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  _T_1537_27 = _RAND_219[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  _T_1537_28 = _RAND_220[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  _T_1537_29 = _RAND_221[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  _T_1537_30 = _RAND_222[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  _T_1537_31 = _RAND_223[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  _T_1537_32 = _RAND_224[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  _T_1537_33 = _RAND_225[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  _T_1537_34 = _RAND_226[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  _T_1537_35 = _RAND_227[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  _T_1537_36 = _RAND_228[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  _T_1537_37 = _RAND_229[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  _T_1537_38 = _RAND_230[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  _T_1537_39 = _RAND_231[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  _T_1537_40 = _RAND_232[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  _T_1537_41 = _RAND_233[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  _T_1537_42 = _RAND_234[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  _T_1537_43 = _RAND_235[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  _T_1537_44 = _RAND_236[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  _T_1537_45 = _RAND_237[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  _T_1537_46 = _RAND_238[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  _T_1537_47 = _RAND_239[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  _T_1537_48 = _RAND_240[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  _T_1537_49 = _RAND_241[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  _T_1537_50 = _RAND_242[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  _T_1537_51 = _RAND_243[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  _T_1537_52 = _RAND_244[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  _T_1537_53 = _RAND_245[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  _T_1537_54 = _RAND_246[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  _T_1537_55 = _RAND_247[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  _T_1537_56 = _RAND_248[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  _T_1537_57 = _RAND_249[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  _T_1537_58 = _RAND_250[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  _T_1537_59 = _RAND_251[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  _T_1537_60 = _RAND_252[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  _T_1537_61 = _RAND_253[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  _T_1537_62 = _RAND_254[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  _T_1537_63 = _RAND_255[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {2{`RANDOM}};
  _T_1866_0 = _RAND_256[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {2{`RANDOM}};
  _T_1866_1 = _RAND_257[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {2{`RANDOM}};
  _T_1866_2 = _RAND_258[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {2{`RANDOM}};
  _T_1866_3 = _RAND_259[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {2{`RANDOM}};
  _T_1866_4 = _RAND_260[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {2{`RANDOM}};
  _T_1866_5 = _RAND_261[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {2{`RANDOM}};
  _T_1866_6 = _RAND_262[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {2{`RANDOM}};
  _T_1866_7 = _RAND_263[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {2{`RANDOM}};
  _T_1866_8 = _RAND_264[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {2{`RANDOM}};
  _T_1866_9 = _RAND_265[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {2{`RANDOM}};
  _T_1866_10 = _RAND_266[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {2{`RANDOM}};
  _T_1866_11 = _RAND_267[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {2{`RANDOM}};
  _T_1866_12 = _RAND_268[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {2{`RANDOM}};
  _T_1866_13 = _RAND_269[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {2{`RANDOM}};
  _T_1866_14 = _RAND_270[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {2{`RANDOM}};
  _T_1866_15 = _RAND_271[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {2{`RANDOM}};
  _T_1866_16 = _RAND_272[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {2{`RANDOM}};
  _T_1866_17 = _RAND_273[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {2{`RANDOM}};
  _T_1866_18 = _RAND_274[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {2{`RANDOM}};
  _T_1866_19 = _RAND_275[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {2{`RANDOM}};
  _T_1866_20 = _RAND_276[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {2{`RANDOM}};
  _T_1866_21 = _RAND_277[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {2{`RANDOM}};
  _T_1866_22 = _RAND_278[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {2{`RANDOM}};
  _T_1866_23 = _RAND_279[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {2{`RANDOM}};
  _T_1866_24 = _RAND_280[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {2{`RANDOM}};
  _T_1866_25 = _RAND_281[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {2{`RANDOM}};
  _T_1866_26 = _RAND_282[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {2{`RANDOM}};
  _T_1866_27 = _RAND_283[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {2{`RANDOM}};
  _T_1866_28 = _RAND_284[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {2{`RANDOM}};
  _T_1866_29 = _RAND_285[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {2{`RANDOM}};
  _T_1866_30 = _RAND_286[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {2{`RANDOM}};
  _T_1866_31 = _RAND_287[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {2{`RANDOM}};
  _T_1866_32 = _RAND_288[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {2{`RANDOM}};
  _T_1866_33 = _RAND_289[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {2{`RANDOM}};
  _T_1866_34 = _RAND_290[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {2{`RANDOM}};
  _T_1866_35 = _RAND_291[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {2{`RANDOM}};
  _T_1866_36 = _RAND_292[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {2{`RANDOM}};
  _T_1866_37 = _RAND_293[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {2{`RANDOM}};
  _T_1866_38 = _RAND_294[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {2{`RANDOM}};
  _T_1866_39 = _RAND_295[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {2{`RANDOM}};
  _T_1866_40 = _RAND_296[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {2{`RANDOM}};
  _T_1866_41 = _RAND_297[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {2{`RANDOM}};
  _T_1866_42 = _RAND_298[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {2{`RANDOM}};
  _T_1866_43 = _RAND_299[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {2{`RANDOM}};
  _T_1866_44 = _RAND_300[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {2{`RANDOM}};
  _T_1866_45 = _RAND_301[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {2{`RANDOM}};
  _T_1866_46 = _RAND_302[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {2{`RANDOM}};
  _T_1866_47 = _RAND_303[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {2{`RANDOM}};
  _T_1866_48 = _RAND_304[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {2{`RANDOM}};
  _T_1866_49 = _RAND_305[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {2{`RANDOM}};
  _T_1866_50 = _RAND_306[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {2{`RANDOM}};
  _T_1866_51 = _RAND_307[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {2{`RANDOM}};
  _T_1866_52 = _RAND_308[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {2{`RANDOM}};
  _T_1866_53 = _RAND_309[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {2{`RANDOM}};
  _T_1866_54 = _RAND_310[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {2{`RANDOM}};
  _T_1866_55 = _RAND_311[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {2{`RANDOM}};
  _T_1866_56 = _RAND_312[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {2{`RANDOM}};
  _T_1866_57 = _RAND_313[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {2{`RANDOM}};
  _T_1866_58 = _RAND_314[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {2{`RANDOM}};
  _T_1866_59 = _RAND_315[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {2{`RANDOM}};
  _T_1866_60 = _RAND_316[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {2{`RANDOM}};
  _T_1866_61 = _RAND_317[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {2{`RANDOM}};
  _T_1866_62 = _RAND_318[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {2{`RANDOM}};
  _T_1866_63 = _RAND_319[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  _T_2195_0 = _RAND_320[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  _T_2195_1 = _RAND_321[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  _T_2195_2 = _RAND_322[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  _T_2195_3 = _RAND_323[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  _T_2195_4 = _RAND_324[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  _T_2195_5 = _RAND_325[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  _T_2195_6 = _RAND_326[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  _T_2195_7 = _RAND_327[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  _T_2195_8 = _RAND_328[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  _T_2195_9 = _RAND_329[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  _T_2195_10 = _RAND_330[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  _T_2195_11 = _RAND_331[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  _T_2195_12 = _RAND_332[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  _T_2195_13 = _RAND_333[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  _T_2195_14 = _RAND_334[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  _T_2195_15 = _RAND_335[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  _T_2195_16 = _RAND_336[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  _T_2195_17 = _RAND_337[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  _T_2195_18 = _RAND_338[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  _T_2195_19 = _RAND_339[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  _T_2195_20 = _RAND_340[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  _T_2195_21 = _RAND_341[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  _T_2195_22 = _RAND_342[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  _T_2195_23 = _RAND_343[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  _T_2195_24 = _RAND_344[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  _T_2195_25 = _RAND_345[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  _T_2195_26 = _RAND_346[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  _T_2195_27 = _RAND_347[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  _T_2195_28 = _RAND_348[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  _T_2195_29 = _RAND_349[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  _T_2195_30 = _RAND_350[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  _T_2195_31 = _RAND_351[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  _T_2195_32 = _RAND_352[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  _T_2195_33 = _RAND_353[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  _T_2195_34 = _RAND_354[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  _T_2195_35 = _RAND_355[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  _T_2195_36 = _RAND_356[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  _T_2195_37 = _RAND_357[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  _T_2195_38 = _RAND_358[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  _T_2195_39 = _RAND_359[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  _T_2195_40 = _RAND_360[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  _T_2195_41 = _RAND_361[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  _T_2195_42 = _RAND_362[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  _T_2195_43 = _RAND_363[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  _T_2195_44 = _RAND_364[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  _T_2195_45 = _RAND_365[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  _T_2195_46 = _RAND_366[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  _T_2195_47 = _RAND_367[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  _T_2195_48 = _RAND_368[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  _T_2195_49 = _RAND_369[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  _T_2195_50 = _RAND_370[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  _T_2195_51 = _RAND_371[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  _T_2195_52 = _RAND_372[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  _T_2195_53 = _RAND_373[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  _T_2195_54 = _RAND_374[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  _T_2195_55 = _RAND_375[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  _T_2195_56 = _RAND_376[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  _T_2195_57 = _RAND_377[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  _T_2195_58 = _RAND_378[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  _T_2195_59 = _RAND_379[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  _T_2195_60 = _RAND_380[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  _T_2195_61 = _RAND_381[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{`RANDOM}};
  _T_2195_62 = _RAND_382[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{`RANDOM}};
  _T_2195_63 = _RAND_383[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    _T_550_0 <= io_inAddr_0;
    _T_550_1 <= io_inAddr_1;
    _T_550_2 <= io_inAddr_2;
    _T_550_3 <= io_inAddr_3;
    _T_550_4 <= io_inAddr_4;
    _T_550_5 <= io_inAddr_5;
    _T_550_6 <= io_inAddr_6;
    _T_550_7 <= io_inAddr_7;
    _T_550_8 <= io_inAddr_8;
    _T_550_9 <= io_inAddr_9;
    _T_550_10 <= io_inAddr_10;
    _T_550_11 <= io_inAddr_11;
    _T_550_12 <= io_inAddr_12;
    _T_550_13 <= io_inAddr_13;
    _T_550_14 <= io_inAddr_14;
    _T_550_15 <= io_inAddr_15;
    _T_550_16 <= io_inAddr_16;
    _T_550_17 <= io_inAddr_17;
    _T_550_18 <= io_inAddr_18;
    _T_550_19 <= io_inAddr_19;
    _T_550_20 <= io_inAddr_20;
    _T_550_21 <= io_inAddr_21;
    _T_550_22 <= io_inAddr_22;
    _T_550_23 <= io_inAddr_23;
    _T_550_24 <= io_inAddr_24;
    _T_550_25 <= io_inAddr_25;
    _T_550_26 <= io_inAddr_26;
    _T_550_27 <= io_inAddr_27;
    _T_550_28 <= io_inAddr_28;
    _T_550_29 <= io_inAddr_29;
    _T_550_30 <= io_inAddr_30;
    _T_550_31 <= io_inAddr_31;
    _T_550_32 <= io_inAddr_32;
    _T_550_33 <= io_inAddr_33;
    _T_550_34 <= io_inAddr_34;
    _T_550_35 <= io_inAddr_35;
    _T_550_36 <= io_inAddr_36;
    _T_550_37 <= io_inAddr_37;
    _T_550_38 <= io_inAddr_38;
    _T_550_39 <= io_inAddr_39;
    _T_550_40 <= io_inAddr_40;
    _T_550_41 <= io_inAddr_41;
    _T_550_42 <= io_inAddr_42;
    _T_550_43 <= io_inAddr_43;
    _T_550_44 <= io_inAddr_44;
    _T_550_45 <= io_inAddr_45;
    _T_550_46 <= io_inAddr_46;
    _T_550_47 <= io_inAddr_47;
    _T_550_48 <= io_inAddr_48;
    _T_550_49 <= io_inAddr_49;
    _T_550_50 <= io_inAddr_50;
    _T_550_51 <= io_inAddr_51;
    _T_550_52 <= io_inAddr_52;
    _T_550_53 <= io_inAddr_53;
    _T_550_54 <= io_inAddr_54;
    _T_550_55 <= io_inAddr_55;
    _T_550_56 <= io_inAddr_56;
    _T_550_57 <= io_inAddr_57;
    _T_550_58 <= io_inAddr_58;
    _T_550_59 <= io_inAddr_59;
    _T_550_60 <= io_inAddr_60;
    _T_550_61 <= io_inAddr_61;
    _T_550_62 <= io_inAddr_62;
    _T_550_63 <= io_inAddr_63;
    _T_879_0 <= io_inData_0;
    _T_879_1 <= io_inData_1;
    _T_879_2 <= io_inData_2;
    _T_879_3 <= io_inData_3;
    _T_879_4 <= io_inData_4;
    _T_879_5 <= io_inData_5;
    _T_879_6 <= io_inData_6;
    _T_879_7 <= io_inData_7;
    _T_879_8 <= io_inData_8;
    _T_879_9 <= io_inData_9;
    _T_879_10 <= io_inData_10;
    _T_879_11 <= io_inData_11;
    _T_879_12 <= io_inData_12;
    _T_879_13 <= io_inData_13;
    _T_879_14 <= io_inData_14;
    _T_879_15 <= io_inData_15;
    _T_879_16 <= io_inData_16;
    _T_879_17 <= io_inData_17;
    _T_879_18 <= io_inData_18;
    _T_879_19 <= io_inData_19;
    _T_879_20 <= io_inData_20;
    _T_879_21 <= io_inData_21;
    _T_879_22 <= io_inData_22;
    _T_879_23 <= io_inData_23;
    _T_879_24 <= io_inData_24;
    _T_879_25 <= io_inData_25;
    _T_879_26 <= io_inData_26;
    _T_879_27 <= io_inData_27;
    _T_879_28 <= io_inData_28;
    _T_879_29 <= io_inData_29;
    _T_879_30 <= io_inData_30;
    _T_879_31 <= io_inData_31;
    _T_879_32 <= io_inData_32;
    _T_879_33 <= io_inData_33;
    _T_879_34 <= io_inData_34;
    _T_879_35 <= io_inData_35;
    _T_879_36 <= io_inData_36;
    _T_879_37 <= io_inData_37;
    _T_879_38 <= io_inData_38;
    _T_879_39 <= io_inData_39;
    _T_879_40 <= io_inData_40;
    _T_879_41 <= io_inData_41;
    _T_879_42 <= io_inData_42;
    _T_879_43 <= io_inData_43;
    _T_879_44 <= io_inData_44;
    _T_879_45 <= io_inData_45;
    _T_879_46 <= io_inData_46;
    _T_879_47 <= io_inData_47;
    _T_879_48 <= io_inData_48;
    _T_879_49 <= io_inData_49;
    _T_879_50 <= io_inData_50;
    _T_879_51 <= io_inData_51;
    _T_879_52 <= io_inData_52;
    _T_879_53 <= io_inData_53;
    _T_879_54 <= io_inData_54;
    _T_879_55 <= io_inData_55;
    _T_879_56 <= io_inData_56;
    _T_879_57 <= io_inData_57;
    _T_879_58 <= io_inData_58;
    _T_879_59 <= io_inData_59;
    _T_879_60 <= io_inData_60;
    _T_879_61 <= io_inData_61;
    _T_879_62 <= io_inData_62;
    _T_879_63 <= io_inData_63;
    _T_1208_0 <= io_inValid_0;
    _T_1208_1 <= io_inValid_1;
    _T_1208_2 <= io_inValid_2;
    _T_1208_3 <= io_inValid_3;
    _T_1208_4 <= io_inValid_4;
    _T_1208_5 <= io_inValid_5;
    _T_1208_6 <= io_inValid_6;
    _T_1208_7 <= io_inValid_7;
    _T_1208_8 <= io_inValid_8;
    _T_1208_9 <= io_inValid_9;
    _T_1208_10 <= io_inValid_10;
    _T_1208_11 <= io_inValid_11;
    _T_1208_12 <= io_inValid_12;
    _T_1208_13 <= io_inValid_13;
    _T_1208_14 <= io_inValid_14;
    _T_1208_15 <= io_inValid_15;
    _T_1208_16 <= io_inValid_16;
    _T_1208_17 <= io_inValid_17;
    _T_1208_18 <= io_inValid_18;
    _T_1208_19 <= io_inValid_19;
    _T_1208_20 <= io_inValid_20;
    _T_1208_21 <= io_inValid_21;
    _T_1208_22 <= io_inValid_22;
    _T_1208_23 <= io_inValid_23;
    _T_1208_24 <= io_inValid_24;
    _T_1208_25 <= io_inValid_25;
    _T_1208_26 <= io_inValid_26;
    _T_1208_27 <= io_inValid_27;
    _T_1208_28 <= io_inValid_28;
    _T_1208_29 <= io_inValid_29;
    _T_1208_30 <= io_inValid_30;
    _T_1208_31 <= io_inValid_31;
    _T_1208_32 <= io_inValid_32;
    _T_1208_33 <= io_inValid_33;
    _T_1208_34 <= io_inValid_34;
    _T_1208_35 <= io_inValid_35;
    _T_1208_36 <= io_inValid_36;
    _T_1208_37 <= io_inValid_37;
    _T_1208_38 <= io_inValid_38;
    _T_1208_39 <= io_inValid_39;
    _T_1208_40 <= io_inValid_40;
    _T_1208_41 <= io_inValid_41;
    _T_1208_42 <= io_inValid_42;
    _T_1208_43 <= io_inValid_43;
    _T_1208_44 <= io_inValid_44;
    _T_1208_45 <= io_inValid_45;
    _T_1208_46 <= io_inValid_46;
    _T_1208_47 <= io_inValid_47;
    _T_1208_48 <= io_inValid_48;
    _T_1208_49 <= io_inValid_49;
    _T_1208_50 <= io_inValid_50;
    _T_1208_51 <= io_inValid_51;
    _T_1208_52 <= io_inValid_52;
    _T_1208_53 <= io_inValid_53;
    _T_1208_54 <= io_inValid_54;
    _T_1208_55 <= io_inValid_55;
    _T_1208_56 <= io_inValid_56;
    _T_1208_57 <= io_inValid_57;
    _T_1208_58 <= io_inValid_58;
    _T_1208_59 <= io_inValid_59;
    _T_1208_60 <= io_inValid_60;
    _T_1208_61 <= io_inValid_61;
    _T_1208_62 <= io_inValid_62;
    _T_1208_63 <= io_inValid_63;
    _T_1537_0 <= switch_io_outAck_0;
    _T_1537_1 <= switch_io_outAck_1;
    _T_1537_2 <= switch_io_outAck_2;
    _T_1537_3 <= switch_io_outAck_3;
    _T_1537_4 <= switch_io_outAck_4;
    _T_1537_5 <= switch_io_outAck_5;
    _T_1537_6 <= switch_io_outAck_6;
    _T_1537_7 <= switch_io_outAck_7;
    _T_1537_8 <= switch_io_outAck_8;
    _T_1537_9 <= switch_io_outAck_9;
    _T_1537_10 <= switch_io_outAck_10;
    _T_1537_11 <= switch_io_outAck_11;
    _T_1537_12 <= switch_io_outAck_12;
    _T_1537_13 <= switch_io_outAck_13;
    _T_1537_14 <= switch_io_outAck_14;
    _T_1537_15 <= switch_io_outAck_15;
    _T_1537_16 <= switch_io_outAck_16;
    _T_1537_17 <= switch_io_outAck_17;
    _T_1537_18 <= switch_io_outAck_18;
    _T_1537_19 <= switch_io_outAck_19;
    _T_1537_20 <= switch_io_outAck_20;
    _T_1537_21 <= switch_io_outAck_21;
    _T_1537_22 <= switch_io_outAck_22;
    _T_1537_23 <= switch_io_outAck_23;
    _T_1537_24 <= switch_io_outAck_24;
    _T_1537_25 <= switch_io_outAck_25;
    _T_1537_26 <= switch_io_outAck_26;
    _T_1537_27 <= switch_io_outAck_27;
    _T_1537_28 <= switch_io_outAck_28;
    _T_1537_29 <= switch_io_outAck_29;
    _T_1537_30 <= switch_io_outAck_30;
    _T_1537_31 <= switch_io_outAck_31;
    _T_1537_32 <= switch_io_outAck_32;
    _T_1537_33 <= switch_io_outAck_33;
    _T_1537_34 <= switch_io_outAck_34;
    _T_1537_35 <= switch_io_outAck_35;
    _T_1537_36 <= switch_io_outAck_36;
    _T_1537_37 <= switch_io_outAck_37;
    _T_1537_38 <= switch_io_outAck_38;
    _T_1537_39 <= switch_io_outAck_39;
    _T_1537_40 <= switch_io_outAck_40;
    _T_1537_41 <= switch_io_outAck_41;
    _T_1537_42 <= switch_io_outAck_42;
    _T_1537_43 <= switch_io_outAck_43;
    _T_1537_44 <= switch_io_outAck_44;
    _T_1537_45 <= switch_io_outAck_45;
    _T_1537_46 <= switch_io_outAck_46;
    _T_1537_47 <= switch_io_outAck_47;
    _T_1537_48 <= switch_io_outAck_48;
    _T_1537_49 <= switch_io_outAck_49;
    _T_1537_50 <= switch_io_outAck_50;
    _T_1537_51 <= switch_io_outAck_51;
    _T_1537_52 <= switch_io_outAck_52;
    _T_1537_53 <= switch_io_outAck_53;
    _T_1537_54 <= switch_io_outAck_54;
    _T_1537_55 <= switch_io_outAck_55;
    _T_1537_56 <= switch_io_outAck_56;
    _T_1537_57 <= switch_io_outAck_57;
    _T_1537_58 <= switch_io_outAck_58;
    _T_1537_59 <= switch_io_outAck_59;
    _T_1537_60 <= switch_io_outAck_60;
    _T_1537_61 <= switch_io_outAck_61;
    _T_1537_62 <= switch_io_outAck_62;
    _T_1537_63 <= switch_io_outAck_63;
    _T_1866_0 <= switch_io_outData_0;
    _T_1866_1 <= switch_io_outData_1;
    _T_1866_2 <= switch_io_outData_2;
    _T_1866_3 <= switch_io_outData_3;
    _T_1866_4 <= switch_io_outData_4;
    _T_1866_5 <= switch_io_outData_5;
    _T_1866_6 <= switch_io_outData_6;
    _T_1866_7 <= switch_io_outData_7;
    _T_1866_8 <= switch_io_outData_8;
    _T_1866_9 <= switch_io_outData_9;
    _T_1866_10 <= switch_io_outData_10;
    _T_1866_11 <= switch_io_outData_11;
    _T_1866_12 <= switch_io_outData_12;
    _T_1866_13 <= switch_io_outData_13;
    _T_1866_14 <= switch_io_outData_14;
    _T_1866_15 <= switch_io_outData_15;
    _T_1866_16 <= switch_io_outData_16;
    _T_1866_17 <= switch_io_outData_17;
    _T_1866_18 <= switch_io_outData_18;
    _T_1866_19 <= switch_io_outData_19;
    _T_1866_20 <= switch_io_outData_20;
    _T_1866_21 <= switch_io_outData_21;
    _T_1866_22 <= switch_io_outData_22;
    _T_1866_23 <= switch_io_outData_23;
    _T_1866_24 <= switch_io_outData_24;
    _T_1866_25 <= switch_io_outData_25;
    _T_1866_26 <= switch_io_outData_26;
    _T_1866_27 <= switch_io_outData_27;
    _T_1866_28 <= switch_io_outData_28;
    _T_1866_29 <= switch_io_outData_29;
    _T_1866_30 <= switch_io_outData_30;
    _T_1866_31 <= switch_io_outData_31;
    _T_1866_32 <= switch_io_outData_32;
    _T_1866_33 <= switch_io_outData_33;
    _T_1866_34 <= switch_io_outData_34;
    _T_1866_35 <= switch_io_outData_35;
    _T_1866_36 <= switch_io_outData_36;
    _T_1866_37 <= switch_io_outData_37;
    _T_1866_38 <= switch_io_outData_38;
    _T_1866_39 <= switch_io_outData_39;
    _T_1866_40 <= switch_io_outData_40;
    _T_1866_41 <= switch_io_outData_41;
    _T_1866_42 <= switch_io_outData_42;
    _T_1866_43 <= switch_io_outData_43;
    _T_1866_44 <= switch_io_outData_44;
    _T_1866_45 <= switch_io_outData_45;
    _T_1866_46 <= switch_io_outData_46;
    _T_1866_47 <= switch_io_outData_47;
    _T_1866_48 <= switch_io_outData_48;
    _T_1866_49 <= switch_io_outData_49;
    _T_1866_50 <= switch_io_outData_50;
    _T_1866_51 <= switch_io_outData_51;
    _T_1866_52 <= switch_io_outData_52;
    _T_1866_53 <= switch_io_outData_53;
    _T_1866_54 <= switch_io_outData_54;
    _T_1866_55 <= switch_io_outData_55;
    _T_1866_56 <= switch_io_outData_56;
    _T_1866_57 <= switch_io_outData_57;
    _T_1866_58 <= switch_io_outData_58;
    _T_1866_59 <= switch_io_outData_59;
    _T_1866_60 <= switch_io_outData_60;
    _T_1866_61 <= switch_io_outData_61;
    _T_1866_62 <= switch_io_outData_62;
    _T_1866_63 <= switch_io_outData_63;
    _T_2195_0 <= switch_io_outValid_0;
    _T_2195_1 <= switch_io_outValid_1;
    _T_2195_2 <= switch_io_outValid_2;
    _T_2195_3 <= switch_io_outValid_3;
    _T_2195_4 <= switch_io_outValid_4;
    _T_2195_5 <= switch_io_outValid_5;
    _T_2195_6 <= switch_io_outValid_6;
    _T_2195_7 <= switch_io_outValid_7;
    _T_2195_8 <= switch_io_outValid_8;
    _T_2195_9 <= switch_io_outValid_9;
    _T_2195_10 <= switch_io_outValid_10;
    _T_2195_11 <= switch_io_outValid_11;
    _T_2195_12 <= switch_io_outValid_12;
    _T_2195_13 <= switch_io_outValid_13;
    _T_2195_14 <= switch_io_outValid_14;
    _T_2195_15 <= switch_io_outValid_15;
    _T_2195_16 <= switch_io_outValid_16;
    _T_2195_17 <= switch_io_outValid_17;
    _T_2195_18 <= switch_io_outValid_18;
    _T_2195_19 <= switch_io_outValid_19;
    _T_2195_20 <= switch_io_outValid_20;
    _T_2195_21 <= switch_io_outValid_21;
    _T_2195_22 <= switch_io_outValid_22;
    _T_2195_23 <= switch_io_outValid_23;
    _T_2195_24 <= switch_io_outValid_24;
    _T_2195_25 <= switch_io_outValid_25;
    _T_2195_26 <= switch_io_outValid_26;
    _T_2195_27 <= switch_io_outValid_27;
    _T_2195_28 <= switch_io_outValid_28;
    _T_2195_29 <= switch_io_outValid_29;
    _T_2195_30 <= switch_io_outValid_30;
    _T_2195_31 <= switch_io_outValid_31;
    _T_2195_32 <= switch_io_outValid_32;
    _T_2195_33 <= switch_io_outValid_33;
    _T_2195_34 <= switch_io_outValid_34;
    _T_2195_35 <= switch_io_outValid_35;
    _T_2195_36 <= switch_io_outValid_36;
    _T_2195_37 <= switch_io_outValid_37;
    _T_2195_38 <= switch_io_outValid_38;
    _T_2195_39 <= switch_io_outValid_39;
    _T_2195_40 <= switch_io_outValid_40;
    _T_2195_41 <= switch_io_outValid_41;
    _T_2195_42 <= switch_io_outValid_42;
    _T_2195_43 <= switch_io_outValid_43;
    _T_2195_44 <= switch_io_outValid_44;
    _T_2195_45 <= switch_io_outValid_45;
    _T_2195_46 <= switch_io_outValid_46;
    _T_2195_47 <= switch_io_outValid_47;
    _T_2195_48 <= switch_io_outValid_48;
    _T_2195_49 <= switch_io_outValid_49;
    _T_2195_50 <= switch_io_outValid_50;
    _T_2195_51 <= switch_io_outValid_51;
    _T_2195_52 <= switch_io_outValid_52;
    _T_2195_53 <= switch_io_outValid_53;
    _T_2195_54 <= switch_io_outValid_54;
    _T_2195_55 <= switch_io_outValid_55;
    _T_2195_56 <= switch_io_outValid_56;
    _T_2195_57 <= switch_io_outValid_57;
    _T_2195_58 <= switch_io_outValid_58;
    _T_2195_59 <= switch_io_outValid_59;
    _T_2195_60 <= switch_io_outValid_60;
    _T_2195_61 <= switch_io_outValid_61;
    _T_2195_62 <= switch_io_outValid_62;
    _T_2195_63 <= switch_io_outValid_63;
  end
endmodule
