module Switch( // @[:@3.2]
  input  [2:0]  io_inAddr_0, // @[:@6.4]
  input  [2:0]  io_inAddr_1, // @[:@6.4]
  input  [2:0]  io_inAddr_2, // @[:@6.4]
  input  [2:0]  io_inAddr_3, // @[:@6.4]
  input  [2:0]  io_inAddr_4, // @[:@6.4]
  input  [2:0]  io_inAddr_5, // @[:@6.4]
  input  [2:0]  io_inAddr_6, // @[:@6.4]
  input  [2:0]  io_inAddr_7, // @[:@6.4]
  input  [47:0] io_inData_0, // @[:@6.4]
  input  [47:0] io_inData_1, // @[:@6.4]
  input  [47:0] io_inData_2, // @[:@6.4]
  input  [47:0] io_inData_3, // @[:@6.4]
  input  [47:0] io_inData_4, // @[:@6.4]
  input  [47:0] io_inData_5, // @[:@6.4]
  input  [47:0] io_inData_6, // @[:@6.4]
  input  [47:0] io_inData_7, // @[:@6.4]
  input         io_inValid_0, // @[:@6.4]
  input         io_inValid_1, // @[:@6.4]
  input         io_inValid_2, // @[:@6.4]
  input         io_inValid_3, // @[:@6.4]
  input         io_inValid_4, // @[:@6.4]
  input         io_inValid_5, // @[:@6.4]
  input         io_inValid_6, // @[:@6.4]
  input         io_inValid_7, // @[:@6.4]
  output        io_outAck_0, // @[:@6.4]
  output        io_outAck_1, // @[:@6.4]
  output        io_outAck_2, // @[:@6.4]
  output        io_outAck_3, // @[:@6.4]
  output        io_outAck_4, // @[:@6.4]
  output        io_outAck_5, // @[:@6.4]
  output        io_outAck_6, // @[:@6.4]
  output        io_outAck_7, // @[:@6.4]
  output [47:0] io_outData_0, // @[:@6.4]
  output [47:0] io_outData_1, // @[:@6.4]
  output [47:0] io_outData_2, // @[:@6.4]
  output [47:0] io_outData_3, // @[:@6.4]
  output [47:0] io_outData_4, // @[:@6.4]
  output [47:0] io_outData_5, // @[:@6.4]
  output [47:0] io_outData_6, // @[:@6.4]
  output [47:0] io_outData_7, // @[:@6.4]
  output        io_outValid_0, // @[:@6.4]
  output        io_outValid_1, // @[:@6.4]
  output        io_outValid_2, // @[:@6.4]
  output        io_outValid_3, // @[:@6.4]
  output        io_outValid_4, // @[:@6.4]
  output        io_outValid_5, // @[:@6.4]
  output        io_outValid_6, // @[:@6.4]
  output        io_outValid_7 // @[:@6.4]
);
  wire  _T_462; // @[Switch.scala 30:53:@10.4]
  wire  valid_0_0; // @[Switch.scala 30:36:@11.4]
  wire  _T_465; // @[Switch.scala 30:53:@13.4]
  wire  valid_0_1; // @[Switch.scala 30:36:@14.4]
  wire  _T_468; // @[Switch.scala 30:53:@16.4]
  wire  valid_0_2; // @[Switch.scala 30:36:@17.4]
  wire  _T_471; // @[Switch.scala 30:53:@19.4]
  wire  valid_0_3; // @[Switch.scala 30:36:@20.4]
  wire  _T_474; // @[Switch.scala 30:53:@22.4]
  wire  valid_0_4; // @[Switch.scala 30:36:@23.4]
  wire  _T_477; // @[Switch.scala 30:53:@25.4]
  wire  valid_0_5; // @[Switch.scala 30:36:@26.4]
  wire  _T_480; // @[Switch.scala 30:53:@28.4]
  wire  valid_0_6; // @[Switch.scala 30:36:@29.4]
  wire  _T_483; // @[Switch.scala 30:53:@31.4]
  wire  valid_0_7; // @[Switch.scala 30:36:@32.4]
  wire [2:0] _T_493; // @[Mux.scala 31:69:@34.4]
  wire [2:0] _T_494; // @[Mux.scala 31:69:@35.4]
  wire [2:0] _T_495; // @[Mux.scala 31:69:@36.4]
  wire [2:0] _T_496; // @[Mux.scala 31:69:@37.4]
  wire [2:0] _T_497; // @[Mux.scala 31:69:@38.4]
  wire [2:0] _T_498; // @[Mux.scala 31:69:@39.4]
  wire [2:0] select_0; // @[Mux.scala 31:69:@40.4]
  wire [47:0] _GEN_1; // @[Switch.scala 33:19:@42.4]
  wire [47:0] _GEN_2; // @[Switch.scala 33:19:@42.4]
  wire [47:0] _GEN_3; // @[Switch.scala 33:19:@42.4]
  wire [47:0] _GEN_4; // @[Switch.scala 33:19:@42.4]
  wire [47:0] _GEN_5; // @[Switch.scala 33:19:@42.4]
  wire [47:0] _GEN_6; // @[Switch.scala 33:19:@42.4]
  wire [7:0] _T_507; // @[Switch.scala 34:32:@49.4]
  wire  _T_511; // @[Switch.scala 30:53:@52.4]
  wire  valid_1_0; // @[Switch.scala 30:36:@53.4]
  wire  _T_514; // @[Switch.scala 30:53:@55.4]
  wire  valid_1_1; // @[Switch.scala 30:36:@56.4]
  wire  _T_517; // @[Switch.scala 30:53:@58.4]
  wire  valid_1_2; // @[Switch.scala 30:36:@59.4]
  wire  _T_520; // @[Switch.scala 30:53:@61.4]
  wire  valid_1_3; // @[Switch.scala 30:36:@62.4]
  wire  _T_523; // @[Switch.scala 30:53:@64.4]
  wire  valid_1_4; // @[Switch.scala 30:36:@65.4]
  wire  _T_526; // @[Switch.scala 30:53:@67.4]
  wire  valid_1_5; // @[Switch.scala 30:36:@68.4]
  wire  _T_529; // @[Switch.scala 30:53:@70.4]
  wire  valid_1_6; // @[Switch.scala 30:36:@71.4]
  wire  _T_532; // @[Switch.scala 30:53:@73.4]
  wire  valid_1_7; // @[Switch.scala 30:36:@74.4]
  wire [2:0] _T_542; // @[Mux.scala 31:69:@76.4]
  wire [2:0] _T_543; // @[Mux.scala 31:69:@77.4]
  wire [2:0] _T_544; // @[Mux.scala 31:69:@78.4]
  wire [2:0] _T_545; // @[Mux.scala 31:69:@79.4]
  wire [2:0] _T_546; // @[Mux.scala 31:69:@80.4]
  wire [2:0] _T_547; // @[Mux.scala 31:69:@81.4]
  wire [2:0] select_1; // @[Mux.scala 31:69:@82.4]
  wire [47:0] _GEN_9; // @[Switch.scala 33:19:@84.4]
  wire [47:0] _GEN_10; // @[Switch.scala 33:19:@84.4]
  wire [47:0] _GEN_11; // @[Switch.scala 33:19:@84.4]
  wire [47:0] _GEN_12; // @[Switch.scala 33:19:@84.4]
  wire [47:0] _GEN_13; // @[Switch.scala 33:19:@84.4]
  wire [47:0] _GEN_14; // @[Switch.scala 33:19:@84.4]
  wire [7:0] _T_556; // @[Switch.scala 34:32:@91.4]
  wire  _T_560; // @[Switch.scala 30:53:@94.4]
  wire  valid_2_0; // @[Switch.scala 30:36:@95.4]
  wire  _T_563; // @[Switch.scala 30:53:@97.4]
  wire  valid_2_1; // @[Switch.scala 30:36:@98.4]
  wire  _T_566; // @[Switch.scala 30:53:@100.4]
  wire  valid_2_2; // @[Switch.scala 30:36:@101.4]
  wire  _T_569; // @[Switch.scala 30:53:@103.4]
  wire  valid_2_3; // @[Switch.scala 30:36:@104.4]
  wire  _T_572; // @[Switch.scala 30:53:@106.4]
  wire  valid_2_4; // @[Switch.scala 30:36:@107.4]
  wire  _T_575; // @[Switch.scala 30:53:@109.4]
  wire  valid_2_5; // @[Switch.scala 30:36:@110.4]
  wire  _T_578; // @[Switch.scala 30:53:@112.4]
  wire  valid_2_6; // @[Switch.scala 30:36:@113.4]
  wire  _T_581; // @[Switch.scala 30:53:@115.4]
  wire  valid_2_7; // @[Switch.scala 30:36:@116.4]
  wire [2:0] _T_591; // @[Mux.scala 31:69:@118.4]
  wire [2:0] _T_592; // @[Mux.scala 31:69:@119.4]
  wire [2:0] _T_593; // @[Mux.scala 31:69:@120.4]
  wire [2:0] _T_594; // @[Mux.scala 31:69:@121.4]
  wire [2:0] _T_595; // @[Mux.scala 31:69:@122.4]
  wire [2:0] _T_596; // @[Mux.scala 31:69:@123.4]
  wire [2:0] select_2; // @[Mux.scala 31:69:@124.4]
  wire [47:0] _GEN_17; // @[Switch.scala 33:19:@126.4]
  wire [47:0] _GEN_18; // @[Switch.scala 33:19:@126.4]
  wire [47:0] _GEN_19; // @[Switch.scala 33:19:@126.4]
  wire [47:0] _GEN_20; // @[Switch.scala 33:19:@126.4]
  wire [47:0] _GEN_21; // @[Switch.scala 33:19:@126.4]
  wire [47:0] _GEN_22; // @[Switch.scala 33:19:@126.4]
  wire [7:0] _T_605; // @[Switch.scala 34:32:@133.4]
  wire  _T_609; // @[Switch.scala 30:53:@136.4]
  wire  valid_3_0; // @[Switch.scala 30:36:@137.4]
  wire  _T_612; // @[Switch.scala 30:53:@139.4]
  wire  valid_3_1; // @[Switch.scala 30:36:@140.4]
  wire  _T_615; // @[Switch.scala 30:53:@142.4]
  wire  valid_3_2; // @[Switch.scala 30:36:@143.4]
  wire  _T_618; // @[Switch.scala 30:53:@145.4]
  wire  valid_3_3; // @[Switch.scala 30:36:@146.4]
  wire  _T_621; // @[Switch.scala 30:53:@148.4]
  wire  valid_3_4; // @[Switch.scala 30:36:@149.4]
  wire  _T_624; // @[Switch.scala 30:53:@151.4]
  wire  valid_3_5; // @[Switch.scala 30:36:@152.4]
  wire  _T_627; // @[Switch.scala 30:53:@154.4]
  wire  valid_3_6; // @[Switch.scala 30:36:@155.4]
  wire  _T_630; // @[Switch.scala 30:53:@157.4]
  wire  valid_3_7; // @[Switch.scala 30:36:@158.4]
  wire [2:0] _T_640; // @[Mux.scala 31:69:@160.4]
  wire [2:0] _T_641; // @[Mux.scala 31:69:@161.4]
  wire [2:0] _T_642; // @[Mux.scala 31:69:@162.4]
  wire [2:0] _T_643; // @[Mux.scala 31:69:@163.4]
  wire [2:0] _T_644; // @[Mux.scala 31:69:@164.4]
  wire [2:0] _T_645; // @[Mux.scala 31:69:@165.4]
  wire [2:0] select_3; // @[Mux.scala 31:69:@166.4]
  wire [47:0] _GEN_25; // @[Switch.scala 33:19:@168.4]
  wire [47:0] _GEN_26; // @[Switch.scala 33:19:@168.4]
  wire [47:0] _GEN_27; // @[Switch.scala 33:19:@168.4]
  wire [47:0] _GEN_28; // @[Switch.scala 33:19:@168.4]
  wire [47:0] _GEN_29; // @[Switch.scala 33:19:@168.4]
  wire [47:0] _GEN_30; // @[Switch.scala 33:19:@168.4]
  wire [7:0] _T_654; // @[Switch.scala 34:32:@175.4]
  wire  _T_658; // @[Switch.scala 30:53:@178.4]
  wire  valid_4_0; // @[Switch.scala 30:36:@179.4]
  wire  _T_661; // @[Switch.scala 30:53:@181.4]
  wire  valid_4_1; // @[Switch.scala 30:36:@182.4]
  wire  _T_664; // @[Switch.scala 30:53:@184.4]
  wire  valid_4_2; // @[Switch.scala 30:36:@185.4]
  wire  _T_667; // @[Switch.scala 30:53:@187.4]
  wire  valid_4_3; // @[Switch.scala 30:36:@188.4]
  wire  _T_670; // @[Switch.scala 30:53:@190.4]
  wire  valid_4_4; // @[Switch.scala 30:36:@191.4]
  wire  _T_673; // @[Switch.scala 30:53:@193.4]
  wire  valid_4_5; // @[Switch.scala 30:36:@194.4]
  wire  _T_676; // @[Switch.scala 30:53:@196.4]
  wire  valid_4_6; // @[Switch.scala 30:36:@197.4]
  wire  _T_679; // @[Switch.scala 30:53:@199.4]
  wire  valid_4_7; // @[Switch.scala 30:36:@200.4]
  wire [2:0] _T_689; // @[Mux.scala 31:69:@202.4]
  wire [2:0] _T_690; // @[Mux.scala 31:69:@203.4]
  wire [2:0] _T_691; // @[Mux.scala 31:69:@204.4]
  wire [2:0] _T_692; // @[Mux.scala 31:69:@205.4]
  wire [2:0] _T_693; // @[Mux.scala 31:69:@206.4]
  wire [2:0] _T_694; // @[Mux.scala 31:69:@207.4]
  wire [2:0] select_4; // @[Mux.scala 31:69:@208.4]
  wire [47:0] _GEN_33; // @[Switch.scala 33:19:@210.4]
  wire [47:0] _GEN_34; // @[Switch.scala 33:19:@210.4]
  wire [47:0] _GEN_35; // @[Switch.scala 33:19:@210.4]
  wire [47:0] _GEN_36; // @[Switch.scala 33:19:@210.4]
  wire [47:0] _GEN_37; // @[Switch.scala 33:19:@210.4]
  wire [47:0] _GEN_38; // @[Switch.scala 33:19:@210.4]
  wire [7:0] _T_703; // @[Switch.scala 34:32:@217.4]
  wire  _T_707; // @[Switch.scala 30:53:@220.4]
  wire  valid_5_0; // @[Switch.scala 30:36:@221.4]
  wire  _T_710; // @[Switch.scala 30:53:@223.4]
  wire  valid_5_1; // @[Switch.scala 30:36:@224.4]
  wire  _T_713; // @[Switch.scala 30:53:@226.4]
  wire  valid_5_2; // @[Switch.scala 30:36:@227.4]
  wire  _T_716; // @[Switch.scala 30:53:@229.4]
  wire  valid_5_3; // @[Switch.scala 30:36:@230.4]
  wire  _T_719; // @[Switch.scala 30:53:@232.4]
  wire  valid_5_4; // @[Switch.scala 30:36:@233.4]
  wire  _T_722; // @[Switch.scala 30:53:@235.4]
  wire  valid_5_5; // @[Switch.scala 30:36:@236.4]
  wire  _T_725; // @[Switch.scala 30:53:@238.4]
  wire  valid_5_6; // @[Switch.scala 30:36:@239.4]
  wire  _T_728; // @[Switch.scala 30:53:@241.4]
  wire  valid_5_7; // @[Switch.scala 30:36:@242.4]
  wire [2:0] _T_738; // @[Mux.scala 31:69:@244.4]
  wire [2:0] _T_739; // @[Mux.scala 31:69:@245.4]
  wire [2:0] _T_740; // @[Mux.scala 31:69:@246.4]
  wire [2:0] _T_741; // @[Mux.scala 31:69:@247.4]
  wire [2:0] _T_742; // @[Mux.scala 31:69:@248.4]
  wire [2:0] _T_743; // @[Mux.scala 31:69:@249.4]
  wire [2:0] select_5; // @[Mux.scala 31:69:@250.4]
  wire [47:0] _GEN_41; // @[Switch.scala 33:19:@252.4]
  wire [47:0] _GEN_42; // @[Switch.scala 33:19:@252.4]
  wire [47:0] _GEN_43; // @[Switch.scala 33:19:@252.4]
  wire [47:0] _GEN_44; // @[Switch.scala 33:19:@252.4]
  wire [47:0] _GEN_45; // @[Switch.scala 33:19:@252.4]
  wire [47:0] _GEN_46; // @[Switch.scala 33:19:@252.4]
  wire [7:0] _T_752; // @[Switch.scala 34:32:@259.4]
  wire  _T_756; // @[Switch.scala 30:53:@262.4]
  wire  valid_6_0; // @[Switch.scala 30:36:@263.4]
  wire  _T_759; // @[Switch.scala 30:53:@265.4]
  wire  valid_6_1; // @[Switch.scala 30:36:@266.4]
  wire  _T_762; // @[Switch.scala 30:53:@268.4]
  wire  valid_6_2; // @[Switch.scala 30:36:@269.4]
  wire  _T_765; // @[Switch.scala 30:53:@271.4]
  wire  valid_6_3; // @[Switch.scala 30:36:@272.4]
  wire  _T_768; // @[Switch.scala 30:53:@274.4]
  wire  valid_6_4; // @[Switch.scala 30:36:@275.4]
  wire  _T_771; // @[Switch.scala 30:53:@277.4]
  wire  valid_6_5; // @[Switch.scala 30:36:@278.4]
  wire  _T_774; // @[Switch.scala 30:53:@280.4]
  wire  valid_6_6; // @[Switch.scala 30:36:@281.4]
  wire  _T_777; // @[Switch.scala 30:53:@283.4]
  wire  valid_6_7; // @[Switch.scala 30:36:@284.4]
  wire [2:0] _T_787; // @[Mux.scala 31:69:@286.4]
  wire [2:0] _T_788; // @[Mux.scala 31:69:@287.4]
  wire [2:0] _T_789; // @[Mux.scala 31:69:@288.4]
  wire [2:0] _T_790; // @[Mux.scala 31:69:@289.4]
  wire [2:0] _T_791; // @[Mux.scala 31:69:@290.4]
  wire [2:0] _T_792; // @[Mux.scala 31:69:@291.4]
  wire [2:0] select_6; // @[Mux.scala 31:69:@292.4]
  wire [47:0] _GEN_49; // @[Switch.scala 33:19:@294.4]
  wire [47:0] _GEN_50; // @[Switch.scala 33:19:@294.4]
  wire [47:0] _GEN_51; // @[Switch.scala 33:19:@294.4]
  wire [47:0] _GEN_52; // @[Switch.scala 33:19:@294.4]
  wire [47:0] _GEN_53; // @[Switch.scala 33:19:@294.4]
  wire [47:0] _GEN_54; // @[Switch.scala 33:19:@294.4]
  wire [7:0] _T_801; // @[Switch.scala 34:32:@301.4]
  wire  _T_805; // @[Switch.scala 30:53:@304.4]
  wire  valid_7_0; // @[Switch.scala 30:36:@305.4]
  wire  _T_808; // @[Switch.scala 30:53:@307.4]
  wire  valid_7_1; // @[Switch.scala 30:36:@308.4]
  wire  _T_811; // @[Switch.scala 30:53:@310.4]
  wire  valid_7_2; // @[Switch.scala 30:36:@311.4]
  wire  _T_814; // @[Switch.scala 30:53:@313.4]
  wire  valid_7_3; // @[Switch.scala 30:36:@314.4]
  wire  _T_817; // @[Switch.scala 30:53:@316.4]
  wire  valid_7_4; // @[Switch.scala 30:36:@317.4]
  wire  _T_820; // @[Switch.scala 30:53:@319.4]
  wire  valid_7_5; // @[Switch.scala 30:36:@320.4]
  wire  _T_823; // @[Switch.scala 30:53:@322.4]
  wire  valid_7_6; // @[Switch.scala 30:36:@323.4]
  wire  _T_826; // @[Switch.scala 30:53:@325.4]
  wire  valid_7_7; // @[Switch.scala 30:36:@326.4]
  wire [2:0] _T_836; // @[Mux.scala 31:69:@328.4]
  wire [2:0] _T_837; // @[Mux.scala 31:69:@329.4]
  wire [2:0] _T_838; // @[Mux.scala 31:69:@330.4]
  wire [2:0] _T_839; // @[Mux.scala 31:69:@331.4]
  wire [2:0] _T_840; // @[Mux.scala 31:69:@332.4]
  wire [2:0] _T_841; // @[Mux.scala 31:69:@333.4]
  wire [2:0] select_7; // @[Mux.scala 31:69:@334.4]
  wire [47:0] _GEN_57; // @[Switch.scala 33:19:@336.4]
  wire [47:0] _GEN_58; // @[Switch.scala 33:19:@336.4]
  wire [47:0] _GEN_59; // @[Switch.scala 33:19:@336.4]
  wire [47:0] _GEN_60; // @[Switch.scala 33:19:@336.4]
  wire [47:0] _GEN_61; // @[Switch.scala 33:19:@336.4]
  wire [47:0] _GEN_62; // @[Switch.scala 33:19:@336.4]
  wire [7:0] _T_850; // @[Switch.scala 34:32:@343.4]
  wire  _T_1220; // @[Switch.scala 41:52:@347.4]
  wire  output_0_0; // @[Switch.scala 41:38:@348.4]
  wire  _T_1223; // @[Switch.scala 41:52:@350.4]
  wire  output_0_1; // @[Switch.scala 41:38:@351.4]
  wire  _T_1226; // @[Switch.scala 41:52:@353.4]
  wire  output_0_2; // @[Switch.scala 41:38:@354.4]
  wire  _T_1229; // @[Switch.scala 41:52:@356.4]
  wire  output_0_3; // @[Switch.scala 41:38:@357.4]
  wire  _T_1232; // @[Switch.scala 41:52:@359.4]
  wire  output_0_4; // @[Switch.scala 41:38:@360.4]
  wire  _T_1235; // @[Switch.scala 41:52:@362.4]
  wire  output_0_5; // @[Switch.scala 41:38:@363.4]
  wire  _T_1238; // @[Switch.scala 41:52:@365.4]
  wire  output_0_6; // @[Switch.scala 41:38:@366.4]
  wire  _T_1241; // @[Switch.scala 41:52:@368.4]
  wire  output_0_7; // @[Switch.scala 41:38:@369.4]
  wire [7:0] _T_1249; // @[Switch.scala 43:31:@377.4]
  wire  _T_1253; // @[Switch.scala 41:52:@380.4]
  wire  output_1_0; // @[Switch.scala 41:38:@381.4]
  wire  _T_1256; // @[Switch.scala 41:52:@383.4]
  wire  output_1_1; // @[Switch.scala 41:38:@384.4]
  wire  _T_1259; // @[Switch.scala 41:52:@386.4]
  wire  output_1_2; // @[Switch.scala 41:38:@387.4]
  wire  _T_1262; // @[Switch.scala 41:52:@389.4]
  wire  output_1_3; // @[Switch.scala 41:38:@390.4]
  wire  _T_1265; // @[Switch.scala 41:52:@392.4]
  wire  output_1_4; // @[Switch.scala 41:38:@393.4]
  wire  _T_1268; // @[Switch.scala 41:52:@395.4]
  wire  output_1_5; // @[Switch.scala 41:38:@396.4]
  wire  _T_1271; // @[Switch.scala 41:52:@398.4]
  wire  output_1_6; // @[Switch.scala 41:38:@399.4]
  wire  _T_1274; // @[Switch.scala 41:52:@401.4]
  wire  output_1_7; // @[Switch.scala 41:38:@402.4]
  wire [7:0] _T_1282; // @[Switch.scala 43:31:@410.4]
  wire  _T_1286; // @[Switch.scala 41:52:@413.4]
  wire  output_2_0; // @[Switch.scala 41:38:@414.4]
  wire  _T_1289; // @[Switch.scala 41:52:@416.4]
  wire  output_2_1; // @[Switch.scala 41:38:@417.4]
  wire  _T_1292; // @[Switch.scala 41:52:@419.4]
  wire  output_2_2; // @[Switch.scala 41:38:@420.4]
  wire  _T_1295; // @[Switch.scala 41:52:@422.4]
  wire  output_2_3; // @[Switch.scala 41:38:@423.4]
  wire  _T_1298; // @[Switch.scala 41:52:@425.4]
  wire  output_2_4; // @[Switch.scala 41:38:@426.4]
  wire  _T_1301; // @[Switch.scala 41:52:@428.4]
  wire  output_2_5; // @[Switch.scala 41:38:@429.4]
  wire  _T_1304; // @[Switch.scala 41:52:@431.4]
  wire  output_2_6; // @[Switch.scala 41:38:@432.4]
  wire  _T_1307; // @[Switch.scala 41:52:@434.4]
  wire  output_2_7; // @[Switch.scala 41:38:@435.4]
  wire [7:0] _T_1315; // @[Switch.scala 43:31:@443.4]
  wire  _T_1319; // @[Switch.scala 41:52:@446.4]
  wire  output_3_0; // @[Switch.scala 41:38:@447.4]
  wire  _T_1322; // @[Switch.scala 41:52:@449.4]
  wire  output_3_1; // @[Switch.scala 41:38:@450.4]
  wire  _T_1325; // @[Switch.scala 41:52:@452.4]
  wire  output_3_2; // @[Switch.scala 41:38:@453.4]
  wire  _T_1328; // @[Switch.scala 41:52:@455.4]
  wire  output_3_3; // @[Switch.scala 41:38:@456.4]
  wire  _T_1331; // @[Switch.scala 41:52:@458.4]
  wire  output_3_4; // @[Switch.scala 41:38:@459.4]
  wire  _T_1334; // @[Switch.scala 41:52:@461.4]
  wire  output_3_5; // @[Switch.scala 41:38:@462.4]
  wire  _T_1337; // @[Switch.scala 41:52:@464.4]
  wire  output_3_6; // @[Switch.scala 41:38:@465.4]
  wire  _T_1340; // @[Switch.scala 41:52:@467.4]
  wire  output_3_7; // @[Switch.scala 41:38:@468.4]
  wire [7:0] _T_1348; // @[Switch.scala 43:31:@476.4]
  wire  _T_1352; // @[Switch.scala 41:52:@479.4]
  wire  output_4_0; // @[Switch.scala 41:38:@480.4]
  wire  _T_1355; // @[Switch.scala 41:52:@482.4]
  wire  output_4_1; // @[Switch.scala 41:38:@483.4]
  wire  _T_1358; // @[Switch.scala 41:52:@485.4]
  wire  output_4_2; // @[Switch.scala 41:38:@486.4]
  wire  _T_1361; // @[Switch.scala 41:52:@488.4]
  wire  output_4_3; // @[Switch.scala 41:38:@489.4]
  wire  _T_1364; // @[Switch.scala 41:52:@491.4]
  wire  output_4_4; // @[Switch.scala 41:38:@492.4]
  wire  _T_1367; // @[Switch.scala 41:52:@494.4]
  wire  output_4_5; // @[Switch.scala 41:38:@495.4]
  wire  _T_1370; // @[Switch.scala 41:52:@497.4]
  wire  output_4_6; // @[Switch.scala 41:38:@498.4]
  wire  _T_1373; // @[Switch.scala 41:52:@500.4]
  wire  output_4_7; // @[Switch.scala 41:38:@501.4]
  wire [7:0] _T_1381; // @[Switch.scala 43:31:@509.4]
  wire  _T_1385; // @[Switch.scala 41:52:@512.4]
  wire  output_5_0; // @[Switch.scala 41:38:@513.4]
  wire  _T_1388; // @[Switch.scala 41:52:@515.4]
  wire  output_5_1; // @[Switch.scala 41:38:@516.4]
  wire  _T_1391; // @[Switch.scala 41:52:@518.4]
  wire  output_5_2; // @[Switch.scala 41:38:@519.4]
  wire  _T_1394; // @[Switch.scala 41:52:@521.4]
  wire  output_5_3; // @[Switch.scala 41:38:@522.4]
  wire  _T_1397; // @[Switch.scala 41:52:@524.4]
  wire  output_5_4; // @[Switch.scala 41:38:@525.4]
  wire  _T_1400; // @[Switch.scala 41:52:@527.4]
  wire  output_5_5; // @[Switch.scala 41:38:@528.4]
  wire  _T_1403; // @[Switch.scala 41:52:@530.4]
  wire  output_5_6; // @[Switch.scala 41:38:@531.4]
  wire  _T_1406; // @[Switch.scala 41:52:@533.4]
  wire  output_5_7; // @[Switch.scala 41:38:@534.4]
  wire [7:0] _T_1414; // @[Switch.scala 43:31:@542.4]
  wire  _T_1418; // @[Switch.scala 41:52:@545.4]
  wire  output_6_0; // @[Switch.scala 41:38:@546.4]
  wire  _T_1421; // @[Switch.scala 41:52:@548.4]
  wire  output_6_1; // @[Switch.scala 41:38:@549.4]
  wire  _T_1424; // @[Switch.scala 41:52:@551.4]
  wire  output_6_2; // @[Switch.scala 41:38:@552.4]
  wire  _T_1427; // @[Switch.scala 41:52:@554.4]
  wire  output_6_3; // @[Switch.scala 41:38:@555.4]
  wire  _T_1430; // @[Switch.scala 41:52:@557.4]
  wire  output_6_4; // @[Switch.scala 41:38:@558.4]
  wire  _T_1433; // @[Switch.scala 41:52:@560.4]
  wire  output_6_5; // @[Switch.scala 41:38:@561.4]
  wire  _T_1436; // @[Switch.scala 41:52:@563.4]
  wire  output_6_6; // @[Switch.scala 41:38:@564.4]
  wire  _T_1439; // @[Switch.scala 41:52:@566.4]
  wire  output_6_7; // @[Switch.scala 41:38:@567.4]
  wire [7:0] _T_1447; // @[Switch.scala 43:31:@575.4]
  wire  _T_1451; // @[Switch.scala 41:52:@578.4]
  wire  output_7_0; // @[Switch.scala 41:38:@579.4]
  wire  _T_1454; // @[Switch.scala 41:52:@581.4]
  wire  output_7_1; // @[Switch.scala 41:38:@582.4]
  wire  _T_1457; // @[Switch.scala 41:52:@584.4]
  wire  output_7_2; // @[Switch.scala 41:38:@585.4]
  wire  _T_1460; // @[Switch.scala 41:52:@587.4]
  wire  output_7_3; // @[Switch.scala 41:38:@588.4]
  wire  _T_1463; // @[Switch.scala 41:52:@590.4]
  wire  output_7_4; // @[Switch.scala 41:38:@591.4]
  wire  _T_1466; // @[Switch.scala 41:52:@593.4]
  wire  output_7_5; // @[Switch.scala 41:38:@594.4]
  wire  _T_1469; // @[Switch.scala 41:52:@596.4]
  wire  output_7_6; // @[Switch.scala 41:38:@597.4]
  wire  _T_1472; // @[Switch.scala 41:52:@599.4]
  wire  output_7_7; // @[Switch.scala 41:38:@600.4]
  wire [7:0] _T_1480; // @[Switch.scala 43:31:@608.4]
  assign _T_462 = io_inAddr_0 == 3'h0; // @[Switch.scala 30:53:@10.4]
  assign valid_0_0 = io_inValid_0 & _T_462; // @[Switch.scala 30:36:@11.4]
  assign _T_465 = io_inAddr_1 == 3'h0; // @[Switch.scala 30:53:@13.4]
  assign valid_0_1 = io_inValid_1 & _T_465; // @[Switch.scala 30:36:@14.4]
  assign _T_468 = io_inAddr_2 == 3'h0; // @[Switch.scala 30:53:@16.4]
  assign valid_0_2 = io_inValid_2 & _T_468; // @[Switch.scala 30:36:@17.4]
  assign _T_471 = io_inAddr_3 == 3'h0; // @[Switch.scala 30:53:@19.4]
  assign valid_0_3 = io_inValid_3 & _T_471; // @[Switch.scala 30:36:@20.4]
  assign _T_474 = io_inAddr_4 == 3'h0; // @[Switch.scala 30:53:@22.4]
  assign valid_0_4 = io_inValid_4 & _T_474; // @[Switch.scala 30:36:@23.4]
  assign _T_477 = io_inAddr_5 == 3'h0; // @[Switch.scala 30:53:@25.4]
  assign valid_0_5 = io_inValid_5 & _T_477; // @[Switch.scala 30:36:@26.4]
  assign _T_480 = io_inAddr_6 == 3'h0; // @[Switch.scala 30:53:@28.4]
  assign valid_0_6 = io_inValid_6 & _T_480; // @[Switch.scala 30:36:@29.4]
  assign _T_483 = io_inAddr_7 == 3'h0; // @[Switch.scala 30:53:@31.4]
  assign valid_0_7 = io_inValid_7 & _T_483; // @[Switch.scala 30:36:@32.4]
  assign _T_493 = valid_0_6 ? 3'h6 : 3'h7; // @[Mux.scala 31:69:@34.4]
  assign _T_494 = valid_0_5 ? 3'h5 : _T_493; // @[Mux.scala 31:69:@35.4]
  assign _T_495 = valid_0_4 ? 3'h4 : _T_494; // @[Mux.scala 31:69:@36.4]
  assign _T_496 = valid_0_3 ? 3'h3 : _T_495; // @[Mux.scala 31:69:@37.4]
  assign _T_497 = valid_0_2 ? 3'h2 : _T_496; // @[Mux.scala 31:69:@38.4]
  assign _T_498 = valid_0_1 ? 3'h1 : _T_497; // @[Mux.scala 31:69:@39.4]
  assign select_0 = valid_0_0 ? 3'h0 : _T_498; // @[Mux.scala 31:69:@40.4]
  assign _GEN_1 = 3'h1 == select_0 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@42.4]
  assign _GEN_2 = 3'h2 == select_0 ? io_inData_2 : _GEN_1; // @[Switch.scala 33:19:@42.4]
  assign _GEN_3 = 3'h3 == select_0 ? io_inData_3 : _GEN_2; // @[Switch.scala 33:19:@42.4]
  assign _GEN_4 = 3'h4 == select_0 ? io_inData_4 : _GEN_3; // @[Switch.scala 33:19:@42.4]
  assign _GEN_5 = 3'h5 == select_0 ? io_inData_5 : _GEN_4; // @[Switch.scala 33:19:@42.4]
  assign _GEN_6 = 3'h6 == select_0 ? io_inData_6 : _GEN_5; // @[Switch.scala 33:19:@42.4]
  assign _T_507 = {valid_0_7,valid_0_6,valid_0_5,valid_0_4,valid_0_3,valid_0_2,valid_0_1,valid_0_0}; // @[Switch.scala 34:32:@49.4]
  assign _T_511 = io_inAddr_0 == 3'h1; // @[Switch.scala 30:53:@52.4]
  assign valid_1_0 = io_inValid_0 & _T_511; // @[Switch.scala 30:36:@53.4]
  assign _T_514 = io_inAddr_1 == 3'h1; // @[Switch.scala 30:53:@55.4]
  assign valid_1_1 = io_inValid_1 & _T_514; // @[Switch.scala 30:36:@56.4]
  assign _T_517 = io_inAddr_2 == 3'h1; // @[Switch.scala 30:53:@58.4]
  assign valid_1_2 = io_inValid_2 & _T_517; // @[Switch.scala 30:36:@59.4]
  assign _T_520 = io_inAddr_3 == 3'h1; // @[Switch.scala 30:53:@61.4]
  assign valid_1_3 = io_inValid_3 & _T_520; // @[Switch.scala 30:36:@62.4]
  assign _T_523 = io_inAddr_4 == 3'h1; // @[Switch.scala 30:53:@64.4]
  assign valid_1_4 = io_inValid_4 & _T_523; // @[Switch.scala 30:36:@65.4]
  assign _T_526 = io_inAddr_5 == 3'h1; // @[Switch.scala 30:53:@67.4]
  assign valid_1_5 = io_inValid_5 & _T_526; // @[Switch.scala 30:36:@68.4]
  assign _T_529 = io_inAddr_6 == 3'h1; // @[Switch.scala 30:53:@70.4]
  assign valid_1_6 = io_inValid_6 & _T_529; // @[Switch.scala 30:36:@71.4]
  assign _T_532 = io_inAddr_7 == 3'h1; // @[Switch.scala 30:53:@73.4]
  assign valid_1_7 = io_inValid_7 & _T_532; // @[Switch.scala 30:36:@74.4]
  assign _T_542 = valid_1_6 ? 3'h6 : 3'h7; // @[Mux.scala 31:69:@76.4]
  assign _T_543 = valid_1_5 ? 3'h5 : _T_542; // @[Mux.scala 31:69:@77.4]
  assign _T_544 = valid_1_4 ? 3'h4 : _T_543; // @[Mux.scala 31:69:@78.4]
  assign _T_545 = valid_1_3 ? 3'h3 : _T_544; // @[Mux.scala 31:69:@79.4]
  assign _T_546 = valid_1_2 ? 3'h2 : _T_545; // @[Mux.scala 31:69:@80.4]
  assign _T_547 = valid_1_1 ? 3'h1 : _T_546; // @[Mux.scala 31:69:@81.4]
  assign select_1 = valid_1_0 ? 3'h0 : _T_547; // @[Mux.scala 31:69:@82.4]
  assign _GEN_9 = 3'h1 == select_1 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@84.4]
  assign _GEN_10 = 3'h2 == select_1 ? io_inData_2 : _GEN_9; // @[Switch.scala 33:19:@84.4]
  assign _GEN_11 = 3'h3 == select_1 ? io_inData_3 : _GEN_10; // @[Switch.scala 33:19:@84.4]
  assign _GEN_12 = 3'h4 == select_1 ? io_inData_4 : _GEN_11; // @[Switch.scala 33:19:@84.4]
  assign _GEN_13 = 3'h5 == select_1 ? io_inData_5 : _GEN_12; // @[Switch.scala 33:19:@84.4]
  assign _GEN_14 = 3'h6 == select_1 ? io_inData_6 : _GEN_13; // @[Switch.scala 33:19:@84.4]
  assign _T_556 = {valid_1_7,valid_1_6,valid_1_5,valid_1_4,valid_1_3,valid_1_2,valid_1_1,valid_1_0}; // @[Switch.scala 34:32:@91.4]
  assign _T_560 = io_inAddr_0 == 3'h2; // @[Switch.scala 30:53:@94.4]
  assign valid_2_0 = io_inValid_0 & _T_560; // @[Switch.scala 30:36:@95.4]
  assign _T_563 = io_inAddr_1 == 3'h2; // @[Switch.scala 30:53:@97.4]
  assign valid_2_1 = io_inValid_1 & _T_563; // @[Switch.scala 30:36:@98.4]
  assign _T_566 = io_inAddr_2 == 3'h2; // @[Switch.scala 30:53:@100.4]
  assign valid_2_2 = io_inValid_2 & _T_566; // @[Switch.scala 30:36:@101.4]
  assign _T_569 = io_inAddr_3 == 3'h2; // @[Switch.scala 30:53:@103.4]
  assign valid_2_3 = io_inValid_3 & _T_569; // @[Switch.scala 30:36:@104.4]
  assign _T_572 = io_inAddr_4 == 3'h2; // @[Switch.scala 30:53:@106.4]
  assign valid_2_4 = io_inValid_4 & _T_572; // @[Switch.scala 30:36:@107.4]
  assign _T_575 = io_inAddr_5 == 3'h2; // @[Switch.scala 30:53:@109.4]
  assign valid_2_5 = io_inValid_5 & _T_575; // @[Switch.scala 30:36:@110.4]
  assign _T_578 = io_inAddr_6 == 3'h2; // @[Switch.scala 30:53:@112.4]
  assign valid_2_6 = io_inValid_6 & _T_578; // @[Switch.scala 30:36:@113.4]
  assign _T_581 = io_inAddr_7 == 3'h2; // @[Switch.scala 30:53:@115.4]
  assign valid_2_7 = io_inValid_7 & _T_581; // @[Switch.scala 30:36:@116.4]
  assign _T_591 = valid_2_6 ? 3'h6 : 3'h7; // @[Mux.scala 31:69:@118.4]
  assign _T_592 = valid_2_5 ? 3'h5 : _T_591; // @[Mux.scala 31:69:@119.4]
  assign _T_593 = valid_2_4 ? 3'h4 : _T_592; // @[Mux.scala 31:69:@120.4]
  assign _T_594 = valid_2_3 ? 3'h3 : _T_593; // @[Mux.scala 31:69:@121.4]
  assign _T_595 = valid_2_2 ? 3'h2 : _T_594; // @[Mux.scala 31:69:@122.4]
  assign _T_596 = valid_2_1 ? 3'h1 : _T_595; // @[Mux.scala 31:69:@123.4]
  assign select_2 = valid_2_0 ? 3'h0 : _T_596; // @[Mux.scala 31:69:@124.4]
  assign _GEN_17 = 3'h1 == select_2 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@126.4]
  assign _GEN_18 = 3'h2 == select_2 ? io_inData_2 : _GEN_17; // @[Switch.scala 33:19:@126.4]
  assign _GEN_19 = 3'h3 == select_2 ? io_inData_3 : _GEN_18; // @[Switch.scala 33:19:@126.4]
  assign _GEN_20 = 3'h4 == select_2 ? io_inData_4 : _GEN_19; // @[Switch.scala 33:19:@126.4]
  assign _GEN_21 = 3'h5 == select_2 ? io_inData_5 : _GEN_20; // @[Switch.scala 33:19:@126.4]
  assign _GEN_22 = 3'h6 == select_2 ? io_inData_6 : _GEN_21; // @[Switch.scala 33:19:@126.4]
  assign _T_605 = {valid_2_7,valid_2_6,valid_2_5,valid_2_4,valid_2_3,valid_2_2,valid_2_1,valid_2_0}; // @[Switch.scala 34:32:@133.4]
  assign _T_609 = io_inAddr_0 == 3'h3; // @[Switch.scala 30:53:@136.4]
  assign valid_3_0 = io_inValid_0 & _T_609; // @[Switch.scala 30:36:@137.4]
  assign _T_612 = io_inAddr_1 == 3'h3; // @[Switch.scala 30:53:@139.4]
  assign valid_3_1 = io_inValid_1 & _T_612; // @[Switch.scala 30:36:@140.4]
  assign _T_615 = io_inAddr_2 == 3'h3; // @[Switch.scala 30:53:@142.4]
  assign valid_3_2 = io_inValid_2 & _T_615; // @[Switch.scala 30:36:@143.4]
  assign _T_618 = io_inAddr_3 == 3'h3; // @[Switch.scala 30:53:@145.4]
  assign valid_3_3 = io_inValid_3 & _T_618; // @[Switch.scala 30:36:@146.4]
  assign _T_621 = io_inAddr_4 == 3'h3; // @[Switch.scala 30:53:@148.4]
  assign valid_3_4 = io_inValid_4 & _T_621; // @[Switch.scala 30:36:@149.4]
  assign _T_624 = io_inAddr_5 == 3'h3; // @[Switch.scala 30:53:@151.4]
  assign valid_3_5 = io_inValid_5 & _T_624; // @[Switch.scala 30:36:@152.4]
  assign _T_627 = io_inAddr_6 == 3'h3; // @[Switch.scala 30:53:@154.4]
  assign valid_3_6 = io_inValid_6 & _T_627; // @[Switch.scala 30:36:@155.4]
  assign _T_630 = io_inAddr_7 == 3'h3; // @[Switch.scala 30:53:@157.4]
  assign valid_3_7 = io_inValid_7 & _T_630; // @[Switch.scala 30:36:@158.4]
  assign _T_640 = valid_3_6 ? 3'h6 : 3'h7; // @[Mux.scala 31:69:@160.4]
  assign _T_641 = valid_3_5 ? 3'h5 : _T_640; // @[Mux.scala 31:69:@161.4]
  assign _T_642 = valid_3_4 ? 3'h4 : _T_641; // @[Mux.scala 31:69:@162.4]
  assign _T_643 = valid_3_3 ? 3'h3 : _T_642; // @[Mux.scala 31:69:@163.4]
  assign _T_644 = valid_3_2 ? 3'h2 : _T_643; // @[Mux.scala 31:69:@164.4]
  assign _T_645 = valid_3_1 ? 3'h1 : _T_644; // @[Mux.scala 31:69:@165.4]
  assign select_3 = valid_3_0 ? 3'h0 : _T_645; // @[Mux.scala 31:69:@166.4]
  assign _GEN_25 = 3'h1 == select_3 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@168.4]
  assign _GEN_26 = 3'h2 == select_3 ? io_inData_2 : _GEN_25; // @[Switch.scala 33:19:@168.4]
  assign _GEN_27 = 3'h3 == select_3 ? io_inData_3 : _GEN_26; // @[Switch.scala 33:19:@168.4]
  assign _GEN_28 = 3'h4 == select_3 ? io_inData_4 : _GEN_27; // @[Switch.scala 33:19:@168.4]
  assign _GEN_29 = 3'h5 == select_3 ? io_inData_5 : _GEN_28; // @[Switch.scala 33:19:@168.4]
  assign _GEN_30 = 3'h6 == select_3 ? io_inData_6 : _GEN_29; // @[Switch.scala 33:19:@168.4]
  assign _T_654 = {valid_3_7,valid_3_6,valid_3_5,valid_3_4,valid_3_3,valid_3_2,valid_3_1,valid_3_0}; // @[Switch.scala 34:32:@175.4]
  assign _T_658 = io_inAddr_0 == 3'h4; // @[Switch.scala 30:53:@178.4]
  assign valid_4_0 = io_inValid_0 & _T_658; // @[Switch.scala 30:36:@179.4]
  assign _T_661 = io_inAddr_1 == 3'h4; // @[Switch.scala 30:53:@181.4]
  assign valid_4_1 = io_inValid_1 & _T_661; // @[Switch.scala 30:36:@182.4]
  assign _T_664 = io_inAddr_2 == 3'h4; // @[Switch.scala 30:53:@184.4]
  assign valid_4_2 = io_inValid_2 & _T_664; // @[Switch.scala 30:36:@185.4]
  assign _T_667 = io_inAddr_3 == 3'h4; // @[Switch.scala 30:53:@187.4]
  assign valid_4_3 = io_inValid_3 & _T_667; // @[Switch.scala 30:36:@188.4]
  assign _T_670 = io_inAddr_4 == 3'h4; // @[Switch.scala 30:53:@190.4]
  assign valid_4_4 = io_inValid_4 & _T_670; // @[Switch.scala 30:36:@191.4]
  assign _T_673 = io_inAddr_5 == 3'h4; // @[Switch.scala 30:53:@193.4]
  assign valid_4_5 = io_inValid_5 & _T_673; // @[Switch.scala 30:36:@194.4]
  assign _T_676 = io_inAddr_6 == 3'h4; // @[Switch.scala 30:53:@196.4]
  assign valid_4_6 = io_inValid_6 & _T_676; // @[Switch.scala 30:36:@197.4]
  assign _T_679 = io_inAddr_7 == 3'h4; // @[Switch.scala 30:53:@199.4]
  assign valid_4_7 = io_inValid_7 & _T_679; // @[Switch.scala 30:36:@200.4]
  assign _T_689 = valid_4_6 ? 3'h6 : 3'h7; // @[Mux.scala 31:69:@202.4]
  assign _T_690 = valid_4_5 ? 3'h5 : _T_689; // @[Mux.scala 31:69:@203.4]
  assign _T_691 = valid_4_4 ? 3'h4 : _T_690; // @[Mux.scala 31:69:@204.4]
  assign _T_692 = valid_4_3 ? 3'h3 : _T_691; // @[Mux.scala 31:69:@205.4]
  assign _T_693 = valid_4_2 ? 3'h2 : _T_692; // @[Mux.scala 31:69:@206.4]
  assign _T_694 = valid_4_1 ? 3'h1 : _T_693; // @[Mux.scala 31:69:@207.4]
  assign select_4 = valid_4_0 ? 3'h0 : _T_694; // @[Mux.scala 31:69:@208.4]
  assign _GEN_33 = 3'h1 == select_4 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@210.4]
  assign _GEN_34 = 3'h2 == select_4 ? io_inData_2 : _GEN_33; // @[Switch.scala 33:19:@210.4]
  assign _GEN_35 = 3'h3 == select_4 ? io_inData_3 : _GEN_34; // @[Switch.scala 33:19:@210.4]
  assign _GEN_36 = 3'h4 == select_4 ? io_inData_4 : _GEN_35; // @[Switch.scala 33:19:@210.4]
  assign _GEN_37 = 3'h5 == select_4 ? io_inData_5 : _GEN_36; // @[Switch.scala 33:19:@210.4]
  assign _GEN_38 = 3'h6 == select_4 ? io_inData_6 : _GEN_37; // @[Switch.scala 33:19:@210.4]
  assign _T_703 = {valid_4_7,valid_4_6,valid_4_5,valid_4_4,valid_4_3,valid_4_2,valid_4_1,valid_4_0}; // @[Switch.scala 34:32:@217.4]
  assign _T_707 = io_inAddr_0 == 3'h5; // @[Switch.scala 30:53:@220.4]
  assign valid_5_0 = io_inValid_0 & _T_707; // @[Switch.scala 30:36:@221.4]
  assign _T_710 = io_inAddr_1 == 3'h5; // @[Switch.scala 30:53:@223.4]
  assign valid_5_1 = io_inValid_1 & _T_710; // @[Switch.scala 30:36:@224.4]
  assign _T_713 = io_inAddr_2 == 3'h5; // @[Switch.scala 30:53:@226.4]
  assign valid_5_2 = io_inValid_2 & _T_713; // @[Switch.scala 30:36:@227.4]
  assign _T_716 = io_inAddr_3 == 3'h5; // @[Switch.scala 30:53:@229.4]
  assign valid_5_3 = io_inValid_3 & _T_716; // @[Switch.scala 30:36:@230.4]
  assign _T_719 = io_inAddr_4 == 3'h5; // @[Switch.scala 30:53:@232.4]
  assign valid_5_4 = io_inValid_4 & _T_719; // @[Switch.scala 30:36:@233.4]
  assign _T_722 = io_inAddr_5 == 3'h5; // @[Switch.scala 30:53:@235.4]
  assign valid_5_5 = io_inValid_5 & _T_722; // @[Switch.scala 30:36:@236.4]
  assign _T_725 = io_inAddr_6 == 3'h5; // @[Switch.scala 30:53:@238.4]
  assign valid_5_6 = io_inValid_6 & _T_725; // @[Switch.scala 30:36:@239.4]
  assign _T_728 = io_inAddr_7 == 3'h5; // @[Switch.scala 30:53:@241.4]
  assign valid_5_7 = io_inValid_7 & _T_728; // @[Switch.scala 30:36:@242.4]
  assign _T_738 = valid_5_6 ? 3'h6 : 3'h7; // @[Mux.scala 31:69:@244.4]
  assign _T_739 = valid_5_5 ? 3'h5 : _T_738; // @[Mux.scala 31:69:@245.4]
  assign _T_740 = valid_5_4 ? 3'h4 : _T_739; // @[Mux.scala 31:69:@246.4]
  assign _T_741 = valid_5_3 ? 3'h3 : _T_740; // @[Mux.scala 31:69:@247.4]
  assign _T_742 = valid_5_2 ? 3'h2 : _T_741; // @[Mux.scala 31:69:@248.4]
  assign _T_743 = valid_5_1 ? 3'h1 : _T_742; // @[Mux.scala 31:69:@249.4]
  assign select_5 = valid_5_0 ? 3'h0 : _T_743; // @[Mux.scala 31:69:@250.4]
  assign _GEN_41 = 3'h1 == select_5 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@252.4]
  assign _GEN_42 = 3'h2 == select_5 ? io_inData_2 : _GEN_41; // @[Switch.scala 33:19:@252.4]
  assign _GEN_43 = 3'h3 == select_5 ? io_inData_3 : _GEN_42; // @[Switch.scala 33:19:@252.4]
  assign _GEN_44 = 3'h4 == select_5 ? io_inData_4 : _GEN_43; // @[Switch.scala 33:19:@252.4]
  assign _GEN_45 = 3'h5 == select_5 ? io_inData_5 : _GEN_44; // @[Switch.scala 33:19:@252.4]
  assign _GEN_46 = 3'h6 == select_5 ? io_inData_6 : _GEN_45; // @[Switch.scala 33:19:@252.4]
  assign _T_752 = {valid_5_7,valid_5_6,valid_5_5,valid_5_4,valid_5_3,valid_5_2,valid_5_1,valid_5_0}; // @[Switch.scala 34:32:@259.4]
  assign _T_756 = io_inAddr_0 == 3'h6; // @[Switch.scala 30:53:@262.4]
  assign valid_6_0 = io_inValid_0 & _T_756; // @[Switch.scala 30:36:@263.4]
  assign _T_759 = io_inAddr_1 == 3'h6; // @[Switch.scala 30:53:@265.4]
  assign valid_6_1 = io_inValid_1 & _T_759; // @[Switch.scala 30:36:@266.4]
  assign _T_762 = io_inAddr_2 == 3'h6; // @[Switch.scala 30:53:@268.4]
  assign valid_6_2 = io_inValid_2 & _T_762; // @[Switch.scala 30:36:@269.4]
  assign _T_765 = io_inAddr_3 == 3'h6; // @[Switch.scala 30:53:@271.4]
  assign valid_6_3 = io_inValid_3 & _T_765; // @[Switch.scala 30:36:@272.4]
  assign _T_768 = io_inAddr_4 == 3'h6; // @[Switch.scala 30:53:@274.4]
  assign valid_6_4 = io_inValid_4 & _T_768; // @[Switch.scala 30:36:@275.4]
  assign _T_771 = io_inAddr_5 == 3'h6; // @[Switch.scala 30:53:@277.4]
  assign valid_6_5 = io_inValid_5 & _T_771; // @[Switch.scala 30:36:@278.4]
  assign _T_774 = io_inAddr_6 == 3'h6; // @[Switch.scala 30:53:@280.4]
  assign valid_6_6 = io_inValid_6 & _T_774; // @[Switch.scala 30:36:@281.4]
  assign _T_777 = io_inAddr_7 == 3'h6; // @[Switch.scala 30:53:@283.4]
  assign valid_6_7 = io_inValid_7 & _T_777; // @[Switch.scala 30:36:@284.4]
  assign _T_787 = valid_6_6 ? 3'h6 : 3'h7; // @[Mux.scala 31:69:@286.4]
  assign _T_788 = valid_6_5 ? 3'h5 : _T_787; // @[Mux.scala 31:69:@287.4]
  assign _T_789 = valid_6_4 ? 3'h4 : _T_788; // @[Mux.scala 31:69:@288.4]
  assign _T_790 = valid_6_3 ? 3'h3 : _T_789; // @[Mux.scala 31:69:@289.4]
  assign _T_791 = valid_6_2 ? 3'h2 : _T_790; // @[Mux.scala 31:69:@290.4]
  assign _T_792 = valid_6_1 ? 3'h1 : _T_791; // @[Mux.scala 31:69:@291.4]
  assign select_6 = valid_6_0 ? 3'h0 : _T_792; // @[Mux.scala 31:69:@292.4]
  assign _GEN_49 = 3'h1 == select_6 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@294.4]
  assign _GEN_50 = 3'h2 == select_6 ? io_inData_2 : _GEN_49; // @[Switch.scala 33:19:@294.4]
  assign _GEN_51 = 3'h3 == select_6 ? io_inData_3 : _GEN_50; // @[Switch.scala 33:19:@294.4]
  assign _GEN_52 = 3'h4 == select_6 ? io_inData_4 : _GEN_51; // @[Switch.scala 33:19:@294.4]
  assign _GEN_53 = 3'h5 == select_6 ? io_inData_5 : _GEN_52; // @[Switch.scala 33:19:@294.4]
  assign _GEN_54 = 3'h6 == select_6 ? io_inData_6 : _GEN_53; // @[Switch.scala 33:19:@294.4]
  assign _T_801 = {valid_6_7,valid_6_6,valid_6_5,valid_6_4,valid_6_3,valid_6_2,valid_6_1,valid_6_0}; // @[Switch.scala 34:32:@301.4]
  assign _T_805 = io_inAddr_0 == 3'h7; // @[Switch.scala 30:53:@304.4]
  assign valid_7_0 = io_inValid_0 & _T_805; // @[Switch.scala 30:36:@305.4]
  assign _T_808 = io_inAddr_1 == 3'h7; // @[Switch.scala 30:53:@307.4]
  assign valid_7_1 = io_inValid_1 & _T_808; // @[Switch.scala 30:36:@308.4]
  assign _T_811 = io_inAddr_2 == 3'h7; // @[Switch.scala 30:53:@310.4]
  assign valid_7_2 = io_inValid_2 & _T_811; // @[Switch.scala 30:36:@311.4]
  assign _T_814 = io_inAddr_3 == 3'h7; // @[Switch.scala 30:53:@313.4]
  assign valid_7_3 = io_inValid_3 & _T_814; // @[Switch.scala 30:36:@314.4]
  assign _T_817 = io_inAddr_4 == 3'h7; // @[Switch.scala 30:53:@316.4]
  assign valid_7_4 = io_inValid_4 & _T_817; // @[Switch.scala 30:36:@317.4]
  assign _T_820 = io_inAddr_5 == 3'h7; // @[Switch.scala 30:53:@319.4]
  assign valid_7_5 = io_inValid_5 & _T_820; // @[Switch.scala 30:36:@320.4]
  assign _T_823 = io_inAddr_6 == 3'h7; // @[Switch.scala 30:53:@322.4]
  assign valid_7_6 = io_inValid_6 & _T_823; // @[Switch.scala 30:36:@323.4]
  assign _T_826 = io_inAddr_7 == 3'h7; // @[Switch.scala 30:53:@325.4]
  assign valid_7_7 = io_inValid_7 & _T_826; // @[Switch.scala 30:36:@326.4]
  assign _T_836 = valid_7_6 ? 3'h6 : 3'h7; // @[Mux.scala 31:69:@328.4]
  assign _T_837 = valid_7_5 ? 3'h5 : _T_836; // @[Mux.scala 31:69:@329.4]
  assign _T_838 = valid_7_4 ? 3'h4 : _T_837; // @[Mux.scala 31:69:@330.4]
  assign _T_839 = valid_7_3 ? 3'h3 : _T_838; // @[Mux.scala 31:69:@331.4]
  assign _T_840 = valid_7_2 ? 3'h2 : _T_839; // @[Mux.scala 31:69:@332.4]
  assign _T_841 = valid_7_1 ? 3'h1 : _T_840; // @[Mux.scala 31:69:@333.4]
  assign select_7 = valid_7_0 ? 3'h0 : _T_841; // @[Mux.scala 31:69:@334.4]
  assign _GEN_57 = 3'h1 == select_7 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@336.4]
  assign _GEN_58 = 3'h2 == select_7 ? io_inData_2 : _GEN_57; // @[Switch.scala 33:19:@336.4]
  assign _GEN_59 = 3'h3 == select_7 ? io_inData_3 : _GEN_58; // @[Switch.scala 33:19:@336.4]
  assign _GEN_60 = 3'h4 == select_7 ? io_inData_4 : _GEN_59; // @[Switch.scala 33:19:@336.4]
  assign _GEN_61 = 3'h5 == select_7 ? io_inData_5 : _GEN_60; // @[Switch.scala 33:19:@336.4]
  assign _GEN_62 = 3'h6 == select_7 ? io_inData_6 : _GEN_61; // @[Switch.scala 33:19:@336.4]
  assign _T_850 = {valid_7_7,valid_7_6,valid_7_5,valid_7_4,valid_7_3,valid_7_2,valid_7_1,valid_7_0}; // @[Switch.scala 34:32:@343.4]
  assign _T_1220 = select_0 == 3'h0; // @[Switch.scala 41:52:@347.4]
  assign output_0_0 = io_outValid_0 & _T_1220; // @[Switch.scala 41:38:@348.4]
  assign _T_1223 = select_1 == 3'h0; // @[Switch.scala 41:52:@350.4]
  assign output_0_1 = io_outValid_1 & _T_1223; // @[Switch.scala 41:38:@351.4]
  assign _T_1226 = select_2 == 3'h0; // @[Switch.scala 41:52:@353.4]
  assign output_0_2 = io_outValid_2 & _T_1226; // @[Switch.scala 41:38:@354.4]
  assign _T_1229 = select_3 == 3'h0; // @[Switch.scala 41:52:@356.4]
  assign output_0_3 = io_outValid_3 & _T_1229; // @[Switch.scala 41:38:@357.4]
  assign _T_1232 = select_4 == 3'h0; // @[Switch.scala 41:52:@359.4]
  assign output_0_4 = io_outValid_4 & _T_1232; // @[Switch.scala 41:38:@360.4]
  assign _T_1235 = select_5 == 3'h0; // @[Switch.scala 41:52:@362.4]
  assign output_0_5 = io_outValid_5 & _T_1235; // @[Switch.scala 41:38:@363.4]
  assign _T_1238 = select_6 == 3'h0; // @[Switch.scala 41:52:@365.4]
  assign output_0_6 = io_outValid_6 & _T_1238; // @[Switch.scala 41:38:@366.4]
  assign _T_1241 = select_7 == 3'h0; // @[Switch.scala 41:52:@368.4]
  assign output_0_7 = io_outValid_7 & _T_1241; // @[Switch.scala 41:38:@369.4]
  assign _T_1249 = {output_0_7,output_0_6,output_0_5,output_0_4,output_0_3,output_0_2,output_0_1,output_0_0}; // @[Switch.scala 43:31:@377.4]
  assign _T_1253 = select_0 == 3'h1; // @[Switch.scala 41:52:@380.4]
  assign output_1_0 = io_outValid_0 & _T_1253; // @[Switch.scala 41:38:@381.4]
  assign _T_1256 = select_1 == 3'h1; // @[Switch.scala 41:52:@383.4]
  assign output_1_1 = io_outValid_1 & _T_1256; // @[Switch.scala 41:38:@384.4]
  assign _T_1259 = select_2 == 3'h1; // @[Switch.scala 41:52:@386.4]
  assign output_1_2 = io_outValid_2 & _T_1259; // @[Switch.scala 41:38:@387.4]
  assign _T_1262 = select_3 == 3'h1; // @[Switch.scala 41:52:@389.4]
  assign output_1_3 = io_outValid_3 & _T_1262; // @[Switch.scala 41:38:@390.4]
  assign _T_1265 = select_4 == 3'h1; // @[Switch.scala 41:52:@392.4]
  assign output_1_4 = io_outValid_4 & _T_1265; // @[Switch.scala 41:38:@393.4]
  assign _T_1268 = select_5 == 3'h1; // @[Switch.scala 41:52:@395.4]
  assign output_1_5 = io_outValid_5 & _T_1268; // @[Switch.scala 41:38:@396.4]
  assign _T_1271 = select_6 == 3'h1; // @[Switch.scala 41:52:@398.4]
  assign output_1_6 = io_outValid_6 & _T_1271; // @[Switch.scala 41:38:@399.4]
  assign _T_1274 = select_7 == 3'h1; // @[Switch.scala 41:52:@401.4]
  assign output_1_7 = io_outValid_7 & _T_1274; // @[Switch.scala 41:38:@402.4]
  assign _T_1282 = {output_1_7,output_1_6,output_1_5,output_1_4,output_1_3,output_1_2,output_1_1,output_1_0}; // @[Switch.scala 43:31:@410.4]
  assign _T_1286 = select_0 == 3'h2; // @[Switch.scala 41:52:@413.4]
  assign output_2_0 = io_outValid_0 & _T_1286; // @[Switch.scala 41:38:@414.4]
  assign _T_1289 = select_1 == 3'h2; // @[Switch.scala 41:52:@416.4]
  assign output_2_1 = io_outValid_1 & _T_1289; // @[Switch.scala 41:38:@417.4]
  assign _T_1292 = select_2 == 3'h2; // @[Switch.scala 41:52:@419.4]
  assign output_2_2 = io_outValid_2 & _T_1292; // @[Switch.scala 41:38:@420.4]
  assign _T_1295 = select_3 == 3'h2; // @[Switch.scala 41:52:@422.4]
  assign output_2_3 = io_outValid_3 & _T_1295; // @[Switch.scala 41:38:@423.4]
  assign _T_1298 = select_4 == 3'h2; // @[Switch.scala 41:52:@425.4]
  assign output_2_4 = io_outValid_4 & _T_1298; // @[Switch.scala 41:38:@426.4]
  assign _T_1301 = select_5 == 3'h2; // @[Switch.scala 41:52:@428.4]
  assign output_2_5 = io_outValid_5 & _T_1301; // @[Switch.scala 41:38:@429.4]
  assign _T_1304 = select_6 == 3'h2; // @[Switch.scala 41:52:@431.4]
  assign output_2_6 = io_outValid_6 & _T_1304; // @[Switch.scala 41:38:@432.4]
  assign _T_1307 = select_7 == 3'h2; // @[Switch.scala 41:52:@434.4]
  assign output_2_7 = io_outValid_7 & _T_1307; // @[Switch.scala 41:38:@435.4]
  assign _T_1315 = {output_2_7,output_2_6,output_2_5,output_2_4,output_2_3,output_2_2,output_2_1,output_2_0}; // @[Switch.scala 43:31:@443.4]
  assign _T_1319 = select_0 == 3'h3; // @[Switch.scala 41:52:@446.4]
  assign output_3_0 = io_outValid_0 & _T_1319; // @[Switch.scala 41:38:@447.4]
  assign _T_1322 = select_1 == 3'h3; // @[Switch.scala 41:52:@449.4]
  assign output_3_1 = io_outValid_1 & _T_1322; // @[Switch.scala 41:38:@450.4]
  assign _T_1325 = select_2 == 3'h3; // @[Switch.scala 41:52:@452.4]
  assign output_3_2 = io_outValid_2 & _T_1325; // @[Switch.scala 41:38:@453.4]
  assign _T_1328 = select_3 == 3'h3; // @[Switch.scala 41:52:@455.4]
  assign output_3_3 = io_outValid_3 & _T_1328; // @[Switch.scala 41:38:@456.4]
  assign _T_1331 = select_4 == 3'h3; // @[Switch.scala 41:52:@458.4]
  assign output_3_4 = io_outValid_4 & _T_1331; // @[Switch.scala 41:38:@459.4]
  assign _T_1334 = select_5 == 3'h3; // @[Switch.scala 41:52:@461.4]
  assign output_3_5 = io_outValid_5 & _T_1334; // @[Switch.scala 41:38:@462.4]
  assign _T_1337 = select_6 == 3'h3; // @[Switch.scala 41:52:@464.4]
  assign output_3_6 = io_outValid_6 & _T_1337; // @[Switch.scala 41:38:@465.4]
  assign _T_1340 = select_7 == 3'h3; // @[Switch.scala 41:52:@467.4]
  assign output_3_7 = io_outValid_7 & _T_1340; // @[Switch.scala 41:38:@468.4]
  assign _T_1348 = {output_3_7,output_3_6,output_3_5,output_3_4,output_3_3,output_3_2,output_3_1,output_3_0}; // @[Switch.scala 43:31:@476.4]
  assign _T_1352 = select_0 == 3'h4; // @[Switch.scala 41:52:@479.4]
  assign output_4_0 = io_outValid_0 & _T_1352; // @[Switch.scala 41:38:@480.4]
  assign _T_1355 = select_1 == 3'h4; // @[Switch.scala 41:52:@482.4]
  assign output_4_1 = io_outValid_1 & _T_1355; // @[Switch.scala 41:38:@483.4]
  assign _T_1358 = select_2 == 3'h4; // @[Switch.scala 41:52:@485.4]
  assign output_4_2 = io_outValid_2 & _T_1358; // @[Switch.scala 41:38:@486.4]
  assign _T_1361 = select_3 == 3'h4; // @[Switch.scala 41:52:@488.4]
  assign output_4_3 = io_outValid_3 & _T_1361; // @[Switch.scala 41:38:@489.4]
  assign _T_1364 = select_4 == 3'h4; // @[Switch.scala 41:52:@491.4]
  assign output_4_4 = io_outValid_4 & _T_1364; // @[Switch.scala 41:38:@492.4]
  assign _T_1367 = select_5 == 3'h4; // @[Switch.scala 41:52:@494.4]
  assign output_4_5 = io_outValid_5 & _T_1367; // @[Switch.scala 41:38:@495.4]
  assign _T_1370 = select_6 == 3'h4; // @[Switch.scala 41:52:@497.4]
  assign output_4_6 = io_outValid_6 & _T_1370; // @[Switch.scala 41:38:@498.4]
  assign _T_1373 = select_7 == 3'h4; // @[Switch.scala 41:52:@500.4]
  assign output_4_7 = io_outValid_7 & _T_1373; // @[Switch.scala 41:38:@501.4]
  assign _T_1381 = {output_4_7,output_4_6,output_4_5,output_4_4,output_4_3,output_4_2,output_4_1,output_4_0}; // @[Switch.scala 43:31:@509.4]
  assign _T_1385 = select_0 == 3'h5; // @[Switch.scala 41:52:@512.4]
  assign output_5_0 = io_outValid_0 & _T_1385; // @[Switch.scala 41:38:@513.4]
  assign _T_1388 = select_1 == 3'h5; // @[Switch.scala 41:52:@515.4]
  assign output_5_1 = io_outValid_1 & _T_1388; // @[Switch.scala 41:38:@516.4]
  assign _T_1391 = select_2 == 3'h5; // @[Switch.scala 41:52:@518.4]
  assign output_5_2 = io_outValid_2 & _T_1391; // @[Switch.scala 41:38:@519.4]
  assign _T_1394 = select_3 == 3'h5; // @[Switch.scala 41:52:@521.4]
  assign output_5_3 = io_outValid_3 & _T_1394; // @[Switch.scala 41:38:@522.4]
  assign _T_1397 = select_4 == 3'h5; // @[Switch.scala 41:52:@524.4]
  assign output_5_4 = io_outValid_4 & _T_1397; // @[Switch.scala 41:38:@525.4]
  assign _T_1400 = select_5 == 3'h5; // @[Switch.scala 41:52:@527.4]
  assign output_5_5 = io_outValid_5 & _T_1400; // @[Switch.scala 41:38:@528.4]
  assign _T_1403 = select_6 == 3'h5; // @[Switch.scala 41:52:@530.4]
  assign output_5_6 = io_outValid_6 & _T_1403; // @[Switch.scala 41:38:@531.4]
  assign _T_1406 = select_7 == 3'h5; // @[Switch.scala 41:52:@533.4]
  assign output_5_7 = io_outValid_7 & _T_1406; // @[Switch.scala 41:38:@534.4]
  assign _T_1414 = {output_5_7,output_5_6,output_5_5,output_5_4,output_5_3,output_5_2,output_5_1,output_5_0}; // @[Switch.scala 43:31:@542.4]
  assign _T_1418 = select_0 == 3'h6; // @[Switch.scala 41:52:@545.4]
  assign output_6_0 = io_outValid_0 & _T_1418; // @[Switch.scala 41:38:@546.4]
  assign _T_1421 = select_1 == 3'h6; // @[Switch.scala 41:52:@548.4]
  assign output_6_1 = io_outValid_1 & _T_1421; // @[Switch.scala 41:38:@549.4]
  assign _T_1424 = select_2 == 3'h6; // @[Switch.scala 41:52:@551.4]
  assign output_6_2 = io_outValid_2 & _T_1424; // @[Switch.scala 41:38:@552.4]
  assign _T_1427 = select_3 == 3'h6; // @[Switch.scala 41:52:@554.4]
  assign output_6_3 = io_outValid_3 & _T_1427; // @[Switch.scala 41:38:@555.4]
  assign _T_1430 = select_4 == 3'h6; // @[Switch.scala 41:52:@557.4]
  assign output_6_4 = io_outValid_4 & _T_1430; // @[Switch.scala 41:38:@558.4]
  assign _T_1433 = select_5 == 3'h6; // @[Switch.scala 41:52:@560.4]
  assign output_6_5 = io_outValid_5 & _T_1433; // @[Switch.scala 41:38:@561.4]
  assign _T_1436 = select_6 == 3'h6; // @[Switch.scala 41:52:@563.4]
  assign output_6_6 = io_outValid_6 & _T_1436; // @[Switch.scala 41:38:@564.4]
  assign _T_1439 = select_7 == 3'h6; // @[Switch.scala 41:52:@566.4]
  assign output_6_7 = io_outValid_7 & _T_1439; // @[Switch.scala 41:38:@567.4]
  assign _T_1447 = {output_6_7,output_6_6,output_6_5,output_6_4,output_6_3,output_6_2,output_6_1,output_6_0}; // @[Switch.scala 43:31:@575.4]
  assign _T_1451 = select_0 == 3'h7; // @[Switch.scala 41:52:@578.4]
  assign output_7_0 = io_outValid_0 & _T_1451; // @[Switch.scala 41:38:@579.4]
  assign _T_1454 = select_1 == 3'h7; // @[Switch.scala 41:52:@581.4]
  assign output_7_1 = io_outValid_1 & _T_1454; // @[Switch.scala 41:38:@582.4]
  assign _T_1457 = select_2 == 3'h7; // @[Switch.scala 41:52:@584.4]
  assign output_7_2 = io_outValid_2 & _T_1457; // @[Switch.scala 41:38:@585.4]
  assign _T_1460 = select_3 == 3'h7; // @[Switch.scala 41:52:@587.4]
  assign output_7_3 = io_outValid_3 & _T_1460; // @[Switch.scala 41:38:@588.4]
  assign _T_1463 = select_4 == 3'h7; // @[Switch.scala 41:52:@590.4]
  assign output_7_4 = io_outValid_4 & _T_1463; // @[Switch.scala 41:38:@591.4]
  assign _T_1466 = select_5 == 3'h7; // @[Switch.scala 41:52:@593.4]
  assign output_7_5 = io_outValid_5 & _T_1466; // @[Switch.scala 41:38:@594.4]
  assign _T_1469 = select_6 == 3'h7; // @[Switch.scala 41:52:@596.4]
  assign output_7_6 = io_outValid_6 & _T_1469; // @[Switch.scala 41:38:@597.4]
  assign _T_1472 = select_7 == 3'h7; // @[Switch.scala 41:52:@599.4]
  assign output_7_7 = io_outValid_7 & _T_1472; // @[Switch.scala 41:38:@600.4]
  assign _T_1480 = {output_7_7,output_7_6,output_7_5,output_7_4,output_7_3,output_7_2,output_7_1,output_7_0}; // @[Switch.scala 43:31:@608.4]
  assign io_outAck_0 = _T_1249 != 8'h0; // @[Switch.scala 43:18:@379.4]
  assign io_outAck_1 = _T_1282 != 8'h0; // @[Switch.scala 43:18:@412.4]
  assign io_outAck_2 = _T_1315 != 8'h0; // @[Switch.scala 43:18:@445.4]
  assign io_outAck_3 = _T_1348 != 8'h0; // @[Switch.scala 43:18:@478.4]
  assign io_outAck_4 = _T_1381 != 8'h0; // @[Switch.scala 43:18:@511.4]
  assign io_outAck_5 = _T_1414 != 8'h0; // @[Switch.scala 43:18:@544.4]
  assign io_outAck_6 = _T_1447 != 8'h0; // @[Switch.scala 43:18:@577.4]
  assign io_outAck_7 = _T_1480 != 8'h0; // @[Switch.scala 43:18:@610.4]
  assign io_outData_0 = 3'h7 == select_0 ? io_inData_7 : _GEN_6; // @[Switch.scala 33:19:@42.4]
  assign io_outData_1 = 3'h7 == select_1 ? io_inData_7 : _GEN_14; // @[Switch.scala 33:19:@84.4]
  assign io_outData_2 = 3'h7 == select_2 ? io_inData_7 : _GEN_22; // @[Switch.scala 33:19:@126.4]
  assign io_outData_3 = 3'h7 == select_3 ? io_inData_7 : _GEN_30; // @[Switch.scala 33:19:@168.4]
  assign io_outData_4 = 3'h7 == select_4 ? io_inData_7 : _GEN_38; // @[Switch.scala 33:19:@210.4]
  assign io_outData_5 = 3'h7 == select_5 ? io_inData_7 : _GEN_46; // @[Switch.scala 33:19:@252.4]
  assign io_outData_6 = 3'h7 == select_6 ? io_inData_7 : _GEN_54; // @[Switch.scala 33:19:@294.4]
  assign io_outData_7 = 3'h7 == select_7 ? io_inData_7 : _GEN_62; // @[Switch.scala 33:19:@336.4]
  assign io_outValid_0 = _T_507 != 8'h0; // @[Switch.scala 34:20:@51.4]
  assign io_outValid_1 = _T_556 != 8'h0; // @[Switch.scala 34:20:@93.4]
  assign io_outValid_2 = _T_605 != 8'h0; // @[Switch.scala 34:20:@135.4]
  assign io_outValid_3 = _T_654 != 8'h0; // @[Switch.scala 34:20:@177.4]
  assign io_outValid_4 = _T_703 != 8'h0; // @[Switch.scala 34:20:@219.4]
  assign io_outValid_5 = _T_752 != 8'h0; // @[Switch.scala 34:20:@261.4]
  assign io_outValid_6 = _T_801 != 8'h0; // @[Switch.scala 34:20:@303.4]
  assign io_outValid_7 = _T_850 != 8'h0; // @[Switch.scala 34:20:@345.4]
endmodule
module SwitchWrapper( // @[:@612.2]
  input         clock, // @[:@613.4]
  input         reset, // @[:@614.4]
  input  [2:0]  io_inAddr_0, // @[:@615.4]
  input  [2:0]  io_inAddr_1, // @[:@615.4]
  input  [2:0]  io_inAddr_2, // @[:@615.4]
  input  [2:0]  io_inAddr_3, // @[:@615.4]
  input  [2:0]  io_inAddr_4, // @[:@615.4]
  input  [2:0]  io_inAddr_5, // @[:@615.4]
  input  [2:0]  io_inAddr_6, // @[:@615.4]
  input  [2:0]  io_inAddr_7, // @[:@615.4]
  input  [47:0] io_inData_0, // @[:@615.4]
  input  [47:0] io_inData_1, // @[:@615.4]
  input  [47:0] io_inData_2, // @[:@615.4]
  input  [47:0] io_inData_3, // @[:@615.4]
  input  [47:0] io_inData_4, // @[:@615.4]
  input  [47:0] io_inData_5, // @[:@615.4]
  input  [47:0] io_inData_6, // @[:@615.4]
  input  [47:0] io_inData_7, // @[:@615.4]
  input         io_inValid_0, // @[:@615.4]
  input         io_inValid_1, // @[:@615.4]
  input         io_inValid_2, // @[:@615.4]
  input         io_inValid_3, // @[:@615.4]
  input         io_inValid_4, // @[:@615.4]
  input         io_inValid_5, // @[:@615.4]
  input         io_inValid_6, // @[:@615.4]
  input         io_inValid_7, // @[:@615.4]
  output        io_outAck_0, // @[:@615.4]
  output        io_outAck_1, // @[:@615.4]
  output        io_outAck_2, // @[:@615.4]
  output        io_outAck_3, // @[:@615.4]
  output        io_outAck_4, // @[:@615.4]
  output        io_outAck_5, // @[:@615.4]
  output        io_outAck_6, // @[:@615.4]
  output        io_outAck_7, // @[:@615.4]
  output [47:0] io_outData_0, // @[:@615.4]
  output [47:0] io_outData_1, // @[:@615.4]
  output [47:0] io_outData_2, // @[:@615.4]
  output [47:0] io_outData_3, // @[:@615.4]
  output [47:0] io_outData_4, // @[:@615.4]
  output [47:0] io_outData_5, // @[:@615.4]
  output [47:0] io_outData_6, // @[:@615.4]
  output [47:0] io_outData_7, // @[:@615.4]
  output        io_outValid_0, // @[:@615.4]
  output        io_outValid_1, // @[:@615.4]
  output        io_outValid_2, // @[:@615.4]
  output        io_outValid_3, // @[:@615.4]
  output        io_outValid_4, // @[:@615.4]
  output        io_outValid_5, // @[:@615.4]
  output        io_outValid_6, // @[:@615.4]
  output        io_outValid_7 // @[:@615.4]
);
  wire [2:0] switch_io_inAddr_0; // @[Switch.scala 50:22:@617.4]
  wire [2:0] switch_io_inAddr_1; // @[Switch.scala 50:22:@617.4]
  wire [2:0] switch_io_inAddr_2; // @[Switch.scala 50:22:@617.4]
  wire [2:0] switch_io_inAddr_3; // @[Switch.scala 50:22:@617.4]
  wire [2:0] switch_io_inAddr_4; // @[Switch.scala 50:22:@617.4]
  wire [2:0] switch_io_inAddr_5; // @[Switch.scala 50:22:@617.4]
  wire [2:0] switch_io_inAddr_6; // @[Switch.scala 50:22:@617.4]
  wire [2:0] switch_io_inAddr_7; // @[Switch.scala 50:22:@617.4]
  wire [47:0] switch_io_inData_0; // @[Switch.scala 50:22:@617.4]
  wire [47:0] switch_io_inData_1; // @[Switch.scala 50:22:@617.4]
  wire [47:0] switch_io_inData_2; // @[Switch.scala 50:22:@617.4]
  wire [47:0] switch_io_inData_3; // @[Switch.scala 50:22:@617.4]
  wire [47:0] switch_io_inData_4; // @[Switch.scala 50:22:@617.4]
  wire [47:0] switch_io_inData_5; // @[Switch.scala 50:22:@617.4]
  wire [47:0] switch_io_inData_6; // @[Switch.scala 50:22:@617.4]
  wire [47:0] switch_io_inData_7; // @[Switch.scala 50:22:@617.4]
  wire  switch_io_inValid_0; // @[Switch.scala 50:22:@617.4]
  wire  switch_io_inValid_1; // @[Switch.scala 50:22:@617.4]
  wire  switch_io_inValid_2; // @[Switch.scala 50:22:@617.4]
  wire  switch_io_inValid_3; // @[Switch.scala 50:22:@617.4]
  wire  switch_io_inValid_4; // @[Switch.scala 50:22:@617.4]
  wire  switch_io_inValid_5; // @[Switch.scala 50:22:@617.4]
  wire  switch_io_inValid_6; // @[Switch.scala 50:22:@617.4]
  wire  switch_io_inValid_7; // @[Switch.scala 50:22:@617.4]
  wire  switch_io_outAck_0; // @[Switch.scala 50:22:@617.4]
  wire  switch_io_outAck_1; // @[Switch.scala 50:22:@617.4]
  wire  switch_io_outAck_2; // @[Switch.scala 50:22:@617.4]
  wire  switch_io_outAck_3; // @[Switch.scala 50:22:@617.4]
  wire  switch_io_outAck_4; // @[Switch.scala 50:22:@617.4]
  wire  switch_io_outAck_5; // @[Switch.scala 50:22:@617.4]
  wire  switch_io_outAck_6; // @[Switch.scala 50:22:@617.4]
  wire  switch_io_outAck_7; // @[Switch.scala 50:22:@617.4]
  wire [47:0] switch_io_outData_0; // @[Switch.scala 50:22:@617.4]
  wire [47:0] switch_io_outData_1; // @[Switch.scala 50:22:@617.4]
  wire [47:0] switch_io_outData_2; // @[Switch.scala 50:22:@617.4]
  wire [47:0] switch_io_outData_3; // @[Switch.scala 50:22:@617.4]
  wire [47:0] switch_io_outData_4; // @[Switch.scala 50:22:@617.4]
  wire [47:0] switch_io_outData_5; // @[Switch.scala 50:22:@617.4]
  wire [47:0] switch_io_outData_6; // @[Switch.scala 50:22:@617.4]
  wire [47:0] switch_io_outData_7; // @[Switch.scala 50:22:@617.4]
  wire  switch_io_outValid_0; // @[Switch.scala 50:22:@617.4]
  wire  switch_io_outValid_1; // @[Switch.scala 50:22:@617.4]
  wire  switch_io_outValid_2; // @[Switch.scala 50:22:@617.4]
  wire  switch_io_outValid_3; // @[Switch.scala 50:22:@617.4]
  wire  switch_io_outValid_4; // @[Switch.scala 50:22:@617.4]
  wire  switch_io_outValid_5; // @[Switch.scala 50:22:@617.4]
  wire  switch_io_outValid_6; // @[Switch.scala 50:22:@617.4]
  wire  switch_io_outValid_7; // @[Switch.scala 50:22:@617.4]
  reg [2:0] _T_102_0; // @[Switch.scala 51:30:@620.4]
  reg [31:0] _RAND_0;
  reg [2:0] _T_102_1; // @[Switch.scala 51:30:@620.4]
  reg [31:0] _RAND_1;
  reg [2:0] _T_102_2; // @[Switch.scala 51:30:@620.4]
  reg [31:0] _RAND_2;
  reg [2:0] _T_102_3; // @[Switch.scala 51:30:@620.4]
  reg [31:0] _RAND_3;
  reg [2:0] _T_102_4; // @[Switch.scala 51:30:@620.4]
  reg [31:0] _RAND_4;
  reg [2:0] _T_102_5; // @[Switch.scala 51:30:@620.4]
  reg [31:0] _RAND_5;
  reg [2:0] _T_102_6; // @[Switch.scala 51:30:@620.4]
  reg [31:0] _RAND_6;
  reg [2:0] _T_102_7; // @[Switch.scala 51:30:@620.4]
  reg [31:0] _RAND_7;
  reg [47:0] _T_151_0; // @[Switch.scala 52:30:@637.4]
  reg [63:0] _RAND_8;
  reg [47:0] _T_151_1; // @[Switch.scala 52:30:@637.4]
  reg [63:0] _RAND_9;
  reg [47:0] _T_151_2; // @[Switch.scala 52:30:@637.4]
  reg [63:0] _RAND_10;
  reg [47:0] _T_151_3; // @[Switch.scala 52:30:@637.4]
  reg [63:0] _RAND_11;
  reg [47:0] _T_151_4; // @[Switch.scala 52:30:@637.4]
  reg [63:0] _RAND_12;
  reg [47:0] _T_151_5; // @[Switch.scala 52:30:@637.4]
  reg [63:0] _RAND_13;
  reg [47:0] _T_151_6; // @[Switch.scala 52:30:@637.4]
  reg [63:0] _RAND_14;
  reg [47:0] _T_151_7; // @[Switch.scala 52:30:@637.4]
  reg [63:0] _RAND_15;
  reg  _T_200_0; // @[Switch.scala 53:31:@654.4]
  reg [31:0] _RAND_16;
  reg  _T_200_1; // @[Switch.scala 53:31:@654.4]
  reg [31:0] _RAND_17;
  reg  _T_200_2; // @[Switch.scala 53:31:@654.4]
  reg [31:0] _RAND_18;
  reg  _T_200_3; // @[Switch.scala 53:31:@654.4]
  reg [31:0] _RAND_19;
  reg  _T_200_4; // @[Switch.scala 53:31:@654.4]
  reg [31:0] _RAND_20;
  reg  _T_200_5; // @[Switch.scala 53:31:@654.4]
  reg [31:0] _RAND_21;
  reg  _T_200_6; // @[Switch.scala 53:31:@654.4]
  reg [31:0] _RAND_22;
  reg  _T_200_7; // @[Switch.scala 53:31:@654.4]
  reg [31:0] _RAND_23;
  reg  _T_249_0; // @[Switch.scala 54:23:@671.4]
  reg [31:0] _RAND_24;
  reg  _T_249_1; // @[Switch.scala 54:23:@671.4]
  reg [31:0] _RAND_25;
  reg  _T_249_2; // @[Switch.scala 54:23:@671.4]
  reg [31:0] _RAND_26;
  reg  _T_249_3; // @[Switch.scala 54:23:@671.4]
  reg [31:0] _RAND_27;
  reg  _T_249_4; // @[Switch.scala 54:23:@671.4]
  reg [31:0] _RAND_28;
  reg  _T_249_5; // @[Switch.scala 54:23:@671.4]
  reg [31:0] _RAND_29;
  reg  _T_249_6; // @[Switch.scala 54:23:@671.4]
  reg [31:0] _RAND_30;
  reg  _T_249_7; // @[Switch.scala 54:23:@671.4]
  reg [31:0] _RAND_31;
  reg [47:0] _T_298_0; // @[Switch.scala 55:24:@688.4]
  reg [63:0] _RAND_32;
  reg [47:0] _T_298_1; // @[Switch.scala 55:24:@688.4]
  reg [63:0] _RAND_33;
  reg [47:0] _T_298_2; // @[Switch.scala 55:24:@688.4]
  reg [63:0] _RAND_34;
  reg [47:0] _T_298_3; // @[Switch.scala 55:24:@688.4]
  reg [63:0] _RAND_35;
  reg [47:0] _T_298_4; // @[Switch.scala 55:24:@688.4]
  reg [63:0] _RAND_36;
  reg [47:0] _T_298_5; // @[Switch.scala 55:24:@688.4]
  reg [63:0] _RAND_37;
  reg [47:0] _T_298_6; // @[Switch.scala 55:24:@688.4]
  reg [63:0] _RAND_38;
  reg [47:0] _T_298_7; // @[Switch.scala 55:24:@688.4]
  reg [63:0] _RAND_39;
  reg  _T_347_0; // @[Switch.scala 56:25:@705.4]
  reg [31:0] _RAND_40;
  reg  _T_347_1; // @[Switch.scala 56:25:@705.4]
  reg [31:0] _RAND_41;
  reg  _T_347_2; // @[Switch.scala 56:25:@705.4]
  reg [31:0] _RAND_42;
  reg  _T_347_3; // @[Switch.scala 56:25:@705.4]
  reg [31:0] _RAND_43;
  reg  _T_347_4; // @[Switch.scala 56:25:@705.4]
  reg [31:0] _RAND_44;
  reg  _T_347_5; // @[Switch.scala 56:25:@705.4]
  reg [31:0] _RAND_45;
  reg  _T_347_6; // @[Switch.scala 56:25:@705.4]
  reg [31:0] _RAND_46;
  reg  _T_347_7; // @[Switch.scala 56:25:@705.4]
  reg [31:0] _RAND_47;
  Switch switch ( // @[Switch.scala 50:22:@617.4]
    .io_inAddr_0(switch_io_inAddr_0),
    .io_inAddr_1(switch_io_inAddr_1),
    .io_inAddr_2(switch_io_inAddr_2),
    .io_inAddr_3(switch_io_inAddr_3),
    .io_inAddr_4(switch_io_inAddr_4),
    .io_inAddr_5(switch_io_inAddr_5),
    .io_inAddr_6(switch_io_inAddr_6),
    .io_inAddr_7(switch_io_inAddr_7),
    .io_inData_0(switch_io_inData_0),
    .io_inData_1(switch_io_inData_1),
    .io_inData_2(switch_io_inData_2),
    .io_inData_3(switch_io_inData_3),
    .io_inData_4(switch_io_inData_4),
    .io_inData_5(switch_io_inData_5),
    .io_inData_6(switch_io_inData_6),
    .io_inData_7(switch_io_inData_7),
    .io_inValid_0(switch_io_inValid_0),
    .io_inValid_1(switch_io_inValid_1),
    .io_inValid_2(switch_io_inValid_2),
    .io_inValid_3(switch_io_inValid_3),
    .io_inValid_4(switch_io_inValid_4),
    .io_inValid_5(switch_io_inValid_5),
    .io_inValid_6(switch_io_inValid_6),
    .io_inValid_7(switch_io_inValid_7),
    .io_outAck_0(switch_io_outAck_0),
    .io_outAck_1(switch_io_outAck_1),
    .io_outAck_2(switch_io_outAck_2),
    .io_outAck_3(switch_io_outAck_3),
    .io_outAck_4(switch_io_outAck_4),
    .io_outAck_5(switch_io_outAck_5),
    .io_outAck_6(switch_io_outAck_6),
    .io_outAck_7(switch_io_outAck_7),
    .io_outData_0(switch_io_outData_0),
    .io_outData_1(switch_io_outData_1),
    .io_outData_2(switch_io_outData_2),
    .io_outData_3(switch_io_outData_3),
    .io_outData_4(switch_io_outData_4),
    .io_outData_5(switch_io_outData_5),
    .io_outData_6(switch_io_outData_6),
    .io_outData_7(switch_io_outData_7),
    .io_outValid_0(switch_io_outValid_0),
    .io_outValid_1(switch_io_outValid_1),
    .io_outValid_2(switch_io_outValid_2),
    .io_outValid_3(switch_io_outValid_3),
    .io_outValid_4(switch_io_outValid_4),
    .io_outValid_5(switch_io_outValid_5),
    .io_outValid_6(switch_io_outValid_6),
    .io_outValid_7(switch_io_outValid_7)
  );
  assign io_outAck_0 = _T_249_0; // @[Switch.scala 54:13:@680.4]
  assign io_outAck_1 = _T_249_1; // @[Switch.scala 54:13:@681.4]
  assign io_outAck_2 = _T_249_2; // @[Switch.scala 54:13:@682.4]
  assign io_outAck_3 = _T_249_3; // @[Switch.scala 54:13:@683.4]
  assign io_outAck_4 = _T_249_4; // @[Switch.scala 54:13:@684.4]
  assign io_outAck_5 = _T_249_5; // @[Switch.scala 54:13:@685.4]
  assign io_outAck_6 = _T_249_6; // @[Switch.scala 54:13:@686.4]
  assign io_outAck_7 = _T_249_7; // @[Switch.scala 54:13:@687.4]
  assign io_outData_0 = _T_298_0; // @[Switch.scala 55:14:@697.4]
  assign io_outData_1 = _T_298_1; // @[Switch.scala 55:14:@698.4]
  assign io_outData_2 = _T_298_2; // @[Switch.scala 55:14:@699.4]
  assign io_outData_3 = _T_298_3; // @[Switch.scala 55:14:@700.4]
  assign io_outData_4 = _T_298_4; // @[Switch.scala 55:14:@701.4]
  assign io_outData_5 = _T_298_5; // @[Switch.scala 55:14:@702.4]
  assign io_outData_6 = _T_298_6; // @[Switch.scala 55:14:@703.4]
  assign io_outData_7 = _T_298_7; // @[Switch.scala 55:14:@704.4]
  assign io_outValid_0 = _T_347_0; // @[Switch.scala 56:15:@714.4]
  assign io_outValid_1 = _T_347_1; // @[Switch.scala 56:15:@715.4]
  assign io_outValid_2 = _T_347_2; // @[Switch.scala 56:15:@716.4]
  assign io_outValid_3 = _T_347_3; // @[Switch.scala 56:15:@717.4]
  assign io_outValid_4 = _T_347_4; // @[Switch.scala 56:15:@718.4]
  assign io_outValid_5 = _T_347_5; // @[Switch.scala 56:15:@719.4]
  assign io_outValid_6 = _T_347_6; // @[Switch.scala 56:15:@720.4]
  assign io_outValid_7 = _T_347_7; // @[Switch.scala 56:15:@721.4]
  assign switch_io_inAddr_0 = _T_102_0; // @[Switch.scala 51:20:@629.4]
  assign switch_io_inAddr_1 = _T_102_1; // @[Switch.scala 51:20:@630.4]
  assign switch_io_inAddr_2 = _T_102_2; // @[Switch.scala 51:20:@631.4]
  assign switch_io_inAddr_3 = _T_102_3; // @[Switch.scala 51:20:@632.4]
  assign switch_io_inAddr_4 = _T_102_4; // @[Switch.scala 51:20:@633.4]
  assign switch_io_inAddr_5 = _T_102_5; // @[Switch.scala 51:20:@634.4]
  assign switch_io_inAddr_6 = _T_102_6; // @[Switch.scala 51:20:@635.4]
  assign switch_io_inAddr_7 = _T_102_7; // @[Switch.scala 51:20:@636.4]
  assign switch_io_inData_0 = _T_151_0; // @[Switch.scala 52:20:@646.4]
  assign switch_io_inData_1 = _T_151_1; // @[Switch.scala 52:20:@647.4]
  assign switch_io_inData_2 = _T_151_2; // @[Switch.scala 52:20:@648.4]
  assign switch_io_inData_3 = _T_151_3; // @[Switch.scala 52:20:@649.4]
  assign switch_io_inData_4 = _T_151_4; // @[Switch.scala 52:20:@650.4]
  assign switch_io_inData_5 = _T_151_5; // @[Switch.scala 52:20:@651.4]
  assign switch_io_inData_6 = _T_151_6; // @[Switch.scala 52:20:@652.4]
  assign switch_io_inData_7 = _T_151_7; // @[Switch.scala 52:20:@653.4]
  assign switch_io_inValid_0 = _T_200_0; // @[Switch.scala 53:21:@663.4]
  assign switch_io_inValid_1 = _T_200_1; // @[Switch.scala 53:21:@664.4]
  assign switch_io_inValid_2 = _T_200_2; // @[Switch.scala 53:21:@665.4]
  assign switch_io_inValid_3 = _T_200_3; // @[Switch.scala 53:21:@666.4]
  assign switch_io_inValid_4 = _T_200_4; // @[Switch.scala 53:21:@667.4]
  assign switch_io_inValid_5 = _T_200_5; // @[Switch.scala 53:21:@668.4]
  assign switch_io_inValid_6 = _T_200_6; // @[Switch.scala 53:21:@669.4]
  assign switch_io_inValid_7 = _T_200_7; // @[Switch.scala 53:21:@670.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_102_0 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_102_1 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_102_2 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_102_3 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_102_4 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_102_5 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_102_6 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_102_7 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {2{`RANDOM}};
  _T_151_0 = _RAND_8[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {2{`RANDOM}};
  _T_151_1 = _RAND_9[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {2{`RANDOM}};
  _T_151_2 = _RAND_10[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {2{`RANDOM}};
  _T_151_3 = _RAND_11[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {2{`RANDOM}};
  _T_151_4 = _RAND_12[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {2{`RANDOM}};
  _T_151_5 = _RAND_13[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {2{`RANDOM}};
  _T_151_6 = _RAND_14[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {2{`RANDOM}};
  _T_151_7 = _RAND_15[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_200_0 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_200_1 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_200_2 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_200_3 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_200_4 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_200_5 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_200_6 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_200_7 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_249_0 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_249_1 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_249_2 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_249_3 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_249_4 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_249_5 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_249_6 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_249_7 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {2{`RANDOM}};
  _T_298_0 = _RAND_32[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {2{`RANDOM}};
  _T_298_1 = _RAND_33[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {2{`RANDOM}};
  _T_298_2 = _RAND_34[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {2{`RANDOM}};
  _T_298_3 = _RAND_35[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {2{`RANDOM}};
  _T_298_4 = _RAND_36[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {2{`RANDOM}};
  _T_298_5 = _RAND_37[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {2{`RANDOM}};
  _T_298_6 = _RAND_38[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {2{`RANDOM}};
  _T_298_7 = _RAND_39[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_347_0 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_347_1 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_347_2 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_347_3 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_347_4 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_347_5 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_347_6 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_347_7 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    _T_102_0 <= io_inAddr_0;
    _T_102_1 <= io_inAddr_1;
    _T_102_2 <= io_inAddr_2;
    _T_102_3 <= io_inAddr_3;
    _T_102_4 <= io_inAddr_4;
    _T_102_5 <= io_inAddr_5;
    _T_102_6 <= io_inAddr_6;
    _T_102_7 <= io_inAddr_7;
    _T_151_0 <= io_inData_0;
    _T_151_1 <= io_inData_1;
    _T_151_2 <= io_inData_2;
    _T_151_3 <= io_inData_3;
    _T_151_4 <= io_inData_4;
    _T_151_5 <= io_inData_5;
    _T_151_6 <= io_inData_6;
    _T_151_7 <= io_inData_7;
    _T_200_0 <= io_inValid_0;
    _T_200_1 <= io_inValid_1;
    _T_200_2 <= io_inValid_2;
    _T_200_3 <= io_inValid_3;
    _T_200_4 <= io_inValid_4;
    _T_200_5 <= io_inValid_5;
    _T_200_6 <= io_inValid_6;
    _T_200_7 <= io_inValid_7;
    _T_249_0 <= switch_io_outAck_0;
    _T_249_1 <= switch_io_outAck_1;
    _T_249_2 <= switch_io_outAck_2;
    _T_249_3 <= switch_io_outAck_3;
    _T_249_4 <= switch_io_outAck_4;
    _T_249_5 <= switch_io_outAck_5;
    _T_249_6 <= switch_io_outAck_6;
    _T_249_7 <= switch_io_outAck_7;
    _T_298_0 <= switch_io_outData_0;
    _T_298_1 <= switch_io_outData_1;
    _T_298_2 <= switch_io_outData_2;
    _T_298_3 <= switch_io_outData_3;
    _T_298_4 <= switch_io_outData_4;
    _T_298_5 <= switch_io_outData_5;
    _T_298_6 <= switch_io_outData_6;
    _T_298_7 <= switch_io_outData_7;
    _T_347_0 <= switch_io_outValid_0;
    _T_347_1 <= switch_io_outValid_1;
    _T_347_2 <= switch_io_outValid_2;
    _T_347_3 <= switch_io_outValid_3;
    _T_347_4 <= switch_io_outValid_4;
    _T_347_5 <= switch_io_outValid_5;
    _T_347_6 <= switch_io_outValid_6;
    _T_347_7 <= switch_io_outValid_7;
  end
endmodule
