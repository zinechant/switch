module Switch( // @[:@3.2]
  input  [4:0]  io_inAddr_0, // @[:@6.4]
  input  [4:0]  io_inAddr_1, // @[:@6.4]
  input  [4:0]  io_inAddr_2, // @[:@6.4]
  input  [4:0]  io_inAddr_3, // @[:@6.4]
  input  [4:0]  io_inAddr_4, // @[:@6.4]
  input  [4:0]  io_inAddr_5, // @[:@6.4]
  input  [4:0]  io_inAddr_6, // @[:@6.4]
  input  [4:0]  io_inAddr_7, // @[:@6.4]
  input  [4:0]  io_inAddr_8, // @[:@6.4]
  input  [4:0]  io_inAddr_9, // @[:@6.4]
  input  [4:0]  io_inAddr_10, // @[:@6.4]
  input  [4:0]  io_inAddr_11, // @[:@6.4]
  input  [4:0]  io_inAddr_12, // @[:@6.4]
  input  [4:0]  io_inAddr_13, // @[:@6.4]
  input  [4:0]  io_inAddr_14, // @[:@6.4]
  input  [4:0]  io_inAddr_15, // @[:@6.4]
  input  [4:0]  io_inAddr_16, // @[:@6.4]
  input  [4:0]  io_inAddr_17, // @[:@6.4]
  input  [4:0]  io_inAddr_18, // @[:@6.4]
  input  [4:0]  io_inAddr_19, // @[:@6.4]
  input  [4:0]  io_inAddr_20, // @[:@6.4]
  input  [4:0]  io_inAddr_21, // @[:@6.4]
  input  [4:0]  io_inAddr_22, // @[:@6.4]
  input  [4:0]  io_inAddr_23, // @[:@6.4]
  input  [4:0]  io_inAddr_24, // @[:@6.4]
  input  [4:0]  io_inAddr_25, // @[:@6.4]
  input  [4:0]  io_inAddr_26, // @[:@6.4]
  input  [4:0]  io_inAddr_27, // @[:@6.4]
  input  [4:0]  io_inAddr_28, // @[:@6.4]
  input  [4:0]  io_inAddr_29, // @[:@6.4]
  input  [4:0]  io_inAddr_30, // @[:@6.4]
  input  [4:0]  io_inAddr_31, // @[:@6.4]
  input  [47:0] io_inData_0, // @[:@6.4]
  input  [47:0] io_inData_1, // @[:@6.4]
  input  [47:0] io_inData_2, // @[:@6.4]
  input  [47:0] io_inData_3, // @[:@6.4]
  input  [47:0] io_inData_4, // @[:@6.4]
  input  [47:0] io_inData_5, // @[:@6.4]
  input  [47:0] io_inData_6, // @[:@6.4]
  input  [47:0] io_inData_7, // @[:@6.4]
  input  [47:0] io_inData_8, // @[:@6.4]
  input  [47:0] io_inData_9, // @[:@6.4]
  input  [47:0] io_inData_10, // @[:@6.4]
  input  [47:0] io_inData_11, // @[:@6.4]
  input  [47:0] io_inData_12, // @[:@6.4]
  input  [47:0] io_inData_13, // @[:@6.4]
  input  [47:0] io_inData_14, // @[:@6.4]
  input  [47:0] io_inData_15, // @[:@6.4]
  input  [47:0] io_inData_16, // @[:@6.4]
  input  [47:0] io_inData_17, // @[:@6.4]
  input  [47:0] io_inData_18, // @[:@6.4]
  input  [47:0] io_inData_19, // @[:@6.4]
  input  [47:0] io_inData_20, // @[:@6.4]
  input  [47:0] io_inData_21, // @[:@6.4]
  input  [47:0] io_inData_22, // @[:@6.4]
  input  [47:0] io_inData_23, // @[:@6.4]
  input  [47:0] io_inData_24, // @[:@6.4]
  input  [47:0] io_inData_25, // @[:@6.4]
  input  [47:0] io_inData_26, // @[:@6.4]
  input  [47:0] io_inData_27, // @[:@6.4]
  input  [47:0] io_inData_28, // @[:@6.4]
  input  [47:0] io_inData_29, // @[:@6.4]
  input  [47:0] io_inData_30, // @[:@6.4]
  input  [47:0] io_inData_31, // @[:@6.4]
  input         io_inValid_0, // @[:@6.4]
  input         io_inValid_1, // @[:@6.4]
  input         io_inValid_2, // @[:@6.4]
  input         io_inValid_3, // @[:@6.4]
  input         io_inValid_4, // @[:@6.4]
  input         io_inValid_5, // @[:@6.4]
  input         io_inValid_6, // @[:@6.4]
  input         io_inValid_7, // @[:@6.4]
  input         io_inValid_8, // @[:@6.4]
  input         io_inValid_9, // @[:@6.4]
  input         io_inValid_10, // @[:@6.4]
  input         io_inValid_11, // @[:@6.4]
  input         io_inValid_12, // @[:@6.4]
  input         io_inValid_13, // @[:@6.4]
  input         io_inValid_14, // @[:@6.4]
  input         io_inValid_15, // @[:@6.4]
  input         io_inValid_16, // @[:@6.4]
  input         io_inValid_17, // @[:@6.4]
  input         io_inValid_18, // @[:@6.4]
  input         io_inValid_19, // @[:@6.4]
  input         io_inValid_20, // @[:@6.4]
  input         io_inValid_21, // @[:@6.4]
  input         io_inValid_22, // @[:@6.4]
  input         io_inValid_23, // @[:@6.4]
  input         io_inValid_24, // @[:@6.4]
  input         io_inValid_25, // @[:@6.4]
  input         io_inValid_26, // @[:@6.4]
  input         io_inValid_27, // @[:@6.4]
  input         io_inValid_28, // @[:@6.4]
  input         io_inValid_29, // @[:@6.4]
  input         io_inValid_30, // @[:@6.4]
  input         io_inValid_31, // @[:@6.4]
  output        io_outAck_0, // @[:@6.4]
  output        io_outAck_1, // @[:@6.4]
  output        io_outAck_2, // @[:@6.4]
  output        io_outAck_3, // @[:@6.4]
  output        io_outAck_4, // @[:@6.4]
  output        io_outAck_5, // @[:@6.4]
  output        io_outAck_6, // @[:@6.4]
  output        io_outAck_7, // @[:@6.4]
  output        io_outAck_8, // @[:@6.4]
  output        io_outAck_9, // @[:@6.4]
  output        io_outAck_10, // @[:@6.4]
  output        io_outAck_11, // @[:@6.4]
  output        io_outAck_12, // @[:@6.4]
  output        io_outAck_13, // @[:@6.4]
  output        io_outAck_14, // @[:@6.4]
  output        io_outAck_15, // @[:@6.4]
  output        io_outAck_16, // @[:@6.4]
  output        io_outAck_17, // @[:@6.4]
  output        io_outAck_18, // @[:@6.4]
  output        io_outAck_19, // @[:@6.4]
  output        io_outAck_20, // @[:@6.4]
  output        io_outAck_21, // @[:@6.4]
  output        io_outAck_22, // @[:@6.4]
  output        io_outAck_23, // @[:@6.4]
  output        io_outAck_24, // @[:@6.4]
  output        io_outAck_25, // @[:@6.4]
  output        io_outAck_26, // @[:@6.4]
  output        io_outAck_27, // @[:@6.4]
  output        io_outAck_28, // @[:@6.4]
  output        io_outAck_29, // @[:@6.4]
  output        io_outAck_30, // @[:@6.4]
  output        io_outAck_31, // @[:@6.4]
  output [47:0] io_outData_0, // @[:@6.4]
  output [47:0] io_outData_1, // @[:@6.4]
  output [47:0] io_outData_2, // @[:@6.4]
  output [47:0] io_outData_3, // @[:@6.4]
  output [47:0] io_outData_4, // @[:@6.4]
  output [47:0] io_outData_5, // @[:@6.4]
  output [47:0] io_outData_6, // @[:@6.4]
  output [47:0] io_outData_7, // @[:@6.4]
  output [47:0] io_outData_8, // @[:@6.4]
  output [47:0] io_outData_9, // @[:@6.4]
  output [47:0] io_outData_10, // @[:@6.4]
  output [47:0] io_outData_11, // @[:@6.4]
  output [47:0] io_outData_12, // @[:@6.4]
  output [47:0] io_outData_13, // @[:@6.4]
  output [47:0] io_outData_14, // @[:@6.4]
  output [47:0] io_outData_15, // @[:@6.4]
  output [47:0] io_outData_16, // @[:@6.4]
  output [47:0] io_outData_17, // @[:@6.4]
  output [47:0] io_outData_18, // @[:@6.4]
  output [47:0] io_outData_19, // @[:@6.4]
  output [47:0] io_outData_20, // @[:@6.4]
  output [47:0] io_outData_21, // @[:@6.4]
  output [47:0] io_outData_22, // @[:@6.4]
  output [47:0] io_outData_23, // @[:@6.4]
  output [47:0] io_outData_24, // @[:@6.4]
  output [47:0] io_outData_25, // @[:@6.4]
  output [47:0] io_outData_26, // @[:@6.4]
  output [47:0] io_outData_27, // @[:@6.4]
  output [47:0] io_outData_28, // @[:@6.4]
  output [47:0] io_outData_29, // @[:@6.4]
  output [47:0] io_outData_30, // @[:@6.4]
  output [47:0] io_outData_31, // @[:@6.4]
  output        io_outValid_0, // @[:@6.4]
  output        io_outValid_1, // @[:@6.4]
  output        io_outValid_2, // @[:@6.4]
  output        io_outValid_3, // @[:@6.4]
  output        io_outValid_4, // @[:@6.4]
  output        io_outValid_5, // @[:@6.4]
  output        io_outValid_6, // @[:@6.4]
  output        io_outValid_7, // @[:@6.4]
  output        io_outValid_8, // @[:@6.4]
  output        io_outValid_9, // @[:@6.4]
  output        io_outValid_10, // @[:@6.4]
  output        io_outValid_11, // @[:@6.4]
  output        io_outValid_12, // @[:@6.4]
  output        io_outValid_13, // @[:@6.4]
  output        io_outValid_14, // @[:@6.4]
  output        io_outValid_15, // @[:@6.4]
  output        io_outValid_16, // @[:@6.4]
  output        io_outValid_17, // @[:@6.4]
  output        io_outValid_18, // @[:@6.4]
  output        io_outValid_19, // @[:@6.4]
  output        io_outValid_20, // @[:@6.4]
  output        io_outValid_21, // @[:@6.4]
  output        io_outValid_22, // @[:@6.4]
  output        io_outValid_23, // @[:@6.4]
  output        io_outValid_24, // @[:@6.4]
  output        io_outValid_25, // @[:@6.4]
  output        io_outValid_26, // @[:@6.4]
  output        io_outValid_27, // @[:@6.4]
  output        io_outValid_28, // @[:@6.4]
  output        io_outValid_29, // @[:@6.4]
  output        io_outValid_30, // @[:@6.4]
  output        io_outValid_31 // @[:@6.4]
);
  wire  _T_4758; // @[Switch.scala 30:53:@10.4]
  wire  valid_0_0; // @[Switch.scala 30:36:@11.4]
  wire  _T_4761; // @[Switch.scala 30:53:@13.4]
  wire  valid_0_1; // @[Switch.scala 30:36:@14.4]
  wire  _T_4764; // @[Switch.scala 30:53:@16.4]
  wire  valid_0_2; // @[Switch.scala 30:36:@17.4]
  wire  _T_4767; // @[Switch.scala 30:53:@19.4]
  wire  valid_0_3; // @[Switch.scala 30:36:@20.4]
  wire  _T_4770; // @[Switch.scala 30:53:@22.4]
  wire  valid_0_4; // @[Switch.scala 30:36:@23.4]
  wire  _T_4773; // @[Switch.scala 30:53:@25.4]
  wire  valid_0_5; // @[Switch.scala 30:36:@26.4]
  wire  _T_4776; // @[Switch.scala 30:53:@28.4]
  wire  valid_0_6; // @[Switch.scala 30:36:@29.4]
  wire  _T_4779; // @[Switch.scala 30:53:@31.4]
  wire  valid_0_7; // @[Switch.scala 30:36:@32.4]
  wire  _T_4782; // @[Switch.scala 30:53:@34.4]
  wire  valid_0_8; // @[Switch.scala 30:36:@35.4]
  wire  _T_4785; // @[Switch.scala 30:53:@37.4]
  wire  valid_0_9; // @[Switch.scala 30:36:@38.4]
  wire  _T_4788; // @[Switch.scala 30:53:@40.4]
  wire  valid_0_10; // @[Switch.scala 30:36:@41.4]
  wire  _T_4791; // @[Switch.scala 30:53:@43.4]
  wire  valid_0_11; // @[Switch.scala 30:36:@44.4]
  wire  _T_4794; // @[Switch.scala 30:53:@46.4]
  wire  valid_0_12; // @[Switch.scala 30:36:@47.4]
  wire  _T_4797; // @[Switch.scala 30:53:@49.4]
  wire  valid_0_13; // @[Switch.scala 30:36:@50.4]
  wire  _T_4800; // @[Switch.scala 30:53:@52.4]
  wire  valid_0_14; // @[Switch.scala 30:36:@53.4]
  wire  _T_4803; // @[Switch.scala 30:53:@55.4]
  wire  valid_0_15; // @[Switch.scala 30:36:@56.4]
  wire  _T_4806; // @[Switch.scala 30:53:@58.4]
  wire  valid_0_16; // @[Switch.scala 30:36:@59.4]
  wire  _T_4809; // @[Switch.scala 30:53:@61.4]
  wire  valid_0_17; // @[Switch.scala 30:36:@62.4]
  wire  _T_4812; // @[Switch.scala 30:53:@64.4]
  wire  valid_0_18; // @[Switch.scala 30:36:@65.4]
  wire  _T_4815; // @[Switch.scala 30:53:@67.4]
  wire  valid_0_19; // @[Switch.scala 30:36:@68.4]
  wire  _T_4818; // @[Switch.scala 30:53:@70.4]
  wire  valid_0_20; // @[Switch.scala 30:36:@71.4]
  wire  _T_4821; // @[Switch.scala 30:53:@73.4]
  wire  valid_0_21; // @[Switch.scala 30:36:@74.4]
  wire  _T_4824; // @[Switch.scala 30:53:@76.4]
  wire  valid_0_22; // @[Switch.scala 30:36:@77.4]
  wire  _T_4827; // @[Switch.scala 30:53:@79.4]
  wire  valid_0_23; // @[Switch.scala 30:36:@80.4]
  wire  _T_4830; // @[Switch.scala 30:53:@82.4]
  wire  valid_0_24; // @[Switch.scala 30:36:@83.4]
  wire  _T_4833; // @[Switch.scala 30:53:@85.4]
  wire  valid_0_25; // @[Switch.scala 30:36:@86.4]
  wire  _T_4836; // @[Switch.scala 30:53:@88.4]
  wire  valid_0_26; // @[Switch.scala 30:36:@89.4]
  wire  _T_4839; // @[Switch.scala 30:53:@91.4]
  wire  valid_0_27; // @[Switch.scala 30:36:@92.4]
  wire  _T_4842; // @[Switch.scala 30:53:@94.4]
  wire  valid_0_28; // @[Switch.scala 30:36:@95.4]
  wire  _T_4845; // @[Switch.scala 30:53:@97.4]
  wire  valid_0_29; // @[Switch.scala 30:36:@98.4]
  wire  _T_4848; // @[Switch.scala 30:53:@100.4]
  wire  valid_0_30; // @[Switch.scala 30:36:@101.4]
  wire  _T_4851; // @[Switch.scala 30:53:@103.4]
  wire  valid_0_31; // @[Switch.scala 30:36:@104.4]
  wire [4:0] _T_4885; // @[Mux.scala 31:69:@106.4]
  wire [4:0] _T_4886; // @[Mux.scala 31:69:@107.4]
  wire [4:0] _T_4887; // @[Mux.scala 31:69:@108.4]
  wire [4:0] _T_4888; // @[Mux.scala 31:69:@109.4]
  wire [4:0] _T_4889; // @[Mux.scala 31:69:@110.4]
  wire [4:0] _T_4890; // @[Mux.scala 31:69:@111.4]
  wire [4:0] _T_4891; // @[Mux.scala 31:69:@112.4]
  wire [4:0] _T_4892; // @[Mux.scala 31:69:@113.4]
  wire [4:0] _T_4893; // @[Mux.scala 31:69:@114.4]
  wire [4:0] _T_4894; // @[Mux.scala 31:69:@115.4]
  wire [4:0] _T_4895; // @[Mux.scala 31:69:@116.4]
  wire [4:0] _T_4896; // @[Mux.scala 31:69:@117.4]
  wire [4:0] _T_4897; // @[Mux.scala 31:69:@118.4]
  wire [4:0] _T_4898; // @[Mux.scala 31:69:@119.4]
  wire [4:0] _T_4899; // @[Mux.scala 31:69:@120.4]
  wire [4:0] _T_4900; // @[Mux.scala 31:69:@121.4]
  wire [4:0] _T_4901; // @[Mux.scala 31:69:@122.4]
  wire [4:0] _T_4902; // @[Mux.scala 31:69:@123.4]
  wire [4:0] _T_4903; // @[Mux.scala 31:69:@124.4]
  wire [4:0] _T_4904; // @[Mux.scala 31:69:@125.4]
  wire [4:0] _T_4905; // @[Mux.scala 31:69:@126.4]
  wire [4:0] _T_4906; // @[Mux.scala 31:69:@127.4]
  wire [4:0] _T_4907; // @[Mux.scala 31:69:@128.4]
  wire [4:0] _T_4908; // @[Mux.scala 31:69:@129.4]
  wire [4:0] _T_4909; // @[Mux.scala 31:69:@130.4]
  wire [4:0] _T_4910; // @[Mux.scala 31:69:@131.4]
  wire [4:0] _T_4911; // @[Mux.scala 31:69:@132.4]
  wire [4:0] _T_4912; // @[Mux.scala 31:69:@133.4]
  wire [4:0] _T_4913; // @[Mux.scala 31:69:@134.4]
  wire [4:0] _T_4914; // @[Mux.scala 31:69:@135.4]
  wire [4:0] select_0; // @[Mux.scala 31:69:@136.4]
  wire [47:0] _GEN_1; // @[Switch.scala 33:19:@138.4]
  wire [47:0] _GEN_2; // @[Switch.scala 33:19:@138.4]
  wire [47:0] _GEN_3; // @[Switch.scala 33:19:@138.4]
  wire [47:0] _GEN_4; // @[Switch.scala 33:19:@138.4]
  wire [47:0] _GEN_5; // @[Switch.scala 33:19:@138.4]
  wire [47:0] _GEN_6; // @[Switch.scala 33:19:@138.4]
  wire [47:0] _GEN_7; // @[Switch.scala 33:19:@138.4]
  wire [47:0] _GEN_8; // @[Switch.scala 33:19:@138.4]
  wire [47:0] _GEN_9; // @[Switch.scala 33:19:@138.4]
  wire [47:0] _GEN_10; // @[Switch.scala 33:19:@138.4]
  wire [47:0] _GEN_11; // @[Switch.scala 33:19:@138.4]
  wire [47:0] _GEN_12; // @[Switch.scala 33:19:@138.4]
  wire [47:0] _GEN_13; // @[Switch.scala 33:19:@138.4]
  wire [47:0] _GEN_14; // @[Switch.scala 33:19:@138.4]
  wire [47:0] _GEN_15; // @[Switch.scala 33:19:@138.4]
  wire [47:0] _GEN_16; // @[Switch.scala 33:19:@138.4]
  wire [47:0] _GEN_17; // @[Switch.scala 33:19:@138.4]
  wire [47:0] _GEN_18; // @[Switch.scala 33:19:@138.4]
  wire [47:0] _GEN_19; // @[Switch.scala 33:19:@138.4]
  wire [47:0] _GEN_20; // @[Switch.scala 33:19:@138.4]
  wire [47:0] _GEN_21; // @[Switch.scala 33:19:@138.4]
  wire [47:0] _GEN_22; // @[Switch.scala 33:19:@138.4]
  wire [47:0] _GEN_23; // @[Switch.scala 33:19:@138.4]
  wire [47:0] _GEN_24; // @[Switch.scala 33:19:@138.4]
  wire [47:0] _GEN_25; // @[Switch.scala 33:19:@138.4]
  wire [47:0] _GEN_26; // @[Switch.scala 33:19:@138.4]
  wire [47:0] _GEN_27; // @[Switch.scala 33:19:@138.4]
  wire [47:0] _GEN_28; // @[Switch.scala 33:19:@138.4]
  wire [47:0] _GEN_29; // @[Switch.scala 33:19:@138.4]
  wire [47:0] _GEN_30; // @[Switch.scala 33:19:@138.4]
  wire [7:0] _T_4923; // @[Switch.scala 34:32:@145.4]
  wire [15:0] _T_4931; // @[Switch.scala 34:32:@153.4]
  wire [7:0] _T_4938; // @[Switch.scala 34:32:@160.4]
  wire [31:0] _T_4947; // @[Switch.scala 34:32:@169.4]
  wire  _T_4951; // @[Switch.scala 30:53:@172.4]
  wire  valid_1_0; // @[Switch.scala 30:36:@173.4]
  wire  _T_4954; // @[Switch.scala 30:53:@175.4]
  wire  valid_1_1; // @[Switch.scala 30:36:@176.4]
  wire  _T_4957; // @[Switch.scala 30:53:@178.4]
  wire  valid_1_2; // @[Switch.scala 30:36:@179.4]
  wire  _T_4960; // @[Switch.scala 30:53:@181.4]
  wire  valid_1_3; // @[Switch.scala 30:36:@182.4]
  wire  _T_4963; // @[Switch.scala 30:53:@184.4]
  wire  valid_1_4; // @[Switch.scala 30:36:@185.4]
  wire  _T_4966; // @[Switch.scala 30:53:@187.4]
  wire  valid_1_5; // @[Switch.scala 30:36:@188.4]
  wire  _T_4969; // @[Switch.scala 30:53:@190.4]
  wire  valid_1_6; // @[Switch.scala 30:36:@191.4]
  wire  _T_4972; // @[Switch.scala 30:53:@193.4]
  wire  valid_1_7; // @[Switch.scala 30:36:@194.4]
  wire  _T_4975; // @[Switch.scala 30:53:@196.4]
  wire  valid_1_8; // @[Switch.scala 30:36:@197.4]
  wire  _T_4978; // @[Switch.scala 30:53:@199.4]
  wire  valid_1_9; // @[Switch.scala 30:36:@200.4]
  wire  _T_4981; // @[Switch.scala 30:53:@202.4]
  wire  valid_1_10; // @[Switch.scala 30:36:@203.4]
  wire  _T_4984; // @[Switch.scala 30:53:@205.4]
  wire  valid_1_11; // @[Switch.scala 30:36:@206.4]
  wire  _T_4987; // @[Switch.scala 30:53:@208.4]
  wire  valid_1_12; // @[Switch.scala 30:36:@209.4]
  wire  _T_4990; // @[Switch.scala 30:53:@211.4]
  wire  valid_1_13; // @[Switch.scala 30:36:@212.4]
  wire  _T_4993; // @[Switch.scala 30:53:@214.4]
  wire  valid_1_14; // @[Switch.scala 30:36:@215.4]
  wire  _T_4996; // @[Switch.scala 30:53:@217.4]
  wire  valid_1_15; // @[Switch.scala 30:36:@218.4]
  wire  _T_4999; // @[Switch.scala 30:53:@220.4]
  wire  valid_1_16; // @[Switch.scala 30:36:@221.4]
  wire  _T_5002; // @[Switch.scala 30:53:@223.4]
  wire  valid_1_17; // @[Switch.scala 30:36:@224.4]
  wire  _T_5005; // @[Switch.scala 30:53:@226.4]
  wire  valid_1_18; // @[Switch.scala 30:36:@227.4]
  wire  _T_5008; // @[Switch.scala 30:53:@229.4]
  wire  valid_1_19; // @[Switch.scala 30:36:@230.4]
  wire  _T_5011; // @[Switch.scala 30:53:@232.4]
  wire  valid_1_20; // @[Switch.scala 30:36:@233.4]
  wire  _T_5014; // @[Switch.scala 30:53:@235.4]
  wire  valid_1_21; // @[Switch.scala 30:36:@236.4]
  wire  _T_5017; // @[Switch.scala 30:53:@238.4]
  wire  valid_1_22; // @[Switch.scala 30:36:@239.4]
  wire  _T_5020; // @[Switch.scala 30:53:@241.4]
  wire  valid_1_23; // @[Switch.scala 30:36:@242.4]
  wire  _T_5023; // @[Switch.scala 30:53:@244.4]
  wire  valid_1_24; // @[Switch.scala 30:36:@245.4]
  wire  _T_5026; // @[Switch.scala 30:53:@247.4]
  wire  valid_1_25; // @[Switch.scala 30:36:@248.4]
  wire  _T_5029; // @[Switch.scala 30:53:@250.4]
  wire  valid_1_26; // @[Switch.scala 30:36:@251.4]
  wire  _T_5032; // @[Switch.scala 30:53:@253.4]
  wire  valid_1_27; // @[Switch.scala 30:36:@254.4]
  wire  _T_5035; // @[Switch.scala 30:53:@256.4]
  wire  valid_1_28; // @[Switch.scala 30:36:@257.4]
  wire  _T_5038; // @[Switch.scala 30:53:@259.4]
  wire  valid_1_29; // @[Switch.scala 30:36:@260.4]
  wire  _T_5041; // @[Switch.scala 30:53:@262.4]
  wire  valid_1_30; // @[Switch.scala 30:36:@263.4]
  wire  _T_5044; // @[Switch.scala 30:53:@265.4]
  wire  valid_1_31; // @[Switch.scala 30:36:@266.4]
  wire [4:0] _T_5078; // @[Mux.scala 31:69:@268.4]
  wire [4:0] _T_5079; // @[Mux.scala 31:69:@269.4]
  wire [4:0] _T_5080; // @[Mux.scala 31:69:@270.4]
  wire [4:0] _T_5081; // @[Mux.scala 31:69:@271.4]
  wire [4:0] _T_5082; // @[Mux.scala 31:69:@272.4]
  wire [4:0] _T_5083; // @[Mux.scala 31:69:@273.4]
  wire [4:0] _T_5084; // @[Mux.scala 31:69:@274.4]
  wire [4:0] _T_5085; // @[Mux.scala 31:69:@275.4]
  wire [4:0] _T_5086; // @[Mux.scala 31:69:@276.4]
  wire [4:0] _T_5087; // @[Mux.scala 31:69:@277.4]
  wire [4:0] _T_5088; // @[Mux.scala 31:69:@278.4]
  wire [4:0] _T_5089; // @[Mux.scala 31:69:@279.4]
  wire [4:0] _T_5090; // @[Mux.scala 31:69:@280.4]
  wire [4:0] _T_5091; // @[Mux.scala 31:69:@281.4]
  wire [4:0] _T_5092; // @[Mux.scala 31:69:@282.4]
  wire [4:0] _T_5093; // @[Mux.scala 31:69:@283.4]
  wire [4:0] _T_5094; // @[Mux.scala 31:69:@284.4]
  wire [4:0] _T_5095; // @[Mux.scala 31:69:@285.4]
  wire [4:0] _T_5096; // @[Mux.scala 31:69:@286.4]
  wire [4:0] _T_5097; // @[Mux.scala 31:69:@287.4]
  wire [4:0] _T_5098; // @[Mux.scala 31:69:@288.4]
  wire [4:0] _T_5099; // @[Mux.scala 31:69:@289.4]
  wire [4:0] _T_5100; // @[Mux.scala 31:69:@290.4]
  wire [4:0] _T_5101; // @[Mux.scala 31:69:@291.4]
  wire [4:0] _T_5102; // @[Mux.scala 31:69:@292.4]
  wire [4:0] _T_5103; // @[Mux.scala 31:69:@293.4]
  wire [4:0] _T_5104; // @[Mux.scala 31:69:@294.4]
  wire [4:0] _T_5105; // @[Mux.scala 31:69:@295.4]
  wire [4:0] _T_5106; // @[Mux.scala 31:69:@296.4]
  wire [4:0] _T_5107; // @[Mux.scala 31:69:@297.4]
  wire [4:0] select_1; // @[Mux.scala 31:69:@298.4]
  wire [47:0] _GEN_33; // @[Switch.scala 33:19:@300.4]
  wire [47:0] _GEN_34; // @[Switch.scala 33:19:@300.4]
  wire [47:0] _GEN_35; // @[Switch.scala 33:19:@300.4]
  wire [47:0] _GEN_36; // @[Switch.scala 33:19:@300.4]
  wire [47:0] _GEN_37; // @[Switch.scala 33:19:@300.4]
  wire [47:0] _GEN_38; // @[Switch.scala 33:19:@300.4]
  wire [47:0] _GEN_39; // @[Switch.scala 33:19:@300.4]
  wire [47:0] _GEN_40; // @[Switch.scala 33:19:@300.4]
  wire [47:0] _GEN_41; // @[Switch.scala 33:19:@300.4]
  wire [47:0] _GEN_42; // @[Switch.scala 33:19:@300.4]
  wire [47:0] _GEN_43; // @[Switch.scala 33:19:@300.4]
  wire [47:0] _GEN_44; // @[Switch.scala 33:19:@300.4]
  wire [47:0] _GEN_45; // @[Switch.scala 33:19:@300.4]
  wire [47:0] _GEN_46; // @[Switch.scala 33:19:@300.4]
  wire [47:0] _GEN_47; // @[Switch.scala 33:19:@300.4]
  wire [47:0] _GEN_48; // @[Switch.scala 33:19:@300.4]
  wire [47:0] _GEN_49; // @[Switch.scala 33:19:@300.4]
  wire [47:0] _GEN_50; // @[Switch.scala 33:19:@300.4]
  wire [47:0] _GEN_51; // @[Switch.scala 33:19:@300.4]
  wire [47:0] _GEN_52; // @[Switch.scala 33:19:@300.4]
  wire [47:0] _GEN_53; // @[Switch.scala 33:19:@300.4]
  wire [47:0] _GEN_54; // @[Switch.scala 33:19:@300.4]
  wire [47:0] _GEN_55; // @[Switch.scala 33:19:@300.4]
  wire [47:0] _GEN_56; // @[Switch.scala 33:19:@300.4]
  wire [47:0] _GEN_57; // @[Switch.scala 33:19:@300.4]
  wire [47:0] _GEN_58; // @[Switch.scala 33:19:@300.4]
  wire [47:0] _GEN_59; // @[Switch.scala 33:19:@300.4]
  wire [47:0] _GEN_60; // @[Switch.scala 33:19:@300.4]
  wire [47:0] _GEN_61; // @[Switch.scala 33:19:@300.4]
  wire [47:0] _GEN_62; // @[Switch.scala 33:19:@300.4]
  wire [7:0] _T_5116; // @[Switch.scala 34:32:@307.4]
  wire [15:0] _T_5124; // @[Switch.scala 34:32:@315.4]
  wire [7:0] _T_5131; // @[Switch.scala 34:32:@322.4]
  wire [31:0] _T_5140; // @[Switch.scala 34:32:@331.4]
  wire  _T_5144; // @[Switch.scala 30:53:@334.4]
  wire  valid_2_0; // @[Switch.scala 30:36:@335.4]
  wire  _T_5147; // @[Switch.scala 30:53:@337.4]
  wire  valid_2_1; // @[Switch.scala 30:36:@338.4]
  wire  _T_5150; // @[Switch.scala 30:53:@340.4]
  wire  valid_2_2; // @[Switch.scala 30:36:@341.4]
  wire  _T_5153; // @[Switch.scala 30:53:@343.4]
  wire  valid_2_3; // @[Switch.scala 30:36:@344.4]
  wire  _T_5156; // @[Switch.scala 30:53:@346.4]
  wire  valid_2_4; // @[Switch.scala 30:36:@347.4]
  wire  _T_5159; // @[Switch.scala 30:53:@349.4]
  wire  valid_2_5; // @[Switch.scala 30:36:@350.4]
  wire  _T_5162; // @[Switch.scala 30:53:@352.4]
  wire  valid_2_6; // @[Switch.scala 30:36:@353.4]
  wire  _T_5165; // @[Switch.scala 30:53:@355.4]
  wire  valid_2_7; // @[Switch.scala 30:36:@356.4]
  wire  _T_5168; // @[Switch.scala 30:53:@358.4]
  wire  valid_2_8; // @[Switch.scala 30:36:@359.4]
  wire  _T_5171; // @[Switch.scala 30:53:@361.4]
  wire  valid_2_9; // @[Switch.scala 30:36:@362.4]
  wire  _T_5174; // @[Switch.scala 30:53:@364.4]
  wire  valid_2_10; // @[Switch.scala 30:36:@365.4]
  wire  _T_5177; // @[Switch.scala 30:53:@367.4]
  wire  valid_2_11; // @[Switch.scala 30:36:@368.4]
  wire  _T_5180; // @[Switch.scala 30:53:@370.4]
  wire  valid_2_12; // @[Switch.scala 30:36:@371.4]
  wire  _T_5183; // @[Switch.scala 30:53:@373.4]
  wire  valid_2_13; // @[Switch.scala 30:36:@374.4]
  wire  _T_5186; // @[Switch.scala 30:53:@376.4]
  wire  valid_2_14; // @[Switch.scala 30:36:@377.4]
  wire  _T_5189; // @[Switch.scala 30:53:@379.4]
  wire  valid_2_15; // @[Switch.scala 30:36:@380.4]
  wire  _T_5192; // @[Switch.scala 30:53:@382.4]
  wire  valid_2_16; // @[Switch.scala 30:36:@383.4]
  wire  _T_5195; // @[Switch.scala 30:53:@385.4]
  wire  valid_2_17; // @[Switch.scala 30:36:@386.4]
  wire  _T_5198; // @[Switch.scala 30:53:@388.4]
  wire  valid_2_18; // @[Switch.scala 30:36:@389.4]
  wire  _T_5201; // @[Switch.scala 30:53:@391.4]
  wire  valid_2_19; // @[Switch.scala 30:36:@392.4]
  wire  _T_5204; // @[Switch.scala 30:53:@394.4]
  wire  valid_2_20; // @[Switch.scala 30:36:@395.4]
  wire  _T_5207; // @[Switch.scala 30:53:@397.4]
  wire  valid_2_21; // @[Switch.scala 30:36:@398.4]
  wire  _T_5210; // @[Switch.scala 30:53:@400.4]
  wire  valid_2_22; // @[Switch.scala 30:36:@401.4]
  wire  _T_5213; // @[Switch.scala 30:53:@403.4]
  wire  valid_2_23; // @[Switch.scala 30:36:@404.4]
  wire  _T_5216; // @[Switch.scala 30:53:@406.4]
  wire  valid_2_24; // @[Switch.scala 30:36:@407.4]
  wire  _T_5219; // @[Switch.scala 30:53:@409.4]
  wire  valid_2_25; // @[Switch.scala 30:36:@410.4]
  wire  _T_5222; // @[Switch.scala 30:53:@412.4]
  wire  valid_2_26; // @[Switch.scala 30:36:@413.4]
  wire  _T_5225; // @[Switch.scala 30:53:@415.4]
  wire  valid_2_27; // @[Switch.scala 30:36:@416.4]
  wire  _T_5228; // @[Switch.scala 30:53:@418.4]
  wire  valid_2_28; // @[Switch.scala 30:36:@419.4]
  wire  _T_5231; // @[Switch.scala 30:53:@421.4]
  wire  valid_2_29; // @[Switch.scala 30:36:@422.4]
  wire  _T_5234; // @[Switch.scala 30:53:@424.4]
  wire  valid_2_30; // @[Switch.scala 30:36:@425.4]
  wire  _T_5237; // @[Switch.scala 30:53:@427.4]
  wire  valid_2_31; // @[Switch.scala 30:36:@428.4]
  wire [4:0] _T_5271; // @[Mux.scala 31:69:@430.4]
  wire [4:0] _T_5272; // @[Mux.scala 31:69:@431.4]
  wire [4:0] _T_5273; // @[Mux.scala 31:69:@432.4]
  wire [4:0] _T_5274; // @[Mux.scala 31:69:@433.4]
  wire [4:0] _T_5275; // @[Mux.scala 31:69:@434.4]
  wire [4:0] _T_5276; // @[Mux.scala 31:69:@435.4]
  wire [4:0] _T_5277; // @[Mux.scala 31:69:@436.4]
  wire [4:0] _T_5278; // @[Mux.scala 31:69:@437.4]
  wire [4:0] _T_5279; // @[Mux.scala 31:69:@438.4]
  wire [4:0] _T_5280; // @[Mux.scala 31:69:@439.4]
  wire [4:0] _T_5281; // @[Mux.scala 31:69:@440.4]
  wire [4:0] _T_5282; // @[Mux.scala 31:69:@441.4]
  wire [4:0] _T_5283; // @[Mux.scala 31:69:@442.4]
  wire [4:0] _T_5284; // @[Mux.scala 31:69:@443.4]
  wire [4:0] _T_5285; // @[Mux.scala 31:69:@444.4]
  wire [4:0] _T_5286; // @[Mux.scala 31:69:@445.4]
  wire [4:0] _T_5287; // @[Mux.scala 31:69:@446.4]
  wire [4:0] _T_5288; // @[Mux.scala 31:69:@447.4]
  wire [4:0] _T_5289; // @[Mux.scala 31:69:@448.4]
  wire [4:0] _T_5290; // @[Mux.scala 31:69:@449.4]
  wire [4:0] _T_5291; // @[Mux.scala 31:69:@450.4]
  wire [4:0] _T_5292; // @[Mux.scala 31:69:@451.4]
  wire [4:0] _T_5293; // @[Mux.scala 31:69:@452.4]
  wire [4:0] _T_5294; // @[Mux.scala 31:69:@453.4]
  wire [4:0] _T_5295; // @[Mux.scala 31:69:@454.4]
  wire [4:0] _T_5296; // @[Mux.scala 31:69:@455.4]
  wire [4:0] _T_5297; // @[Mux.scala 31:69:@456.4]
  wire [4:0] _T_5298; // @[Mux.scala 31:69:@457.4]
  wire [4:0] _T_5299; // @[Mux.scala 31:69:@458.4]
  wire [4:0] _T_5300; // @[Mux.scala 31:69:@459.4]
  wire [4:0] select_2; // @[Mux.scala 31:69:@460.4]
  wire [47:0] _GEN_65; // @[Switch.scala 33:19:@462.4]
  wire [47:0] _GEN_66; // @[Switch.scala 33:19:@462.4]
  wire [47:0] _GEN_67; // @[Switch.scala 33:19:@462.4]
  wire [47:0] _GEN_68; // @[Switch.scala 33:19:@462.4]
  wire [47:0] _GEN_69; // @[Switch.scala 33:19:@462.4]
  wire [47:0] _GEN_70; // @[Switch.scala 33:19:@462.4]
  wire [47:0] _GEN_71; // @[Switch.scala 33:19:@462.4]
  wire [47:0] _GEN_72; // @[Switch.scala 33:19:@462.4]
  wire [47:0] _GEN_73; // @[Switch.scala 33:19:@462.4]
  wire [47:0] _GEN_74; // @[Switch.scala 33:19:@462.4]
  wire [47:0] _GEN_75; // @[Switch.scala 33:19:@462.4]
  wire [47:0] _GEN_76; // @[Switch.scala 33:19:@462.4]
  wire [47:0] _GEN_77; // @[Switch.scala 33:19:@462.4]
  wire [47:0] _GEN_78; // @[Switch.scala 33:19:@462.4]
  wire [47:0] _GEN_79; // @[Switch.scala 33:19:@462.4]
  wire [47:0] _GEN_80; // @[Switch.scala 33:19:@462.4]
  wire [47:0] _GEN_81; // @[Switch.scala 33:19:@462.4]
  wire [47:0] _GEN_82; // @[Switch.scala 33:19:@462.4]
  wire [47:0] _GEN_83; // @[Switch.scala 33:19:@462.4]
  wire [47:0] _GEN_84; // @[Switch.scala 33:19:@462.4]
  wire [47:0] _GEN_85; // @[Switch.scala 33:19:@462.4]
  wire [47:0] _GEN_86; // @[Switch.scala 33:19:@462.4]
  wire [47:0] _GEN_87; // @[Switch.scala 33:19:@462.4]
  wire [47:0] _GEN_88; // @[Switch.scala 33:19:@462.4]
  wire [47:0] _GEN_89; // @[Switch.scala 33:19:@462.4]
  wire [47:0] _GEN_90; // @[Switch.scala 33:19:@462.4]
  wire [47:0] _GEN_91; // @[Switch.scala 33:19:@462.4]
  wire [47:0] _GEN_92; // @[Switch.scala 33:19:@462.4]
  wire [47:0] _GEN_93; // @[Switch.scala 33:19:@462.4]
  wire [47:0] _GEN_94; // @[Switch.scala 33:19:@462.4]
  wire [7:0] _T_5309; // @[Switch.scala 34:32:@469.4]
  wire [15:0] _T_5317; // @[Switch.scala 34:32:@477.4]
  wire [7:0] _T_5324; // @[Switch.scala 34:32:@484.4]
  wire [31:0] _T_5333; // @[Switch.scala 34:32:@493.4]
  wire  _T_5337; // @[Switch.scala 30:53:@496.4]
  wire  valid_3_0; // @[Switch.scala 30:36:@497.4]
  wire  _T_5340; // @[Switch.scala 30:53:@499.4]
  wire  valid_3_1; // @[Switch.scala 30:36:@500.4]
  wire  _T_5343; // @[Switch.scala 30:53:@502.4]
  wire  valid_3_2; // @[Switch.scala 30:36:@503.4]
  wire  _T_5346; // @[Switch.scala 30:53:@505.4]
  wire  valid_3_3; // @[Switch.scala 30:36:@506.4]
  wire  _T_5349; // @[Switch.scala 30:53:@508.4]
  wire  valid_3_4; // @[Switch.scala 30:36:@509.4]
  wire  _T_5352; // @[Switch.scala 30:53:@511.4]
  wire  valid_3_5; // @[Switch.scala 30:36:@512.4]
  wire  _T_5355; // @[Switch.scala 30:53:@514.4]
  wire  valid_3_6; // @[Switch.scala 30:36:@515.4]
  wire  _T_5358; // @[Switch.scala 30:53:@517.4]
  wire  valid_3_7; // @[Switch.scala 30:36:@518.4]
  wire  _T_5361; // @[Switch.scala 30:53:@520.4]
  wire  valid_3_8; // @[Switch.scala 30:36:@521.4]
  wire  _T_5364; // @[Switch.scala 30:53:@523.4]
  wire  valid_3_9; // @[Switch.scala 30:36:@524.4]
  wire  _T_5367; // @[Switch.scala 30:53:@526.4]
  wire  valid_3_10; // @[Switch.scala 30:36:@527.4]
  wire  _T_5370; // @[Switch.scala 30:53:@529.4]
  wire  valid_3_11; // @[Switch.scala 30:36:@530.4]
  wire  _T_5373; // @[Switch.scala 30:53:@532.4]
  wire  valid_3_12; // @[Switch.scala 30:36:@533.4]
  wire  _T_5376; // @[Switch.scala 30:53:@535.4]
  wire  valid_3_13; // @[Switch.scala 30:36:@536.4]
  wire  _T_5379; // @[Switch.scala 30:53:@538.4]
  wire  valid_3_14; // @[Switch.scala 30:36:@539.4]
  wire  _T_5382; // @[Switch.scala 30:53:@541.4]
  wire  valid_3_15; // @[Switch.scala 30:36:@542.4]
  wire  _T_5385; // @[Switch.scala 30:53:@544.4]
  wire  valid_3_16; // @[Switch.scala 30:36:@545.4]
  wire  _T_5388; // @[Switch.scala 30:53:@547.4]
  wire  valid_3_17; // @[Switch.scala 30:36:@548.4]
  wire  _T_5391; // @[Switch.scala 30:53:@550.4]
  wire  valid_3_18; // @[Switch.scala 30:36:@551.4]
  wire  _T_5394; // @[Switch.scala 30:53:@553.4]
  wire  valid_3_19; // @[Switch.scala 30:36:@554.4]
  wire  _T_5397; // @[Switch.scala 30:53:@556.4]
  wire  valid_3_20; // @[Switch.scala 30:36:@557.4]
  wire  _T_5400; // @[Switch.scala 30:53:@559.4]
  wire  valid_3_21; // @[Switch.scala 30:36:@560.4]
  wire  _T_5403; // @[Switch.scala 30:53:@562.4]
  wire  valid_3_22; // @[Switch.scala 30:36:@563.4]
  wire  _T_5406; // @[Switch.scala 30:53:@565.4]
  wire  valid_3_23; // @[Switch.scala 30:36:@566.4]
  wire  _T_5409; // @[Switch.scala 30:53:@568.4]
  wire  valid_3_24; // @[Switch.scala 30:36:@569.4]
  wire  _T_5412; // @[Switch.scala 30:53:@571.4]
  wire  valid_3_25; // @[Switch.scala 30:36:@572.4]
  wire  _T_5415; // @[Switch.scala 30:53:@574.4]
  wire  valid_3_26; // @[Switch.scala 30:36:@575.4]
  wire  _T_5418; // @[Switch.scala 30:53:@577.4]
  wire  valid_3_27; // @[Switch.scala 30:36:@578.4]
  wire  _T_5421; // @[Switch.scala 30:53:@580.4]
  wire  valid_3_28; // @[Switch.scala 30:36:@581.4]
  wire  _T_5424; // @[Switch.scala 30:53:@583.4]
  wire  valid_3_29; // @[Switch.scala 30:36:@584.4]
  wire  _T_5427; // @[Switch.scala 30:53:@586.4]
  wire  valid_3_30; // @[Switch.scala 30:36:@587.4]
  wire  _T_5430; // @[Switch.scala 30:53:@589.4]
  wire  valid_3_31; // @[Switch.scala 30:36:@590.4]
  wire [4:0] _T_5464; // @[Mux.scala 31:69:@592.4]
  wire [4:0] _T_5465; // @[Mux.scala 31:69:@593.4]
  wire [4:0] _T_5466; // @[Mux.scala 31:69:@594.4]
  wire [4:0] _T_5467; // @[Mux.scala 31:69:@595.4]
  wire [4:0] _T_5468; // @[Mux.scala 31:69:@596.4]
  wire [4:0] _T_5469; // @[Mux.scala 31:69:@597.4]
  wire [4:0] _T_5470; // @[Mux.scala 31:69:@598.4]
  wire [4:0] _T_5471; // @[Mux.scala 31:69:@599.4]
  wire [4:0] _T_5472; // @[Mux.scala 31:69:@600.4]
  wire [4:0] _T_5473; // @[Mux.scala 31:69:@601.4]
  wire [4:0] _T_5474; // @[Mux.scala 31:69:@602.4]
  wire [4:0] _T_5475; // @[Mux.scala 31:69:@603.4]
  wire [4:0] _T_5476; // @[Mux.scala 31:69:@604.4]
  wire [4:0] _T_5477; // @[Mux.scala 31:69:@605.4]
  wire [4:0] _T_5478; // @[Mux.scala 31:69:@606.4]
  wire [4:0] _T_5479; // @[Mux.scala 31:69:@607.4]
  wire [4:0] _T_5480; // @[Mux.scala 31:69:@608.4]
  wire [4:0] _T_5481; // @[Mux.scala 31:69:@609.4]
  wire [4:0] _T_5482; // @[Mux.scala 31:69:@610.4]
  wire [4:0] _T_5483; // @[Mux.scala 31:69:@611.4]
  wire [4:0] _T_5484; // @[Mux.scala 31:69:@612.4]
  wire [4:0] _T_5485; // @[Mux.scala 31:69:@613.4]
  wire [4:0] _T_5486; // @[Mux.scala 31:69:@614.4]
  wire [4:0] _T_5487; // @[Mux.scala 31:69:@615.4]
  wire [4:0] _T_5488; // @[Mux.scala 31:69:@616.4]
  wire [4:0] _T_5489; // @[Mux.scala 31:69:@617.4]
  wire [4:0] _T_5490; // @[Mux.scala 31:69:@618.4]
  wire [4:0] _T_5491; // @[Mux.scala 31:69:@619.4]
  wire [4:0] _T_5492; // @[Mux.scala 31:69:@620.4]
  wire [4:0] _T_5493; // @[Mux.scala 31:69:@621.4]
  wire [4:0] select_3; // @[Mux.scala 31:69:@622.4]
  wire [47:0] _GEN_97; // @[Switch.scala 33:19:@624.4]
  wire [47:0] _GEN_98; // @[Switch.scala 33:19:@624.4]
  wire [47:0] _GEN_99; // @[Switch.scala 33:19:@624.4]
  wire [47:0] _GEN_100; // @[Switch.scala 33:19:@624.4]
  wire [47:0] _GEN_101; // @[Switch.scala 33:19:@624.4]
  wire [47:0] _GEN_102; // @[Switch.scala 33:19:@624.4]
  wire [47:0] _GEN_103; // @[Switch.scala 33:19:@624.4]
  wire [47:0] _GEN_104; // @[Switch.scala 33:19:@624.4]
  wire [47:0] _GEN_105; // @[Switch.scala 33:19:@624.4]
  wire [47:0] _GEN_106; // @[Switch.scala 33:19:@624.4]
  wire [47:0] _GEN_107; // @[Switch.scala 33:19:@624.4]
  wire [47:0] _GEN_108; // @[Switch.scala 33:19:@624.4]
  wire [47:0] _GEN_109; // @[Switch.scala 33:19:@624.4]
  wire [47:0] _GEN_110; // @[Switch.scala 33:19:@624.4]
  wire [47:0] _GEN_111; // @[Switch.scala 33:19:@624.4]
  wire [47:0] _GEN_112; // @[Switch.scala 33:19:@624.4]
  wire [47:0] _GEN_113; // @[Switch.scala 33:19:@624.4]
  wire [47:0] _GEN_114; // @[Switch.scala 33:19:@624.4]
  wire [47:0] _GEN_115; // @[Switch.scala 33:19:@624.4]
  wire [47:0] _GEN_116; // @[Switch.scala 33:19:@624.4]
  wire [47:0] _GEN_117; // @[Switch.scala 33:19:@624.4]
  wire [47:0] _GEN_118; // @[Switch.scala 33:19:@624.4]
  wire [47:0] _GEN_119; // @[Switch.scala 33:19:@624.4]
  wire [47:0] _GEN_120; // @[Switch.scala 33:19:@624.4]
  wire [47:0] _GEN_121; // @[Switch.scala 33:19:@624.4]
  wire [47:0] _GEN_122; // @[Switch.scala 33:19:@624.4]
  wire [47:0] _GEN_123; // @[Switch.scala 33:19:@624.4]
  wire [47:0] _GEN_124; // @[Switch.scala 33:19:@624.4]
  wire [47:0] _GEN_125; // @[Switch.scala 33:19:@624.4]
  wire [47:0] _GEN_126; // @[Switch.scala 33:19:@624.4]
  wire [7:0] _T_5502; // @[Switch.scala 34:32:@631.4]
  wire [15:0] _T_5510; // @[Switch.scala 34:32:@639.4]
  wire [7:0] _T_5517; // @[Switch.scala 34:32:@646.4]
  wire [31:0] _T_5526; // @[Switch.scala 34:32:@655.4]
  wire  _T_5530; // @[Switch.scala 30:53:@658.4]
  wire  valid_4_0; // @[Switch.scala 30:36:@659.4]
  wire  _T_5533; // @[Switch.scala 30:53:@661.4]
  wire  valid_4_1; // @[Switch.scala 30:36:@662.4]
  wire  _T_5536; // @[Switch.scala 30:53:@664.4]
  wire  valid_4_2; // @[Switch.scala 30:36:@665.4]
  wire  _T_5539; // @[Switch.scala 30:53:@667.4]
  wire  valid_4_3; // @[Switch.scala 30:36:@668.4]
  wire  _T_5542; // @[Switch.scala 30:53:@670.4]
  wire  valid_4_4; // @[Switch.scala 30:36:@671.4]
  wire  _T_5545; // @[Switch.scala 30:53:@673.4]
  wire  valid_4_5; // @[Switch.scala 30:36:@674.4]
  wire  _T_5548; // @[Switch.scala 30:53:@676.4]
  wire  valid_4_6; // @[Switch.scala 30:36:@677.4]
  wire  _T_5551; // @[Switch.scala 30:53:@679.4]
  wire  valid_4_7; // @[Switch.scala 30:36:@680.4]
  wire  _T_5554; // @[Switch.scala 30:53:@682.4]
  wire  valid_4_8; // @[Switch.scala 30:36:@683.4]
  wire  _T_5557; // @[Switch.scala 30:53:@685.4]
  wire  valid_4_9; // @[Switch.scala 30:36:@686.4]
  wire  _T_5560; // @[Switch.scala 30:53:@688.4]
  wire  valid_4_10; // @[Switch.scala 30:36:@689.4]
  wire  _T_5563; // @[Switch.scala 30:53:@691.4]
  wire  valid_4_11; // @[Switch.scala 30:36:@692.4]
  wire  _T_5566; // @[Switch.scala 30:53:@694.4]
  wire  valid_4_12; // @[Switch.scala 30:36:@695.4]
  wire  _T_5569; // @[Switch.scala 30:53:@697.4]
  wire  valid_4_13; // @[Switch.scala 30:36:@698.4]
  wire  _T_5572; // @[Switch.scala 30:53:@700.4]
  wire  valid_4_14; // @[Switch.scala 30:36:@701.4]
  wire  _T_5575; // @[Switch.scala 30:53:@703.4]
  wire  valid_4_15; // @[Switch.scala 30:36:@704.4]
  wire  _T_5578; // @[Switch.scala 30:53:@706.4]
  wire  valid_4_16; // @[Switch.scala 30:36:@707.4]
  wire  _T_5581; // @[Switch.scala 30:53:@709.4]
  wire  valid_4_17; // @[Switch.scala 30:36:@710.4]
  wire  _T_5584; // @[Switch.scala 30:53:@712.4]
  wire  valid_4_18; // @[Switch.scala 30:36:@713.4]
  wire  _T_5587; // @[Switch.scala 30:53:@715.4]
  wire  valid_4_19; // @[Switch.scala 30:36:@716.4]
  wire  _T_5590; // @[Switch.scala 30:53:@718.4]
  wire  valid_4_20; // @[Switch.scala 30:36:@719.4]
  wire  _T_5593; // @[Switch.scala 30:53:@721.4]
  wire  valid_4_21; // @[Switch.scala 30:36:@722.4]
  wire  _T_5596; // @[Switch.scala 30:53:@724.4]
  wire  valid_4_22; // @[Switch.scala 30:36:@725.4]
  wire  _T_5599; // @[Switch.scala 30:53:@727.4]
  wire  valid_4_23; // @[Switch.scala 30:36:@728.4]
  wire  _T_5602; // @[Switch.scala 30:53:@730.4]
  wire  valid_4_24; // @[Switch.scala 30:36:@731.4]
  wire  _T_5605; // @[Switch.scala 30:53:@733.4]
  wire  valid_4_25; // @[Switch.scala 30:36:@734.4]
  wire  _T_5608; // @[Switch.scala 30:53:@736.4]
  wire  valid_4_26; // @[Switch.scala 30:36:@737.4]
  wire  _T_5611; // @[Switch.scala 30:53:@739.4]
  wire  valid_4_27; // @[Switch.scala 30:36:@740.4]
  wire  _T_5614; // @[Switch.scala 30:53:@742.4]
  wire  valid_4_28; // @[Switch.scala 30:36:@743.4]
  wire  _T_5617; // @[Switch.scala 30:53:@745.4]
  wire  valid_4_29; // @[Switch.scala 30:36:@746.4]
  wire  _T_5620; // @[Switch.scala 30:53:@748.4]
  wire  valid_4_30; // @[Switch.scala 30:36:@749.4]
  wire  _T_5623; // @[Switch.scala 30:53:@751.4]
  wire  valid_4_31; // @[Switch.scala 30:36:@752.4]
  wire [4:0] _T_5657; // @[Mux.scala 31:69:@754.4]
  wire [4:0] _T_5658; // @[Mux.scala 31:69:@755.4]
  wire [4:0] _T_5659; // @[Mux.scala 31:69:@756.4]
  wire [4:0] _T_5660; // @[Mux.scala 31:69:@757.4]
  wire [4:0] _T_5661; // @[Mux.scala 31:69:@758.4]
  wire [4:0] _T_5662; // @[Mux.scala 31:69:@759.4]
  wire [4:0] _T_5663; // @[Mux.scala 31:69:@760.4]
  wire [4:0] _T_5664; // @[Mux.scala 31:69:@761.4]
  wire [4:0] _T_5665; // @[Mux.scala 31:69:@762.4]
  wire [4:0] _T_5666; // @[Mux.scala 31:69:@763.4]
  wire [4:0] _T_5667; // @[Mux.scala 31:69:@764.4]
  wire [4:0] _T_5668; // @[Mux.scala 31:69:@765.4]
  wire [4:0] _T_5669; // @[Mux.scala 31:69:@766.4]
  wire [4:0] _T_5670; // @[Mux.scala 31:69:@767.4]
  wire [4:0] _T_5671; // @[Mux.scala 31:69:@768.4]
  wire [4:0] _T_5672; // @[Mux.scala 31:69:@769.4]
  wire [4:0] _T_5673; // @[Mux.scala 31:69:@770.4]
  wire [4:0] _T_5674; // @[Mux.scala 31:69:@771.4]
  wire [4:0] _T_5675; // @[Mux.scala 31:69:@772.4]
  wire [4:0] _T_5676; // @[Mux.scala 31:69:@773.4]
  wire [4:0] _T_5677; // @[Mux.scala 31:69:@774.4]
  wire [4:0] _T_5678; // @[Mux.scala 31:69:@775.4]
  wire [4:0] _T_5679; // @[Mux.scala 31:69:@776.4]
  wire [4:0] _T_5680; // @[Mux.scala 31:69:@777.4]
  wire [4:0] _T_5681; // @[Mux.scala 31:69:@778.4]
  wire [4:0] _T_5682; // @[Mux.scala 31:69:@779.4]
  wire [4:0] _T_5683; // @[Mux.scala 31:69:@780.4]
  wire [4:0] _T_5684; // @[Mux.scala 31:69:@781.4]
  wire [4:0] _T_5685; // @[Mux.scala 31:69:@782.4]
  wire [4:0] _T_5686; // @[Mux.scala 31:69:@783.4]
  wire [4:0] select_4; // @[Mux.scala 31:69:@784.4]
  wire [47:0] _GEN_129; // @[Switch.scala 33:19:@786.4]
  wire [47:0] _GEN_130; // @[Switch.scala 33:19:@786.4]
  wire [47:0] _GEN_131; // @[Switch.scala 33:19:@786.4]
  wire [47:0] _GEN_132; // @[Switch.scala 33:19:@786.4]
  wire [47:0] _GEN_133; // @[Switch.scala 33:19:@786.4]
  wire [47:0] _GEN_134; // @[Switch.scala 33:19:@786.4]
  wire [47:0] _GEN_135; // @[Switch.scala 33:19:@786.4]
  wire [47:0] _GEN_136; // @[Switch.scala 33:19:@786.4]
  wire [47:0] _GEN_137; // @[Switch.scala 33:19:@786.4]
  wire [47:0] _GEN_138; // @[Switch.scala 33:19:@786.4]
  wire [47:0] _GEN_139; // @[Switch.scala 33:19:@786.4]
  wire [47:0] _GEN_140; // @[Switch.scala 33:19:@786.4]
  wire [47:0] _GEN_141; // @[Switch.scala 33:19:@786.4]
  wire [47:0] _GEN_142; // @[Switch.scala 33:19:@786.4]
  wire [47:0] _GEN_143; // @[Switch.scala 33:19:@786.4]
  wire [47:0] _GEN_144; // @[Switch.scala 33:19:@786.4]
  wire [47:0] _GEN_145; // @[Switch.scala 33:19:@786.4]
  wire [47:0] _GEN_146; // @[Switch.scala 33:19:@786.4]
  wire [47:0] _GEN_147; // @[Switch.scala 33:19:@786.4]
  wire [47:0] _GEN_148; // @[Switch.scala 33:19:@786.4]
  wire [47:0] _GEN_149; // @[Switch.scala 33:19:@786.4]
  wire [47:0] _GEN_150; // @[Switch.scala 33:19:@786.4]
  wire [47:0] _GEN_151; // @[Switch.scala 33:19:@786.4]
  wire [47:0] _GEN_152; // @[Switch.scala 33:19:@786.4]
  wire [47:0] _GEN_153; // @[Switch.scala 33:19:@786.4]
  wire [47:0] _GEN_154; // @[Switch.scala 33:19:@786.4]
  wire [47:0] _GEN_155; // @[Switch.scala 33:19:@786.4]
  wire [47:0] _GEN_156; // @[Switch.scala 33:19:@786.4]
  wire [47:0] _GEN_157; // @[Switch.scala 33:19:@786.4]
  wire [47:0] _GEN_158; // @[Switch.scala 33:19:@786.4]
  wire [7:0] _T_5695; // @[Switch.scala 34:32:@793.4]
  wire [15:0] _T_5703; // @[Switch.scala 34:32:@801.4]
  wire [7:0] _T_5710; // @[Switch.scala 34:32:@808.4]
  wire [31:0] _T_5719; // @[Switch.scala 34:32:@817.4]
  wire  _T_5723; // @[Switch.scala 30:53:@820.4]
  wire  valid_5_0; // @[Switch.scala 30:36:@821.4]
  wire  _T_5726; // @[Switch.scala 30:53:@823.4]
  wire  valid_5_1; // @[Switch.scala 30:36:@824.4]
  wire  _T_5729; // @[Switch.scala 30:53:@826.4]
  wire  valid_5_2; // @[Switch.scala 30:36:@827.4]
  wire  _T_5732; // @[Switch.scala 30:53:@829.4]
  wire  valid_5_3; // @[Switch.scala 30:36:@830.4]
  wire  _T_5735; // @[Switch.scala 30:53:@832.4]
  wire  valid_5_4; // @[Switch.scala 30:36:@833.4]
  wire  _T_5738; // @[Switch.scala 30:53:@835.4]
  wire  valid_5_5; // @[Switch.scala 30:36:@836.4]
  wire  _T_5741; // @[Switch.scala 30:53:@838.4]
  wire  valid_5_6; // @[Switch.scala 30:36:@839.4]
  wire  _T_5744; // @[Switch.scala 30:53:@841.4]
  wire  valid_5_7; // @[Switch.scala 30:36:@842.4]
  wire  _T_5747; // @[Switch.scala 30:53:@844.4]
  wire  valid_5_8; // @[Switch.scala 30:36:@845.4]
  wire  _T_5750; // @[Switch.scala 30:53:@847.4]
  wire  valid_5_9; // @[Switch.scala 30:36:@848.4]
  wire  _T_5753; // @[Switch.scala 30:53:@850.4]
  wire  valid_5_10; // @[Switch.scala 30:36:@851.4]
  wire  _T_5756; // @[Switch.scala 30:53:@853.4]
  wire  valid_5_11; // @[Switch.scala 30:36:@854.4]
  wire  _T_5759; // @[Switch.scala 30:53:@856.4]
  wire  valid_5_12; // @[Switch.scala 30:36:@857.4]
  wire  _T_5762; // @[Switch.scala 30:53:@859.4]
  wire  valid_5_13; // @[Switch.scala 30:36:@860.4]
  wire  _T_5765; // @[Switch.scala 30:53:@862.4]
  wire  valid_5_14; // @[Switch.scala 30:36:@863.4]
  wire  _T_5768; // @[Switch.scala 30:53:@865.4]
  wire  valid_5_15; // @[Switch.scala 30:36:@866.4]
  wire  _T_5771; // @[Switch.scala 30:53:@868.4]
  wire  valid_5_16; // @[Switch.scala 30:36:@869.4]
  wire  _T_5774; // @[Switch.scala 30:53:@871.4]
  wire  valid_5_17; // @[Switch.scala 30:36:@872.4]
  wire  _T_5777; // @[Switch.scala 30:53:@874.4]
  wire  valid_5_18; // @[Switch.scala 30:36:@875.4]
  wire  _T_5780; // @[Switch.scala 30:53:@877.4]
  wire  valid_5_19; // @[Switch.scala 30:36:@878.4]
  wire  _T_5783; // @[Switch.scala 30:53:@880.4]
  wire  valid_5_20; // @[Switch.scala 30:36:@881.4]
  wire  _T_5786; // @[Switch.scala 30:53:@883.4]
  wire  valid_5_21; // @[Switch.scala 30:36:@884.4]
  wire  _T_5789; // @[Switch.scala 30:53:@886.4]
  wire  valid_5_22; // @[Switch.scala 30:36:@887.4]
  wire  _T_5792; // @[Switch.scala 30:53:@889.4]
  wire  valid_5_23; // @[Switch.scala 30:36:@890.4]
  wire  _T_5795; // @[Switch.scala 30:53:@892.4]
  wire  valid_5_24; // @[Switch.scala 30:36:@893.4]
  wire  _T_5798; // @[Switch.scala 30:53:@895.4]
  wire  valid_5_25; // @[Switch.scala 30:36:@896.4]
  wire  _T_5801; // @[Switch.scala 30:53:@898.4]
  wire  valid_5_26; // @[Switch.scala 30:36:@899.4]
  wire  _T_5804; // @[Switch.scala 30:53:@901.4]
  wire  valid_5_27; // @[Switch.scala 30:36:@902.4]
  wire  _T_5807; // @[Switch.scala 30:53:@904.4]
  wire  valid_5_28; // @[Switch.scala 30:36:@905.4]
  wire  _T_5810; // @[Switch.scala 30:53:@907.4]
  wire  valid_5_29; // @[Switch.scala 30:36:@908.4]
  wire  _T_5813; // @[Switch.scala 30:53:@910.4]
  wire  valid_5_30; // @[Switch.scala 30:36:@911.4]
  wire  _T_5816; // @[Switch.scala 30:53:@913.4]
  wire  valid_5_31; // @[Switch.scala 30:36:@914.4]
  wire [4:0] _T_5850; // @[Mux.scala 31:69:@916.4]
  wire [4:0] _T_5851; // @[Mux.scala 31:69:@917.4]
  wire [4:0] _T_5852; // @[Mux.scala 31:69:@918.4]
  wire [4:0] _T_5853; // @[Mux.scala 31:69:@919.4]
  wire [4:0] _T_5854; // @[Mux.scala 31:69:@920.4]
  wire [4:0] _T_5855; // @[Mux.scala 31:69:@921.4]
  wire [4:0] _T_5856; // @[Mux.scala 31:69:@922.4]
  wire [4:0] _T_5857; // @[Mux.scala 31:69:@923.4]
  wire [4:0] _T_5858; // @[Mux.scala 31:69:@924.4]
  wire [4:0] _T_5859; // @[Mux.scala 31:69:@925.4]
  wire [4:0] _T_5860; // @[Mux.scala 31:69:@926.4]
  wire [4:0] _T_5861; // @[Mux.scala 31:69:@927.4]
  wire [4:0] _T_5862; // @[Mux.scala 31:69:@928.4]
  wire [4:0] _T_5863; // @[Mux.scala 31:69:@929.4]
  wire [4:0] _T_5864; // @[Mux.scala 31:69:@930.4]
  wire [4:0] _T_5865; // @[Mux.scala 31:69:@931.4]
  wire [4:0] _T_5866; // @[Mux.scala 31:69:@932.4]
  wire [4:0] _T_5867; // @[Mux.scala 31:69:@933.4]
  wire [4:0] _T_5868; // @[Mux.scala 31:69:@934.4]
  wire [4:0] _T_5869; // @[Mux.scala 31:69:@935.4]
  wire [4:0] _T_5870; // @[Mux.scala 31:69:@936.4]
  wire [4:0] _T_5871; // @[Mux.scala 31:69:@937.4]
  wire [4:0] _T_5872; // @[Mux.scala 31:69:@938.4]
  wire [4:0] _T_5873; // @[Mux.scala 31:69:@939.4]
  wire [4:0] _T_5874; // @[Mux.scala 31:69:@940.4]
  wire [4:0] _T_5875; // @[Mux.scala 31:69:@941.4]
  wire [4:0] _T_5876; // @[Mux.scala 31:69:@942.4]
  wire [4:0] _T_5877; // @[Mux.scala 31:69:@943.4]
  wire [4:0] _T_5878; // @[Mux.scala 31:69:@944.4]
  wire [4:0] _T_5879; // @[Mux.scala 31:69:@945.4]
  wire [4:0] select_5; // @[Mux.scala 31:69:@946.4]
  wire [47:0] _GEN_161; // @[Switch.scala 33:19:@948.4]
  wire [47:0] _GEN_162; // @[Switch.scala 33:19:@948.4]
  wire [47:0] _GEN_163; // @[Switch.scala 33:19:@948.4]
  wire [47:0] _GEN_164; // @[Switch.scala 33:19:@948.4]
  wire [47:0] _GEN_165; // @[Switch.scala 33:19:@948.4]
  wire [47:0] _GEN_166; // @[Switch.scala 33:19:@948.4]
  wire [47:0] _GEN_167; // @[Switch.scala 33:19:@948.4]
  wire [47:0] _GEN_168; // @[Switch.scala 33:19:@948.4]
  wire [47:0] _GEN_169; // @[Switch.scala 33:19:@948.4]
  wire [47:0] _GEN_170; // @[Switch.scala 33:19:@948.4]
  wire [47:0] _GEN_171; // @[Switch.scala 33:19:@948.4]
  wire [47:0] _GEN_172; // @[Switch.scala 33:19:@948.4]
  wire [47:0] _GEN_173; // @[Switch.scala 33:19:@948.4]
  wire [47:0] _GEN_174; // @[Switch.scala 33:19:@948.4]
  wire [47:0] _GEN_175; // @[Switch.scala 33:19:@948.4]
  wire [47:0] _GEN_176; // @[Switch.scala 33:19:@948.4]
  wire [47:0] _GEN_177; // @[Switch.scala 33:19:@948.4]
  wire [47:0] _GEN_178; // @[Switch.scala 33:19:@948.4]
  wire [47:0] _GEN_179; // @[Switch.scala 33:19:@948.4]
  wire [47:0] _GEN_180; // @[Switch.scala 33:19:@948.4]
  wire [47:0] _GEN_181; // @[Switch.scala 33:19:@948.4]
  wire [47:0] _GEN_182; // @[Switch.scala 33:19:@948.4]
  wire [47:0] _GEN_183; // @[Switch.scala 33:19:@948.4]
  wire [47:0] _GEN_184; // @[Switch.scala 33:19:@948.4]
  wire [47:0] _GEN_185; // @[Switch.scala 33:19:@948.4]
  wire [47:0] _GEN_186; // @[Switch.scala 33:19:@948.4]
  wire [47:0] _GEN_187; // @[Switch.scala 33:19:@948.4]
  wire [47:0] _GEN_188; // @[Switch.scala 33:19:@948.4]
  wire [47:0] _GEN_189; // @[Switch.scala 33:19:@948.4]
  wire [47:0] _GEN_190; // @[Switch.scala 33:19:@948.4]
  wire [7:0] _T_5888; // @[Switch.scala 34:32:@955.4]
  wire [15:0] _T_5896; // @[Switch.scala 34:32:@963.4]
  wire [7:0] _T_5903; // @[Switch.scala 34:32:@970.4]
  wire [31:0] _T_5912; // @[Switch.scala 34:32:@979.4]
  wire  _T_5916; // @[Switch.scala 30:53:@982.4]
  wire  valid_6_0; // @[Switch.scala 30:36:@983.4]
  wire  _T_5919; // @[Switch.scala 30:53:@985.4]
  wire  valid_6_1; // @[Switch.scala 30:36:@986.4]
  wire  _T_5922; // @[Switch.scala 30:53:@988.4]
  wire  valid_6_2; // @[Switch.scala 30:36:@989.4]
  wire  _T_5925; // @[Switch.scala 30:53:@991.4]
  wire  valid_6_3; // @[Switch.scala 30:36:@992.4]
  wire  _T_5928; // @[Switch.scala 30:53:@994.4]
  wire  valid_6_4; // @[Switch.scala 30:36:@995.4]
  wire  _T_5931; // @[Switch.scala 30:53:@997.4]
  wire  valid_6_5; // @[Switch.scala 30:36:@998.4]
  wire  _T_5934; // @[Switch.scala 30:53:@1000.4]
  wire  valid_6_6; // @[Switch.scala 30:36:@1001.4]
  wire  _T_5937; // @[Switch.scala 30:53:@1003.4]
  wire  valid_6_7; // @[Switch.scala 30:36:@1004.4]
  wire  _T_5940; // @[Switch.scala 30:53:@1006.4]
  wire  valid_6_8; // @[Switch.scala 30:36:@1007.4]
  wire  _T_5943; // @[Switch.scala 30:53:@1009.4]
  wire  valid_6_9; // @[Switch.scala 30:36:@1010.4]
  wire  _T_5946; // @[Switch.scala 30:53:@1012.4]
  wire  valid_6_10; // @[Switch.scala 30:36:@1013.4]
  wire  _T_5949; // @[Switch.scala 30:53:@1015.4]
  wire  valid_6_11; // @[Switch.scala 30:36:@1016.4]
  wire  _T_5952; // @[Switch.scala 30:53:@1018.4]
  wire  valid_6_12; // @[Switch.scala 30:36:@1019.4]
  wire  _T_5955; // @[Switch.scala 30:53:@1021.4]
  wire  valid_6_13; // @[Switch.scala 30:36:@1022.4]
  wire  _T_5958; // @[Switch.scala 30:53:@1024.4]
  wire  valid_6_14; // @[Switch.scala 30:36:@1025.4]
  wire  _T_5961; // @[Switch.scala 30:53:@1027.4]
  wire  valid_6_15; // @[Switch.scala 30:36:@1028.4]
  wire  _T_5964; // @[Switch.scala 30:53:@1030.4]
  wire  valid_6_16; // @[Switch.scala 30:36:@1031.4]
  wire  _T_5967; // @[Switch.scala 30:53:@1033.4]
  wire  valid_6_17; // @[Switch.scala 30:36:@1034.4]
  wire  _T_5970; // @[Switch.scala 30:53:@1036.4]
  wire  valid_6_18; // @[Switch.scala 30:36:@1037.4]
  wire  _T_5973; // @[Switch.scala 30:53:@1039.4]
  wire  valid_6_19; // @[Switch.scala 30:36:@1040.4]
  wire  _T_5976; // @[Switch.scala 30:53:@1042.4]
  wire  valid_6_20; // @[Switch.scala 30:36:@1043.4]
  wire  _T_5979; // @[Switch.scala 30:53:@1045.4]
  wire  valid_6_21; // @[Switch.scala 30:36:@1046.4]
  wire  _T_5982; // @[Switch.scala 30:53:@1048.4]
  wire  valid_6_22; // @[Switch.scala 30:36:@1049.4]
  wire  _T_5985; // @[Switch.scala 30:53:@1051.4]
  wire  valid_6_23; // @[Switch.scala 30:36:@1052.4]
  wire  _T_5988; // @[Switch.scala 30:53:@1054.4]
  wire  valid_6_24; // @[Switch.scala 30:36:@1055.4]
  wire  _T_5991; // @[Switch.scala 30:53:@1057.4]
  wire  valid_6_25; // @[Switch.scala 30:36:@1058.4]
  wire  _T_5994; // @[Switch.scala 30:53:@1060.4]
  wire  valid_6_26; // @[Switch.scala 30:36:@1061.4]
  wire  _T_5997; // @[Switch.scala 30:53:@1063.4]
  wire  valid_6_27; // @[Switch.scala 30:36:@1064.4]
  wire  _T_6000; // @[Switch.scala 30:53:@1066.4]
  wire  valid_6_28; // @[Switch.scala 30:36:@1067.4]
  wire  _T_6003; // @[Switch.scala 30:53:@1069.4]
  wire  valid_6_29; // @[Switch.scala 30:36:@1070.4]
  wire  _T_6006; // @[Switch.scala 30:53:@1072.4]
  wire  valid_6_30; // @[Switch.scala 30:36:@1073.4]
  wire  _T_6009; // @[Switch.scala 30:53:@1075.4]
  wire  valid_6_31; // @[Switch.scala 30:36:@1076.4]
  wire [4:0] _T_6043; // @[Mux.scala 31:69:@1078.4]
  wire [4:0] _T_6044; // @[Mux.scala 31:69:@1079.4]
  wire [4:0] _T_6045; // @[Mux.scala 31:69:@1080.4]
  wire [4:0] _T_6046; // @[Mux.scala 31:69:@1081.4]
  wire [4:0] _T_6047; // @[Mux.scala 31:69:@1082.4]
  wire [4:0] _T_6048; // @[Mux.scala 31:69:@1083.4]
  wire [4:0] _T_6049; // @[Mux.scala 31:69:@1084.4]
  wire [4:0] _T_6050; // @[Mux.scala 31:69:@1085.4]
  wire [4:0] _T_6051; // @[Mux.scala 31:69:@1086.4]
  wire [4:0] _T_6052; // @[Mux.scala 31:69:@1087.4]
  wire [4:0] _T_6053; // @[Mux.scala 31:69:@1088.4]
  wire [4:0] _T_6054; // @[Mux.scala 31:69:@1089.4]
  wire [4:0] _T_6055; // @[Mux.scala 31:69:@1090.4]
  wire [4:0] _T_6056; // @[Mux.scala 31:69:@1091.4]
  wire [4:0] _T_6057; // @[Mux.scala 31:69:@1092.4]
  wire [4:0] _T_6058; // @[Mux.scala 31:69:@1093.4]
  wire [4:0] _T_6059; // @[Mux.scala 31:69:@1094.4]
  wire [4:0] _T_6060; // @[Mux.scala 31:69:@1095.4]
  wire [4:0] _T_6061; // @[Mux.scala 31:69:@1096.4]
  wire [4:0] _T_6062; // @[Mux.scala 31:69:@1097.4]
  wire [4:0] _T_6063; // @[Mux.scala 31:69:@1098.4]
  wire [4:0] _T_6064; // @[Mux.scala 31:69:@1099.4]
  wire [4:0] _T_6065; // @[Mux.scala 31:69:@1100.4]
  wire [4:0] _T_6066; // @[Mux.scala 31:69:@1101.4]
  wire [4:0] _T_6067; // @[Mux.scala 31:69:@1102.4]
  wire [4:0] _T_6068; // @[Mux.scala 31:69:@1103.4]
  wire [4:0] _T_6069; // @[Mux.scala 31:69:@1104.4]
  wire [4:0] _T_6070; // @[Mux.scala 31:69:@1105.4]
  wire [4:0] _T_6071; // @[Mux.scala 31:69:@1106.4]
  wire [4:0] _T_6072; // @[Mux.scala 31:69:@1107.4]
  wire [4:0] select_6; // @[Mux.scala 31:69:@1108.4]
  wire [47:0] _GEN_193; // @[Switch.scala 33:19:@1110.4]
  wire [47:0] _GEN_194; // @[Switch.scala 33:19:@1110.4]
  wire [47:0] _GEN_195; // @[Switch.scala 33:19:@1110.4]
  wire [47:0] _GEN_196; // @[Switch.scala 33:19:@1110.4]
  wire [47:0] _GEN_197; // @[Switch.scala 33:19:@1110.4]
  wire [47:0] _GEN_198; // @[Switch.scala 33:19:@1110.4]
  wire [47:0] _GEN_199; // @[Switch.scala 33:19:@1110.4]
  wire [47:0] _GEN_200; // @[Switch.scala 33:19:@1110.4]
  wire [47:0] _GEN_201; // @[Switch.scala 33:19:@1110.4]
  wire [47:0] _GEN_202; // @[Switch.scala 33:19:@1110.4]
  wire [47:0] _GEN_203; // @[Switch.scala 33:19:@1110.4]
  wire [47:0] _GEN_204; // @[Switch.scala 33:19:@1110.4]
  wire [47:0] _GEN_205; // @[Switch.scala 33:19:@1110.4]
  wire [47:0] _GEN_206; // @[Switch.scala 33:19:@1110.4]
  wire [47:0] _GEN_207; // @[Switch.scala 33:19:@1110.4]
  wire [47:0] _GEN_208; // @[Switch.scala 33:19:@1110.4]
  wire [47:0] _GEN_209; // @[Switch.scala 33:19:@1110.4]
  wire [47:0] _GEN_210; // @[Switch.scala 33:19:@1110.4]
  wire [47:0] _GEN_211; // @[Switch.scala 33:19:@1110.4]
  wire [47:0] _GEN_212; // @[Switch.scala 33:19:@1110.4]
  wire [47:0] _GEN_213; // @[Switch.scala 33:19:@1110.4]
  wire [47:0] _GEN_214; // @[Switch.scala 33:19:@1110.4]
  wire [47:0] _GEN_215; // @[Switch.scala 33:19:@1110.4]
  wire [47:0] _GEN_216; // @[Switch.scala 33:19:@1110.4]
  wire [47:0] _GEN_217; // @[Switch.scala 33:19:@1110.4]
  wire [47:0] _GEN_218; // @[Switch.scala 33:19:@1110.4]
  wire [47:0] _GEN_219; // @[Switch.scala 33:19:@1110.4]
  wire [47:0] _GEN_220; // @[Switch.scala 33:19:@1110.4]
  wire [47:0] _GEN_221; // @[Switch.scala 33:19:@1110.4]
  wire [47:0] _GEN_222; // @[Switch.scala 33:19:@1110.4]
  wire [7:0] _T_6081; // @[Switch.scala 34:32:@1117.4]
  wire [15:0] _T_6089; // @[Switch.scala 34:32:@1125.4]
  wire [7:0] _T_6096; // @[Switch.scala 34:32:@1132.4]
  wire [31:0] _T_6105; // @[Switch.scala 34:32:@1141.4]
  wire  _T_6109; // @[Switch.scala 30:53:@1144.4]
  wire  valid_7_0; // @[Switch.scala 30:36:@1145.4]
  wire  _T_6112; // @[Switch.scala 30:53:@1147.4]
  wire  valid_7_1; // @[Switch.scala 30:36:@1148.4]
  wire  _T_6115; // @[Switch.scala 30:53:@1150.4]
  wire  valid_7_2; // @[Switch.scala 30:36:@1151.4]
  wire  _T_6118; // @[Switch.scala 30:53:@1153.4]
  wire  valid_7_3; // @[Switch.scala 30:36:@1154.4]
  wire  _T_6121; // @[Switch.scala 30:53:@1156.4]
  wire  valid_7_4; // @[Switch.scala 30:36:@1157.4]
  wire  _T_6124; // @[Switch.scala 30:53:@1159.4]
  wire  valid_7_5; // @[Switch.scala 30:36:@1160.4]
  wire  _T_6127; // @[Switch.scala 30:53:@1162.4]
  wire  valid_7_6; // @[Switch.scala 30:36:@1163.4]
  wire  _T_6130; // @[Switch.scala 30:53:@1165.4]
  wire  valid_7_7; // @[Switch.scala 30:36:@1166.4]
  wire  _T_6133; // @[Switch.scala 30:53:@1168.4]
  wire  valid_7_8; // @[Switch.scala 30:36:@1169.4]
  wire  _T_6136; // @[Switch.scala 30:53:@1171.4]
  wire  valid_7_9; // @[Switch.scala 30:36:@1172.4]
  wire  _T_6139; // @[Switch.scala 30:53:@1174.4]
  wire  valid_7_10; // @[Switch.scala 30:36:@1175.4]
  wire  _T_6142; // @[Switch.scala 30:53:@1177.4]
  wire  valid_7_11; // @[Switch.scala 30:36:@1178.4]
  wire  _T_6145; // @[Switch.scala 30:53:@1180.4]
  wire  valid_7_12; // @[Switch.scala 30:36:@1181.4]
  wire  _T_6148; // @[Switch.scala 30:53:@1183.4]
  wire  valid_7_13; // @[Switch.scala 30:36:@1184.4]
  wire  _T_6151; // @[Switch.scala 30:53:@1186.4]
  wire  valid_7_14; // @[Switch.scala 30:36:@1187.4]
  wire  _T_6154; // @[Switch.scala 30:53:@1189.4]
  wire  valid_7_15; // @[Switch.scala 30:36:@1190.4]
  wire  _T_6157; // @[Switch.scala 30:53:@1192.4]
  wire  valid_7_16; // @[Switch.scala 30:36:@1193.4]
  wire  _T_6160; // @[Switch.scala 30:53:@1195.4]
  wire  valid_7_17; // @[Switch.scala 30:36:@1196.4]
  wire  _T_6163; // @[Switch.scala 30:53:@1198.4]
  wire  valid_7_18; // @[Switch.scala 30:36:@1199.4]
  wire  _T_6166; // @[Switch.scala 30:53:@1201.4]
  wire  valid_7_19; // @[Switch.scala 30:36:@1202.4]
  wire  _T_6169; // @[Switch.scala 30:53:@1204.4]
  wire  valid_7_20; // @[Switch.scala 30:36:@1205.4]
  wire  _T_6172; // @[Switch.scala 30:53:@1207.4]
  wire  valid_7_21; // @[Switch.scala 30:36:@1208.4]
  wire  _T_6175; // @[Switch.scala 30:53:@1210.4]
  wire  valid_7_22; // @[Switch.scala 30:36:@1211.4]
  wire  _T_6178; // @[Switch.scala 30:53:@1213.4]
  wire  valid_7_23; // @[Switch.scala 30:36:@1214.4]
  wire  _T_6181; // @[Switch.scala 30:53:@1216.4]
  wire  valid_7_24; // @[Switch.scala 30:36:@1217.4]
  wire  _T_6184; // @[Switch.scala 30:53:@1219.4]
  wire  valid_7_25; // @[Switch.scala 30:36:@1220.4]
  wire  _T_6187; // @[Switch.scala 30:53:@1222.4]
  wire  valid_7_26; // @[Switch.scala 30:36:@1223.4]
  wire  _T_6190; // @[Switch.scala 30:53:@1225.4]
  wire  valid_7_27; // @[Switch.scala 30:36:@1226.4]
  wire  _T_6193; // @[Switch.scala 30:53:@1228.4]
  wire  valid_7_28; // @[Switch.scala 30:36:@1229.4]
  wire  _T_6196; // @[Switch.scala 30:53:@1231.4]
  wire  valid_7_29; // @[Switch.scala 30:36:@1232.4]
  wire  _T_6199; // @[Switch.scala 30:53:@1234.4]
  wire  valid_7_30; // @[Switch.scala 30:36:@1235.4]
  wire  _T_6202; // @[Switch.scala 30:53:@1237.4]
  wire  valid_7_31; // @[Switch.scala 30:36:@1238.4]
  wire [4:0] _T_6236; // @[Mux.scala 31:69:@1240.4]
  wire [4:0] _T_6237; // @[Mux.scala 31:69:@1241.4]
  wire [4:0] _T_6238; // @[Mux.scala 31:69:@1242.4]
  wire [4:0] _T_6239; // @[Mux.scala 31:69:@1243.4]
  wire [4:0] _T_6240; // @[Mux.scala 31:69:@1244.4]
  wire [4:0] _T_6241; // @[Mux.scala 31:69:@1245.4]
  wire [4:0] _T_6242; // @[Mux.scala 31:69:@1246.4]
  wire [4:0] _T_6243; // @[Mux.scala 31:69:@1247.4]
  wire [4:0] _T_6244; // @[Mux.scala 31:69:@1248.4]
  wire [4:0] _T_6245; // @[Mux.scala 31:69:@1249.4]
  wire [4:0] _T_6246; // @[Mux.scala 31:69:@1250.4]
  wire [4:0] _T_6247; // @[Mux.scala 31:69:@1251.4]
  wire [4:0] _T_6248; // @[Mux.scala 31:69:@1252.4]
  wire [4:0] _T_6249; // @[Mux.scala 31:69:@1253.4]
  wire [4:0] _T_6250; // @[Mux.scala 31:69:@1254.4]
  wire [4:0] _T_6251; // @[Mux.scala 31:69:@1255.4]
  wire [4:0] _T_6252; // @[Mux.scala 31:69:@1256.4]
  wire [4:0] _T_6253; // @[Mux.scala 31:69:@1257.4]
  wire [4:0] _T_6254; // @[Mux.scala 31:69:@1258.4]
  wire [4:0] _T_6255; // @[Mux.scala 31:69:@1259.4]
  wire [4:0] _T_6256; // @[Mux.scala 31:69:@1260.4]
  wire [4:0] _T_6257; // @[Mux.scala 31:69:@1261.4]
  wire [4:0] _T_6258; // @[Mux.scala 31:69:@1262.4]
  wire [4:0] _T_6259; // @[Mux.scala 31:69:@1263.4]
  wire [4:0] _T_6260; // @[Mux.scala 31:69:@1264.4]
  wire [4:0] _T_6261; // @[Mux.scala 31:69:@1265.4]
  wire [4:0] _T_6262; // @[Mux.scala 31:69:@1266.4]
  wire [4:0] _T_6263; // @[Mux.scala 31:69:@1267.4]
  wire [4:0] _T_6264; // @[Mux.scala 31:69:@1268.4]
  wire [4:0] _T_6265; // @[Mux.scala 31:69:@1269.4]
  wire [4:0] select_7; // @[Mux.scala 31:69:@1270.4]
  wire [47:0] _GEN_225; // @[Switch.scala 33:19:@1272.4]
  wire [47:0] _GEN_226; // @[Switch.scala 33:19:@1272.4]
  wire [47:0] _GEN_227; // @[Switch.scala 33:19:@1272.4]
  wire [47:0] _GEN_228; // @[Switch.scala 33:19:@1272.4]
  wire [47:0] _GEN_229; // @[Switch.scala 33:19:@1272.4]
  wire [47:0] _GEN_230; // @[Switch.scala 33:19:@1272.4]
  wire [47:0] _GEN_231; // @[Switch.scala 33:19:@1272.4]
  wire [47:0] _GEN_232; // @[Switch.scala 33:19:@1272.4]
  wire [47:0] _GEN_233; // @[Switch.scala 33:19:@1272.4]
  wire [47:0] _GEN_234; // @[Switch.scala 33:19:@1272.4]
  wire [47:0] _GEN_235; // @[Switch.scala 33:19:@1272.4]
  wire [47:0] _GEN_236; // @[Switch.scala 33:19:@1272.4]
  wire [47:0] _GEN_237; // @[Switch.scala 33:19:@1272.4]
  wire [47:0] _GEN_238; // @[Switch.scala 33:19:@1272.4]
  wire [47:0] _GEN_239; // @[Switch.scala 33:19:@1272.4]
  wire [47:0] _GEN_240; // @[Switch.scala 33:19:@1272.4]
  wire [47:0] _GEN_241; // @[Switch.scala 33:19:@1272.4]
  wire [47:0] _GEN_242; // @[Switch.scala 33:19:@1272.4]
  wire [47:0] _GEN_243; // @[Switch.scala 33:19:@1272.4]
  wire [47:0] _GEN_244; // @[Switch.scala 33:19:@1272.4]
  wire [47:0] _GEN_245; // @[Switch.scala 33:19:@1272.4]
  wire [47:0] _GEN_246; // @[Switch.scala 33:19:@1272.4]
  wire [47:0] _GEN_247; // @[Switch.scala 33:19:@1272.4]
  wire [47:0] _GEN_248; // @[Switch.scala 33:19:@1272.4]
  wire [47:0] _GEN_249; // @[Switch.scala 33:19:@1272.4]
  wire [47:0] _GEN_250; // @[Switch.scala 33:19:@1272.4]
  wire [47:0] _GEN_251; // @[Switch.scala 33:19:@1272.4]
  wire [47:0] _GEN_252; // @[Switch.scala 33:19:@1272.4]
  wire [47:0] _GEN_253; // @[Switch.scala 33:19:@1272.4]
  wire [47:0] _GEN_254; // @[Switch.scala 33:19:@1272.4]
  wire [7:0] _T_6274; // @[Switch.scala 34:32:@1279.4]
  wire [15:0] _T_6282; // @[Switch.scala 34:32:@1287.4]
  wire [7:0] _T_6289; // @[Switch.scala 34:32:@1294.4]
  wire [31:0] _T_6298; // @[Switch.scala 34:32:@1303.4]
  wire  _T_6302; // @[Switch.scala 30:53:@1306.4]
  wire  valid_8_0; // @[Switch.scala 30:36:@1307.4]
  wire  _T_6305; // @[Switch.scala 30:53:@1309.4]
  wire  valid_8_1; // @[Switch.scala 30:36:@1310.4]
  wire  _T_6308; // @[Switch.scala 30:53:@1312.4]
  wire  valid_8_2; // @[Switch.scala 30:36:@1313.4]
  wire  _T_6311; // @[Switch.scala 30:53:@1315.4]
  wire  valid_8_3; // @[Switch.scala 30:36:@1316.4]
  wire  _T_6314; // @[Switch.scala 30:53:@1318.4]
  wire  valid_8_4; // @[Switch.scala 30:36:@1319.4]
  wire  _T_6317; // @[Switch.scala 30:53:@1321.4]
  wire  valid_8_5; // @[Switch.scala 30:36:@1322.4]
  wire  _T_6320; // @[Switch.scala 30:53:@1324.4]
  wire  valid_8_6; // @[Switch.scala 30:36:@1325.4]
  wire  _T_6323; // @[Switch.scala 30:53:@1327.4]
  wire  valid_8_7; // @[Switch.scala 30:36:@1328.4]
  wire  _T_6326; // @[Switch.scala 30:53:@1330.4]
  wire  valid_8_8; // @[Switch.scala 30:36:@1331.4]
  wire  _T_6329; // @[Switch.scala 30:53:@1333.4]
  wire  valid_8_9; // @[Switch.scala 30:36:@1334.4]
  wire  _T_6332; // @[Switch.scala 30:53:@1336.4]
  wire  valid_8_10; // @[Switch.scala 30:36:@1337.4]
  wire  _T_6335; // @[Switch.scala 30:53:@1339.4]
  wire  valid_8_11; // @[Switch.scala 30:36:@1340.4]
  wire  _T_6338; // @[Switch.scala 30:53:@1342.4]
  wire  valid_8_12; // @[Switch.scala 30:36:@1343.4]
  wire  _T_6341; // @[Switch.scala 30:53:@1345.4]
  wire  valid_8_13; // @[Switch.scala 30:36:@1346.4]
  wire  _T_6344; // @[Switch.scala 30:53:@1348.4]
  wire  valid_8_14; // @[Switch.scala 30:36:@1349.4]
  wire  _T_6347; // @[Switch.scala 30:53:@1351.4]
  wire  valid_8_15; // @[Switch.scala 30:36:@1352.4]
  wire  _T_6350; // @[Switch.scala 30:53:@1354.4]
  wire  valid_8_16; // @[Switch.scala 30:36:@1355.4]
  wire  _T_6353; // @[Switch.scala 30:53:@1357.4]
  wire  valid_8_17; // @[Switch.scala 30:36:@1358.4]
  wire  _T_6356; // @[Switch.scala 30:53:@1360.4]
  wire  valid_8_18; // @[Switch.scala 30:36:@1361.4]
  wire  _T_6359; // @[Switch.scala 30:53:@1363.4]
  wire  valid_8_19; // @[Switch.scala 30:36:@1364.4]
  wire  _T_6362; // @[Switch.scala 30:53:@1366.4]
  wire  valid_8_20; // @[Switch.scala 30:36:@1367.4]
  wire  _T_6365; // @[Switch.scala 30:53:@1369.4]
  wire  valid_8_21; // @[Switch.scala 30:36:@1370.4]
  wire  _T_6368; // @[Switch.scala 30:53:@1372.4]
  wire  valid_8_22; // @[Switch.scala 30:36:@1373.4]
  wire  _T_6371; // @[Switch.scala 30:53:@1375.4]
  wire  valid_8_23; // @[Switch.scala 30:36:@1376.4]
  wire  _T_6374; // @[Switch.scala 30:53:@1378.4]
  wire  valid_8_24; // @[Switch.scala 30:36:@1379.4]
  wire  _T_6377; // @[Switch.scala 30:53:@1381.4]
  wire  valid_8_25; // @[Switch.scala 30:36:@1382.4]
  wire  _T_6380; // @[Switch.scala 30:53:@1384.4]
  wire  valid_8_26; // @[Switch.scala 30:36:@1385.4]
  wire  _T_6383; // @[Switch.scala 30:53:@1387.4]
  wire  valid_8_27; // @[Switch.scala 30:36:@1388.4]
  wire  _T_6386; // @[Switch.scala 30:53:@1390.4]
  wire  valid_8_28; // @[Switch.scala 30:36:@1391.4]
  wire  _T_6389; // @[Switch.scala 30:53:@1393.4]
  wire  valid_8_29; // @[Switch.scala 30:36:@1394.4]
  wire  _T_6392; // @[Switch.scala 30:53:@1396.4]
  wire  valid_8_30; // @[Switch.scala 30:36:@1397.4]
  wire  _T_6395; // @[Switch.scala 30:53:@1399.4]
  wire  valid_8_31; // @[Switch.scala 30:36:@1400.4]
  wire [4:0] _T_6429; // @[Mux.scala 31:69:@1402.4]
  wire [4:0] _T_6430; // @[Mux.scala 31:69:@1403.4]
  wire [4:0] _T_6431; // @[Mux.scala 31:69:@1404.4]
  wire [4:0] _T_6432; // @[Mux.scala 31:69:@1405.4]
  wire [4:0] _T_6433; // @[Mux.scala 31:69:@1406.4]
  wire [4:0] _T_6434; // @[Mux.scala 31:69:@1407.4]
  wire [4:0] _T_6435; // @[Mux.scala 31:69:@1408.4]
  wire [4:0] _T_6436; // @[Mux.scala 31:69:@1409.4]
  wire [4:0] _T_6437; // @[Mux.scala 31:69:@1410.4]
  wire [4:0] _T_6438; // @[Mux.scala 31:69:@1411.4]
  wire [4:0] _T_6439; // @[Mux.scala 31:69:@1412.4]
  wire [4:0] _T_6440; // @[Mux.scala 31:69:@1413.4]
  wire [4:0] _T_6441; // @[Mux.scala 31:69:@1414.4]
  wire [4:0] _T_6442; // @[Mux.scala 31:69:@1415.4]
  wire [4:0] _T_6443; // @[Mux.scala 31:69:@1416.4]
  wire [4:0] _T_6444; // @[Mux.scala 31:69:@1417.4]
  wire [4:0] _T_6445; // @[Mux.scala 31:69:@1418.4]
  wire [4:0] _T_6446; // @[Mux.scala 31:69:@1419.4]
  wire [4:0] _T_6447; // @[Mux.scala 31:69:@1420.4]
  wire [4:0] _T_6448; // @[Mux.scala 31:69:@1421.4]
  wire [4:0] _T_6449; // @[Mux.scala 31:69:@1422.4]
  wire [4:0] _T_6450; // @[Mux.scala 31:69:@1423.4]
  wire [4:0] _T_6451; // @[Mux.scala 31:69:@1424.4]
  wire [4:0] _T_6452; // @[Mux.scala 31:69:@1425.4]
  wire [4:0] _T_6453; // @[Mux.scala 31:69:@1426.4]
  wire [4:0] _T_6454; // @[Mux.scala 31:69:@1427.4]
  wire [4:0] _T_6455; // @[Mux.scala 31:69:@1428.4]
  wire [4:0] _T_6456; // @[Mux.scala 31:69:@1429.4]
  wire [4:0] _T_6457; // @[Mux.scala 31:69:@1430.4]
  wire [4:0] _T_6458; // @[Mux.scala 31:69:@1431.4]
  wire [4:0] select_8; // @[Mux.scala 31:69:@1432.4]
  wire [47:0] _GEN_257; // @[Switch.scala 33:19:@1434.4]
  wire [47:0] _GEN_258; // @[Switch.scala 33:19:@1434.4]
  wire [47:0] _GEN_259; // @[Switch.scala 33:19:@1434.4]
  wire [47:0] _GEN_260; // @[Switch.scala 33:19:@1434.4]
  wire [47:0] _GEN_261; // @[Switch.scala 33:19:@1434.4]
  wire [47:0] _GEN_262; // @[Switch.scala 33:19:@1434.4]
  wire [47:0] _GEN_263; // @[Switch.scala 33:19:@1434.4]
  wire [47:0] _GEN_264; // @[Switch.scala 33:19:@1434.4]
  wire [47:0] _GEN_265; // @[Switch.scala 33:19:@1434.4]
  wire [47:0] _GEN_266; // @[Switch.scala 33:19:@1434.4]
  wire [47:0] _GEN_267; // @[Switch.scala 33:19:@1434.4]
  wire [47:0] _GEN_268; // @[Switch.scala 33:19:@1434.4]
  wire [47:0] _GEN_269; // @[Switch.scala 33:19:@1434.4]
  wire [47:0] _GEN_270; // @[Switch.scala 33:19:@1434.4]
  wire [47:0] _GEN_271; // @[Switch.scala 33:19:@1434.4]
  wire [47:0] _GEN_272; // @[Switch.scala 33:19:@1434.4]
  wire [47:0] _GEN_273; // @[Switch.scala 33:19:@1434.4]
  wire [47:0] _GEN_274; // @[Switch.scala 33:19:@1434.4]
  wire [47:0] _GEN_275; // @[Switch.scala 33:19:@1434.4]
  wire [47:0] _GEN_276; // @[Switch.scala 33:19:@1434.4]
  wire [47:0] _GEN_277; // @[Switch.scala 33:19:@1434.4]
  wire [47:0] _GEN_278; // @[Switch.scala 33:19:@1434.4]
  wire [47:0] _GEN_279; // @[Switch.scala 33:19:@1434.4]
  wire [47:0] _GEN_280; // @[Switch.scala 33:19:@1434.4]
  wire [47:0] _GEN_281; // @[Switch.scala 33:19:@1434.4]
  wire [47:0] _GEN_282; // @[Switch.scala 33:19:@1434.4]
  wire [47:0] _GEN_283; // @[Switch.scala 33:19:@1434.4]
  wire [47:0] _GEN_284; // @[Switch.scala 33:19:@1434.4]
  wire [47:0] _GEN_285; // @[Switch.scala 33:19:@1434.4]
  wire [47:0] _GEN_286; // @[Switch.scala 33:19:@1434.4]
  wire [7:0] _T_6467; // @[Switch.scala 34:32:@1441.4]
  wire [15:0] _T_6475; // @[Switch.scala 34:32:@1449.4]
  wire [7:0] _T_6482; // @[Switch.scala 34:32:@1456.4]
  wire [31:0] _T_6491; // @[Switch.scala 34:32:@1465.4]
  wire  _T_6495; // @[Switch.scala 30:53:@1468.4]
  wire  valid_9_0; // @[Switch.scala 30:36:@1469.4]
  wire  _T_6498; // @[Switch.scala 30:53:@1471.4]
  wire  valid_9_1; // @[Switch.scala 30:36:@1472.4]
  wire  _T_6501; // @[Switch.scala 30:53:@1474.4]
  wire  valid_9_2; // @[Switch.scala 30:36:@1475.4]
  wire  _T_6504; // @[Switch.scala 30:53:@1477.4]
  wire  valid_9_3; // @[Switch.scala 30:36:@1478.4]
  wire  _T_6507; // @[Switch.scala 30:53:@1480.4]
  wire  valid_9_4; // @[Switch.scala 30:36:@1481.4]
  wire  _T_6510; // @[Switch.scala 30:53:@1483.4]
  wire  valid_9_5; // @[Switch.scala 30:36:@1484.4]
  wire  _T_6513; // @[Switch.scala 30:53:@1486.4]
  wire  valid_9_6; // @[Switch.scala 30:36:@1487.4]
  wire  _T_6516; // @[Switch.scala 30:53:@1489.4]
  wire  valid_9_7; // @[Switch.scala 30:36:@1490.4]
  wire  _T_6519; // @[Switch.scala 30:53:@1492.4]
  wire  valid_9_8; // @[Switch.scala 30:36:@1493.4]
  wire  _T_6522; // @[Switch.scala 30:53:@1495.4]
  wire  valid_9_9; // @[Switch.scala 30:36:@1496.4]
  wire  _T_6525; // @[Switch.scala 30:53:@1498.4]
  wire  valid_9_10; // @[Switch.scala 30:36:@1499.4]
  wire  _T_6528; // @[Switch.scala 30:53:@1501.4]
  wire  valid_9_11; // @[Switch.scala 30:36:@1502.4]
  wire  _T_6531; // @[Switch.scala 30:53:@1504.4]
  wire  valid_9_12; // @[Switch.scala 30:36:@1505.4]
  wire  _T_6534; // @[Switch.scala 30:53:@1507.4]
  wire  valid_9_13; // @[Switch.scala 30:36:@1508.4]
  wire  _T_6537; // @[Switch.scala 30:53:@1510.4]
  wire  valid_9_14; // @[Switch.scala 30:36:@1511.4]
  wire  _T_6540; // @[Switch.scala 30:53:@1513.4]
  wire  valid_9_15; // @[Switch.scala 30:36:@1514.4]
  wire  _T_6543; // @[Switch.scala 30:53:@1516.4]
  wire  valid_9_16; // @[Switch.scala 30:36:@1517.4]
  wire  _T_6546; // @[Switch.scala 30:53:@1519.4]
  wire  valid_9_17; // @[Switch.scala 30:36:@1520.4]
  wire  _T_6549; // @[Switch.scala 30:53:@1522.4]
  wire  valid_9_18; // @[Switch.scala 30:36:@1523.4]
  wire  _T_6552; // @[Switch.scala 30:53:@1525.4]
  wire  valid_9_19; // @[Switch.scala 30:36:@1526.4]
  wire  _T_6555; // @[Switch.scala 30:53:@1528.4]
  wire  valid_9_20; // @[Switch.scala 30:36:@1529.4]
  wire  _T_6558; // @[Switch.scala 30:53:@1531.4]
  wire  valid_9_21; // @[Switch.scala 30:36:@1532.4]
  wire  _T_6561; // @[Switch.scala 30:53:@1534.4]
  wire  valid_9_22; // @[Switch.scala 30:36:@1535.4]
  wire  _T_6564; // @[Switch.scala 30:53:@1537.4]
  wire  valid_9_23; // @[Switch.scala 30:36:@1538.4]
  wire  _T_6567; // @[Switch.scala 30:53:@1540.4]
  wire  valid_9_24; // @[Switch.scala 30:36:@1541.4]
  wire  _T_6570; // @[Switch.scala 30:53:@1543.4]
  wire  valid_9_25; // @[Switch.scala 30:36:@1544.4]
  wire  _T_6573; // @[Switch.scala 30:53:@1546.4]
  wire  valid_9_26; // @[Switch.scala 30:36:@1547.4]
  wire  _T_6576; // @[Switch.scala 30:53:@1549.4]
  wire  valid_9_27; // @[Switch.scala 30:36:@1550.4]
  wire  _T_6579; // @[Switch.scala 30:53:@1552.4]
  wire  valid_9_28; // @[Switch.scala 30:36:@1553.4]
  wire  _T_6582; // @[Switch.scala 30:53:@1555.4]
  wire  valid_9_29; // @[Switch.scala 30:36:@1556.4]
  wire  _T_6585; // @[Switch.scala 30:53:@1558.4]
  wire  valid_9_30; // @[Switch.scala 30:36:@1559.4]
  wire  _T_6588; // @[Switch.scala 30:53:@1561.4]
  wire  valid_9_31; // @[Switch.scala 30:36:@1562.4]
  wire [4:0] _T_6622; // @[Mux.scala 31:69:@1564.4]
  wire [4:0] _T_6623; // @[Mux.scala 31:69:@1565.4]
  wire [4:0] _T_6624; // @[Mux.scala 31:69:@1566.4]
  wire [4:0] _T_6625; // @[Mux.scala 31:69:@1567.4]
  wire [4:0] _T_6626; // @[Mux.scala 31:69:@1568.4]
  wire [4:0] _T_6627; // @[Mux.scala 31:69:@1569.4]
  wire [4:0] _T_6628; // @[Mux.scala 31:69:@1570.4]
  wire [4:0] _T_6629; // @[Mux.scala 31:69:@1571.4]
  wire [4:0] _T_6630; // @[Mux.scala 31:69:@1572.4]
  wire [4:0] _T_6631; // @[Mux.scala 31:69:@1573.4]
  wire [4:0] _T_6632; // @[Mux.scala 31:69:@1574.4]
  wire [4:0] _T_6633; // @[Mux.scala 31:69:@1575.4]
  wire [4:0] _T_6634; // @[Mux.scala 31:69:@1576.4]
  wire [4:0] _T_6635; // @[Mux.scala 31:69:@1577.4]
  wire [4:0] _T_6636; // @[Mux.scala 31:69:@1578.4]
  wire [4:0] _T_6637; // @[Mux.scala 31:69:@1579.4]
  wire [4:0] _T_6638; // @[Mux.scala 31:69:@1580.4]
  wire [4:0] _T_6639; // @[Mux.scala 31:69:@1581.4]
  wire [4:0] _T_6640; // @[Mux.scala 31:69:@1582.4]
  wire [4:0] _T_6641; // @[Mux.scala 31:69:@1583.4]
  wire [4:0] _T_6642; // @[Mux.scala 31:69:@1584.4]
  wire [4:0] _T_6643; // @[Mux.scala 31:69:@1585.4]
  wire [4:0] _T_6644; // @[Mux.scala 31:69:@1586.4]
  wire [4:0] _T_6645; // @[Mux.scala 31:69:@1587.4]
  wire [4:0] _T_6646; // @[Mux.scala 31:69:@1588.4]
  wire [4:0] _T_6647; // @[Mux.scala 31:69:@1589.4]
  wire [4:0] _T_6648; // @[Mux.scala 31:69:@1590.4]
  wire [4:0] _T_6649; // @[Mux.scala 31:69:@1591.4]
  wire [4:0] _T_6650; // @[Mux.scala 31:69:@1592.4]
  wire [4:0] _T_6651; // @[Mux.scala 31:69:@1593.4]
  wire [4:0] select_9; // @[Mux.scala 31:69:@1594.4]
  wire [47:0] _GEN_289; // @[Switch.scala 33:19:@1596.4]
  wire [47:0] _GEN_290; // @[Switch.scala 33:19:@1596.4]
  wire [47:0] _GEN_291; // @[Switch.scala 33:19:@1596.4]
  wire [47:0] _GEN_292; // @[Switch.scala 33:19:@1596.4]
  wire [47:0] _GEN_293; // @[Switch.scala 33:19:@1596.4]
  wire [47:0] _GEN_294; // @[Switch.scala 33:19:@1596.4]
  wire [47:0] _GEN_295; // @[Switch.scala 33:19:@1596.4]
  wire [47:0] _GEN_296; // @[Switch.scala 33:19:@1596.4]
  wire [47:0] _GEN_297; // @[Switch.scala 33:19:@1596.4]
  wire [47:0] _GEN_298; // @[Switch.scala 33:19:@1596.4]
  wire [47:0] _GEN_299; // @[Switch.scala 33:19:@1596.4]
  wire [47:0] _GEN_300; // @[Switch.scala 33:19:@1596.4]
  wire [47:0] _GEN_301; // @[Switch.scala 33:19:@1596.4]
  wire [47:0] _GEN_302; // @[Switch.scala 33:19:@1596.4]
  wire [47:0] _GEN_303; // @[Switch.scala 33:19:@1596.4]
  wire [47:0] _GEN_304; // @[Switch.scala 33:19:@1596.4]
  wire [47:0] _GEN_305; // @[Switch.scala 33:19:@1596.4]
  wire [47:0] _GEN_306; // @[Switch.scala 33:19:@1596.4]
  wire [47:0] _GEN_307; // @[Switch.scala 33:19:@1596.4]
  wire [47:0] _GEN_308; // @[Switch.scala 33:19:@1596.4]
  wire [47:0] _GEN_309; // @[Switch.scala 33:19:@1596.4]
  wire [47:0] _GEN_310; // @[Switch.scala 33:19:@1596.4]
  wire [47:0] _GEN_311; // @[Switch.scala 33:19:@1596.4]
  wire [47:0] _GEN_312; // @[Switch.scala 33:19:@1596.4]
  wire [47:0] _GEN_313; // @[Switch.scala 33:19:@1596.4]
  wire [47:0] _GEN_314; // @[Switch.scala 33:19:@1596.4]
  wire [47:0] _GEN_315; // @[Switch.scala 33:19:@1596.4]
  wire [47:0] _GEN_316; // @[Switch.scala 33:19:@1596.4]
  wire [47:0] _GEN_317; // @[Switch.scala 33:19:@1596.4]
  wire [47:0] _GEN_318; // @[Switch.scala 33:19:@1596.4]
  wire [7:0] _T_6660; // @[Switch.scala 34:32:@1603.4]
  wire [15:0] _T_6668; // @[Switch.scala 34:32:@1611.4]
  wire [7:0] _T_6675; // @[Switch.scala 34:32:@1618.4]
  wire [31:0] _T_6684; // @[Switch.scala 34:32:@1627.4]
  wire  _T_6688; // @[Switch.scala 30:53:@1630.4]
  wire  valid_10_0; // @[Switch.scala 30:36:@1631.4]
  wire  _T_6691; // @[Switch.scala 30:53:@1633.4]
  wire  valid_10_1; // @[Switch.scala 30:36:@1634.4]
  wire  _T_6694; // @[Switch.scala 30:53:@1636.4]
  wire  valid_10_2; // @[Switch.scala 30:36:@1637.4]
  wire  _T_6697; // @[Switch.scala 30:53:@1639.4]
  wire  valid_10_3; // @[Switch.scala 30:36:@1640.4]
  wire  _T_6700; // @[Switch.scala 30:53:@1642.4]
  wire  valid_10_4; // @[Switch.scala 30:36:@1643.4]
  wire  _T_6703; // @[Switch.scala 30:53:@1645.4]
  wire  valid_10_5; // @[Switch.scala 30:36:@1646.4]
  wire  _T_6706; // @[Switch.scala 30:53:@1648.4]
  wire  valid_10_6; // @[Switch.scala 30:36:@1649.4]
  wire  _T_6709; // @[Switch.scala 30:53:@1651.4]
  wire  valid_10_7; // @[Switch.scala 30:36:@1652.4]
  wire  _T_6712; // @[Switch.scala 30:53:@1654.4]
  wire  valid_10_8; // @[Switch.scala 30:36:@1655.4]
  wire  _T_6715; // @[Switch.scala 30:53:@1657.4]
  wire  valid_10_9; // @[Switch.scala 30:36:@1658.4]
  wire  _T_6718; // @[Switch.scala 30:53:@1660.4]
  wire  valid_10_10; // @[Switch.scala 30:36:@1661.4]
  wire  _T_6721; // @[Switch.scala 30:53:@1663.4]
  wire  valid_10_11; // @[Switch.scala 30:36:@1664.4]
  wire  _T_6724; // @[Switch.scala 30:53:@1666.4]
  wire  valid_10_12; // @[Switch.scala 30:36:@1667.4]
  wire  _T_6727; // @[Switch.scala 30:53:@1669.4]
  wire  valid_10_13; // @[Switch.scala 30:36:@1670.4]
  wire  _T_6730; // @[Switch.scala 30:53:@1672.4]
  wire  valid_10_14; // @[Switch.scala 30:36:@1673.4]
  wire  _T_6733; // @[Switch.scala 30:53:@1675.4]
  wire  valid_10_15; // @[Switch.scala 30:36:@1676.4]
  wire  _T_6736; // @[Switch.scala 30:53:@1678.4]
  wire  valid_10_16; // @[Switch.scala 30:36:@1679.4]
  wire  _T_6739; // @[Switch.scala 30:53:@1681.4]
  wire  valid_10_17; // @[Switch.scala 30:36:@1682.4]
  wire  _T_6742; // @[Switch.scala 30:53:@1684.4]
  wire  valid_10_18; // @[Switch.scala 30:36:@1685.4]
  wire  _T_6745; // @[Switch.scala 30:53:@1687.4]
  wire  valid_10_19; // @[Switch.scala 30:36:@1688.4]
  wire  _T_6748; // @[Switch.scala 30:53:@1690.4]
  wire  valid_10_20; // @[Switch.scala 30:36:@1691.4]
  wire  _T_6751; // @[Switch.scala 30:53:@1693.4]
  wire  valid_10_21; // @[Switch.scala 30:36:@1694.4]
  wire  _T_6754; // @[Switch.scala 30:53:@1696.4]
  wire  valid_10_22; // @[Switch.scala 30:36:@1697.4]
  wire  _T_6757; // @[Switch.scala 30:53:@1699.4]
  wire  valid_10_23; // @[Switch.scala 30:36:@1700.4]
  wire  _T_6760; // @[Switch.scala 30:53:@1702.4]
  wire  valid_10_24; // @[Switch.scala 30:36:@1703.4]
  wire  _T_6763; // @[Switch.scala 30:53:@1705.4]
  wire  valid_10_25; // @[Switch.scala 30:36:@1706.4]
  wire  _T_6766; // @[Switch.scala 30:53:@1708.4]
  wire  valid_10_26; // @[Switch.scala 30:36:@1709.4]
  wire  _T_6769; // @[Switch.scala 30:53:@1711.4]
  wire  valid_10_27; // @[Switch.scala 30:36:@1712.4]
  wire  _T_6772; // @[Switch.scala 30:53:@1714.4]
  wire  valid_10_28; // @[Switch.scala 30:36:@1715.4]
  wire  _T_6775; // @[Switch.scala 30:53:@1717.4]
  wire  valid_10_29; // @[Switch.scala 30:36:@1718.4]
  wire  _T_6778; // @[Switch.scala 30:53:@1720.4]
  wire  valid_10_30; // @[Switch.scala 30:36:@1721.4]
  wire  _T_6781; // @[Switch.scala 30:53:@1723.4]
  wire  valid_10_31; // @[Switch.scala 30:36:@1724.4]
  wire [4:0] _T_6815; // @[Mux.scala 31:69:@1726.4]
  wire [4:0] _T_6816; // @[Mux.scala 31:69:@1727.4]
  wire [4:0] _T_6817; // @[Mux.scala 31:69:@1728.4]
  wire [4:0] _T_6818; // @[Mux.scala 31:69:@1729.4]
  wire [4:0] _T_6819; // @[Mux.scala 31:69:@1730.4]
  wire [4:0] _T_6820; // @[Mux.scala 31:69:@1731.4]
  wire [4:0] _T_6821; // @[Mux.scala 31:69:@1732.4]
  wire [4:0] _T_6822; // @[Mux.scala 31:69:@1733.4]
  wire [4:0] _T_6823; // @[Mux.scala 31:69:@1734.4]
  wire [4:0] _T_6824; // @[Mux.scala 31:69:@1735.4]
  wire [4:0] _T_6825; // @[Mux.scala 31:69:@1736.4]
  wire [4:0] _T_6826; // @[Mux.scala 31:69:@1737.4]
  wire [4:0] _T_6827; // @[Mux.scala 31:69:@1738.4]
  wire [4:0] _T_6828; // @[Mux.scala 31:69:@1739.4]
  wire [4:0] _T_6829; // @[Mux.scala 31:69:@1740.4]
  wire [4:0] _T_6830; // @[Mux.scala 31:69:@1741.4]
  wire [4:0] _T_6831; // @[Mux.scala 31:69:@1742.4]
  wire [4:0] _T_6832; // @[Mux.scala 31:69:@1743.4]
  wire [4:0] _T_6833; // @[Mux.scala 31:69:@1744.4]
  wire [4:0] _T_6834; // @[Mux.scala 31:69:@1745.4]
  wire [4:0] _T_6835; // @[Mux.scala 31:69:@1746.4]
  wire [4:0] _T_6836; // @[Mux.scala 31:69:@1747.4]
  wire [4:0] _T_6837; // @[Mux.scala 31:69:@1748.4]
  wire [4:0] _T_6838; // @[Mux.scala 31:69:@1749.4]
  wire [4:0] _T_6839; // @[Mux.scala 31:69:@1750.4]
  wire [4:0] _T_6840; // @[Mux.scala 31:69:@1751.4]
  wire [4:0] _T_6841; // @[Mux.scala 31:69:@1752.4]
  wire [4:0] _T_6842; // @[Mux.scala 31:69:@1753.4]
  wire [4:0] _T_6843; // @[Mux.scala 31:69:@1754.4]
  wire [4:0] _T_6844; // @[Mux.scala 31:69:@1755.4]
  wire [4:0] select_10; // @[Mux.scala 31:69:@1756.4]
  wire [47:0] _GEN_321; // @[Switch.scala 33:19:@1758.4]
  wire [47:0] _GEN_322; // @[Switch.scala 33:19:@1758.4]
  wire [47:0] _GEN_323; // @[Switch.scala 33:19:@1758.4]
  wire [47:0] _GEN_324; // @[Switch.scala 33:19:@1758.4]
  wire [47:0] _GEN_325; // @[Switch.scala 33:19:@1758.4]
  wire [47:0] _GEN_326; // @[Switch.scala 33:19:@1758.4]
  wire [47:0] _GEN_327; // @[Switch.scala 33:19:@1758.4]
  wire [47:0] _GEN_328; // @[Switch.scala 33:19:@1758.4]
  wire [47:0] _GEN_329; // @[Switch.scala 33:19:@1758.4]
  wire [47:0] _GEN_330; // @[Switch.scala 33:19:@1758.4]
  wire [47:0] _GEN_331; // @[Switch.scala 33:19:@1758.4]
  wire [47:0] _GEN_332; // @[Switch.scala 33:19:@1758.4]
  wire [47:0] _GEN_333; // @[Switch.scala 33:19:@1758.4]
  wire [47:0] _GEN_334; // @[Switch.scala 33:19:@1758.4]
  wire [47:0] _GEN_335; // @[Switch.scala 33:19:@1758.4]
  wire [47:0] _GEN_336; // @[Switch.scala 33:19:@1758.4]
  wire [47:0] _GEN_337; // @[Switch.scala 33:19:@1758.4]
  wire [47:0] _GEN_338; // @[Switch.scala 33:19:@1758.4]
  wire [47:0] _GEN_339; // @[Switch.scala 33:19:@1758.4]
  wire [47:0] _GEN_340; // @[Switch.scala 33:19:@1758.4]
  wire [47:0] _GEN_341; // @[Switch.scala 33:19:@1758.4]
  wire [47:0] _GEN_342; // @[Switch.scala 33:19:@1758.4]
  wire [47:0] _GEN_343; // @[Switch.scala 33:19:@1758.4]
  wire [47:0] _GEN_344; // @[Switch.scala 33:19:@1758.4]
  wire [47:0] _GEN_345; // @[Switch.scala 33:19:@1758.4]
  wire [47:0] _GEN_346; // @[Switch.scala 33:19:@1758.4]
  wire [47:0] _GEN_347; // @[Switch.scala 33:19:@1758.4]
  wire [47:0] _GEN_348; // @[Switch.scala 33:19:@1758.4]
  wire [47:0] _GEN_349; // @[Switch.scala 33:19:@1758.4]
  wire [47:0] _GEN_350; // @[Switch.scala 33:19:@1758.4]
  wire [7:0] _T_6853; // @[Switch.scala 34:32:@1765.4]
  wire [15:0] _T_6861; // @[Switch.scala 34:32:@1773.4]
  wire [7:0] _T_6868; // @[Switch.scala 34:32:@1780.4]
  wire [31:0] _T_6877; // @[Switch.scala 34:32:@1789.4]
  wire  _T_6881; // @[Switch.scala 30:53:@1792.4]
  wire  valid_11_0; // @[Switch.scala 30:36:@1793.4]
  wire  _T_6884; // @[Switch.scala 30:53:@1795.4]
  wire  valid_11_1; // @[Switch.scala 30:36:@1796.4]
  wire  _T_6887; // @[Switch.scala 30:53:@1798.4]
  wire  valid_11_2; // @[Switch.scala 30:36:@1799.4]
  wire  _T_6890; // @[Switch.scala 30:53:@1801.4]
  wire  valid_11_3; // @[Switch.scala 30:36:@1802.4]
  wire  _T_6893; // @[Switch.scala 30:53:@1804.4]
  wire  valid_11_4; // @[Switch.scala 30:36:@1805.4]
  wire  _T_6896; // @[Switch.scala 30:53:@1807.4]
  wire  valid_11_5; // @[Switch.scala 30:36:@1808.4]
  wire  _T_6899; // @[Switch.scala 30:53:@1810.4]
  wire  valid_11_6; // @[Switch.scala 30:36:@1811.4]
  wire  _T_6902; // @[Switch.scala 30:53:@1813.4]
  wire  valid_11_7; // @[Switch.scala 30:36:@1814.4]
  wire  _T_6905; // @[Switch.scala 30:53:@1816.4]
  wire  valid_11_8; // @[Switch.scala 30:36:@1817.4]
  wire  _T_6908; // @[Switch.scala 30:53:@1819.4]
  wire  valid_11_9; // @[Switch.scala 30:36:@1820.4]
  wire  _T_6911; // @[Switch.scala 30:53:@1822.4]
  wire  valid_11_10; // @[Switch.scala 30:36:@1823.4]
  wire  _T_6914; // @[Switch.scala 30:53:@1825.4]
  wire  valid_11_11; // @[Switch.scala 30:36:@1826.4]
  wire  _T_6917; // @[Switch.scala 30:53:@1828.4]
  wire  valid_11_12; // @[Switch.scala 30:36:@1829.4]
  wire  _T_6920; // @[Switch.scala 30:53:@1831.4]
  wire  valid_11_13; // @[Switch.scala 30:36:@1832.4]
  wire  _T_6923; // @[Switch.scala 30:53:@1834.4]
  wire  valid_11_14; // @[Switch.scala 30:36:@1835.4]
  wire  _T_6926; // @[Switch.scala 30:53:@1837.4]
  wire  valid_11_15; // @[Switch.scala 30:36:@1838.4]
  wire  _T_6929; // @[Switch.scala 30:53:@1840.4]
  wire  valid_11_16; // @[Switch.scala 30:36:@1841.4]
  wire  _T_6932; // @[Switch.scala 30:53:@1843.4]
  wire  valid_11_17; // @[Switch.scala 30:36:@1844.4]
  wire  _T_6935; // @[Switch.scala 30:53:@1846.4]
  wire  valid_11_18; // @[Switch.scala 30:36:@1847.4]
  wire  _T_6938; // @[Switch.scala 30:53:@1849.4]
  wire  valid_11_19; // @[Switch.scala 30:36:@1850.4]
  wire  _T_6941; // @[Switch.scala 30:53:@1852.4]
  wire  valid_11_20; // @[Switch.scala 30:36:@1853.4]
  wire  _T_6944; // @[Switch.scala 30:53:@1855.4]
  wire  valid_11_21; // @[Switch.scala 30:36:@1856.4]
  wire  _T_6947; // @[Switch.scala 30:53:@1858.4]
  wire  valid_11_22; // @[Switch.scala 30:36:@1859.4]
  wire  _T_6950; // @[Switch.scala 30:53:@1861.4]
  wire  valid_11_23; // @[Switch.scala 30:36:@1862.4]
  wire  _T_6953; // @[Switch.scala 30:53:@1864.4]
  wire  valid_11_24; // @[Switch.scala 30:36:@1865.4]
  wire  _T_6956; // @[Switch.scala 30:53:@1867.4]
  wire  valid_11_25; // @[Switch.scala 30:36:@1868.4]
  wire  _T_6959; // @[Switch.scala 30:53:@1870.4]
  wire  valid_11_26; // @[Switch.scala 30:36:@1871.4]
  wire  _T_6962; // @[Switch.scala 30:53:@1873.4]
  wire  valid_11_27; // @[Switch.scala 30:36:@1874.4]
  wire  _T_6965; // @[Switch.scala 30:53:@1876.4]
  wire  valid_11_28; // @[Switch.scala 30:36:@1877.4]
  wire  _T_6968; // @[Switch.scala 30:53:@1879.4]
  wire  valid_11_29; // @[Switch.scala 30:36:@1880.4]
  wire  _T_6971; // @[Switch.scala 30:53:@1882.4]
  wire  valid_11_30; // @[Switch.scala 30:36:@1883.4]
  wire  _T_6974; // @[Switch.scala 30:53:@1885.4]
  wire  valid_11_31; // @[Switch.scala 30:36:@1886.4]
  wire [4:0] _T_7008; // @[Mux.scala 31:69:@1888.4]
  wire [4:0] _T_7009; // @[Mux.scala 31:69:@1889.4]
  wire [4:0] _T_7010; // @[Mux.scala 31:69:@1890.4]
  wire [4:0] _T_7011; // @[Mux.scala 31:69:@1891.4]
  wire [4:0] _T_7012; // @[Mux.scala 31:69:@1892.4]
  wire [4:0] _T_7013; // @[Mux.scala 31:69:@1893.4]
  wire [4:0] _T_7014; // @[Mux.scala 31:69:@1894.4]
  wire [4:0] _T_7015; // @[Mux.scala 31:69:@1895.4]
  wire [4:0] _T_7016; // @[Mux.scala 31:69:@1896.4]
  wire [4:0] _T_7017; // @[Mux.scala 31:69:@1897.4]
  wire [4:0] _T_7018; // @[Mux.scala 31:69:@1898.4]
  wire [4:0] _T_7019; // @[Mux.scala 31:69:@1899.4]
  wire [4:0] _T_7020; // @[Mux.scala 31:69:@1900.4]
  wire [4:0] _T_7021; // @[Mux.scala 31:69:@1901.4]
  wire [4:0] _T_7022; // @[Mux.scala 31:69:@1902.4]
  wire [4:0] _T_7023; // @[Mux.scala 31:69:@1903.4]
  wire [4:0] _T_7024; // @[Mux.scala 31:69:@1904.4]
  wire [4:0] _T_7025; // @[Mux.scala 31:69:@1905.4]
  wire [4:0] _T_7026; // @[Mux.scala 31:69:@1906.4]
  wire [4:0] _T_7027; // @[Mux.scala 31:69:@1907.4]
  wire [4:0] _T_7028; // @[Mux.scala 31:69:@1908.4]
  wire [4:0] _T_7029; // @[Mux.scala 31:69:@1909.4]
  wire [4:0] _T_7030; // @[Mux.scala 31:69:@1910.4]
  wire [4:0] _T_7031; // @[Mux.scala 31:69:@1911.4]
  wire [4:0] _T_7032; // @[Mux.scala 31:69:@1912.4]
  wire [4:0] _T_7033; // @[Mux.scala 31:69:@1913.4]
  wire [4:0] _T_7034; // @[Mux.scala 31:69:@1914.4]
  wire [4:0] _T_7035; // @[Mux.scala 31:69:@1915.4]
  wire [4:0] _T_7036; // @[Mux.scala 31:69:@1916.4]
  wire [4:0] _T_7037; // @[Mux.scala 31:69:@1917.4]
  wire [4:0] select_11; // @[Mux.scala 31:69:@1918.4]
  wire [47:0] _GEN_353; // @[Switch.scala 33:19:@1920.4]
  wire [47:0] _GEN_354; // @[Switch.scala 33:19:@1920.4]
  wire [47:0] _GEN_355; // @[Switch.scala 33:19:@1920.4]
  wire [47:0] _GEN_356; // @[Switch.scala 33:19:@1920.4]
  wire [47:0] _GEN_357; // @[Switch.scala 33:19:@1920.4]
  wire [47:0] _GEN_358; // @[Switch.scala 33:19:@1920.4]
  wire [47:0] _GEN_359; // @[Switch.scala 33:19:@1920.4]
  wire [47:0] _GEN_360; // @[Switch.scala 33:19:@1920.4]
  wire [47:0] _GEN_361; // @[Switch.scala 33:19:@1920.4]
  wire [47:0] _GEN_362; // @[Switch.scala 33:19:@1920.4]
  wire [47:0] _GEN_363; // @[Switch.scala 33:19:@1920.4]
  wire [47:0] _GEN_364; // @[Switch.scala 33:19:@1920.4]
  wire [47:0] _GEN_365; // @[Switch.scala 33:19:@1920.4]
  wire [47:0] _GEN_366; // @[Switch.scala 33:19:@1920.4]
  wire [47:0] _GEN_367; // @[Switch.scala 33:19:@1920.4]
  wire [47:0] _GEN_368; // @[Switch.scala 33:19:@1920.4]
  wire [47:0] _GEN_369; // @[Switch.scala 33:19:@1920.4]
  wire [47:0] _GEN_370; // @[Switch.scala 33:19:@1920.4]
  wire [47:0] _GEN_371; // @[Switch.scala 33:19:@1920.4]
  wire [47:0] _GEN_372; // @[Switch.scala 33:19:@1920.4]
  wire [47:0] _GEN_373; // @[Switch.scala 33:19:@1920.4]
  wire [47:0] _GEN_374; // @[Switch.scala 33:19:@1920.4]
  wire [47:0] _GEN_375; // @[Switch.scala 33:19:@1920.4]
  wire [47:0] _GEN_376; // @[Switch.scala 33:19:@1920.4]
  wire [47:0] _GEN_377; // @[Switch.scala 33:19:@1920.4]
  wire [47:0] _GEN_378; // @[Switch.scala 33:19:@1920.4]
  wire [47:0] _GEN_379; // @[Switch.scala 33:19:@1920.4]
  wire [47:0] _GEN_380; // @[Switch.scala 33:19:@1920.4]
  wire [47:0] _GEN_381; // @[Switch.scala 33:19:@1920.4]
  wire [47:0] _GEN_382; // @[Switch.scala 33:19:@1920.4]
  wire [7:0] _T_7046; // @[Switch.scala 34:32:@1927.4]
  wire [15:0] _T_7054; // @[Switch.scala 34:32:@1935.4]
  wire [7:0] _T_7061; // @[Switch.scala 34:32:@1942.4]
  wire [31:0] _T_7070; // @[Switch.scala 34:32:@1951.4]
  wire  _T_7074; // @[Switch.scala 30:53:@1954.4]
  wire  valid_12_0; // @[Switch.scala 30:36:@1955.4]
  wire  _T_7077; // @[Switch.scala 30:53:@1957.4]
  wire  valid_12_1; // @[Switch.scala 30:36:@1958.4]
  wire  _T_7080; // @[Switch.scala 30:53:@1960.4]
  wire  valid_12_2; // @[Switch.scala 30:36:@1961.4]
  wire  _T_7083; // @[Switch.scala 30:53:@1963.4]
  wire  valid_12_3; // @[Switch.scala 30:36:@1964.4]
  wire  _T_7086; // @[Switch.scala 30:53:@1966.4]
  wire  valid_12_4; // @[Switch.scala 30:36:@1967.4]
  wire  _T_7089; // @[Switch.scala 30:53:@1969.4]
  wire  valid_12_5; // @[Switch.scala 30:36:@1970.4]
  wire  _T_7092; // @[Switch.scala 30:53:@1972.4]
  wire  valid_12_6; // @[Switch.scala 30:36:@1973.4]
  wire  _T_7095; // @[Switch.scala 30:53:@1975.4]
  wire  valid_12_7; // @[Switch.scala 30:36:@1976.4]
  wire  _T_7098; // @[Switch.scala 30:53:@1978.4]
  wire  valid_12_8; // @[Switch.scala 30:36:@1979.4]
  wire  _T_7101; // @[Switch.scala 30:53:@1981.4]
  wire  valid_12_9; // @[Switch.scala 30:36:@1982.4]
  wire  _T_7104; // @[Switch.scala 30:53:@1984.4]
  wire  valid_12_10; // @[Switch.scala 30:36:@1985.4]
  wire  _T_7107; // @[Switch.scala 30:53:@1987.4]
  wire  valid_12_11; // @[Switch.scala 30:36:@1988.4]
  wire  _T_7110; // @[Switch.scala 30:53:@1990.4]
  wire  valid_12_12; // @[Switch.scala 30:36:@1991.4]
  wire  _T_7113; // @[Switch.scala 30:53:@1993.4]
  wire  valid_12_13; // @[Switch.scala 30:36:@1994.4]
  wire  _T_7116; // @[Switch.scala 30:53:@1996.4]
  wire  valid_12_14; // @[Switch.scala 30:36:@1997.4]
  wire  _T_7119; // @[Switch.scala 30:53:@1999.4]
  wire  valid_12_15; // @[Switch.scala 30:36:@2000.4]
  wire  _T_7122; // @[Switch.scala 30:53:@2002.4]
  wire  valid_12_16; // @[Switch.scala 30:36:@2003.4]
  wire  _T_7125; // @[Switch.scala 30:53:@2005.4]
  wire  valid_12_17; // @[Switch.scala 30:36:@2006.4]
  wire  _T_7128; // @[Switch.scala 30:53:@2008.4]
  wire  valid_12_18; // @[Switch.scala 30:36:@2009.4]
  wire  _T_7131; // @[Switch.scala 30:53:@2011.4]
  wire  valid_12_19; // @[Switch.scala 30:36:@2012.4]
  wire  _T_7134; // @[Switch.scala 30:53:@2014.4]
  wire  valid_12_20; // @[Switch.scala 30:36:@2015.4]
  wire  _T_7137; // @[Switch.scala 30:53:@2017.4]
  wire  valid_12_21; // @[Switch.scala 30:36:@2018.4]
  wire  _T_7140; // @[Switch.scala 30:53:@2020.4]
  wire  valid_12_22; // @[Switch.scala 30:36:@2021.4]
  wire  _T_7143; // @[Switch.scala 30:53:@2023.4]
  wire  valid_12_23; // @[Switch.scala 30:36:@2024.4]
  wire  _T_7146; // @[Switch.scala 30:53:@2026.4]
  wire  valid_12_24; // @[Switch.scala 30:36:@2027.4]
  wire  _T_7149; // @[Switch.scala 30:53:@2029.4]
  wire  valid_12_25; // @[Switch.scala 30:36:@2030.4]
  wire  _T_7152; // @[Switch.scala 30:53:@2032.4]
  wire  valid_12_26; // @[Switch.scala 30:36:@2033.4]
  wire  _T_7155; // @[Switch.scala 30:53:@2035.4]
  wire  valid_12_27; // @[Switch.scala 30:36:@2036.4]
  wire  _T_7158; // @[Switch.scala 30:53:@2038.4]
  wire  valid_12_28; // @[Switch.scala 30:36:@2039.4]
  wire  _T_7161; // @[Switch.scala 30:53:@2041.4]
  wire  valid_12_29; // @[Switch.scala 30:36:@2042.4]
  wire  _T_7164; // @[Switch.scala 30:53:@2044.4]
  wire  valid_12_30; // @[Switch.scala 30:36:@2045.4]
  wire  _T_7167; // @[Switch.scala 30:53:@2047.4]
  wire  valid_12_31; // @[Switch.scala 30:36:@2048.4]
  wire [4:0] _T_7201; // @[Mux.scala 31:69:@2050.4]
  wire [4:0] _T_7202; // @[Mux.scala 31:69:@2051.4]
  wire [4:0] _T_7203; // @[Mux.scala 31:69:@2052.4]
  wire [4:0] _T_7204; // @[Mux.scala 31:69:@2053.4]
  wire [4:0] _T_7205; // @[Mux.scala 31:69:@2054.4]
  wire [4:0] _T_7206; // @[Mux.scala 31:69:@2055.4]
  wire [4:0] _T_7207; // @[Mux.scala 31:69:@2056.4]
  wire [4:0] _T_7208; // @[Mux.scala 31:69:@2057.4]
  wire [4:0] _T_7209; // @[Mux.scala 31:69:@2058.4]
  wire [4:0] _T_7210; // @[Mux.scala 31:69:@2059.4]
  wire [4:0] _T_7211; // @[Mux.scala 31:69:@2060.4]
  wire [4:0] _T_7212; // @[Mux.scala 31:69:@2061.4]
  wire [4:0] _T_7213; // @[Mux.scala 31:69:@2062.4]
  wire [4:0] _T_7214; // @[Mux.scala 31:69:@2063.4]
  wire [4:0] _T_7215; // @[Mux.scala 31:69:@2064.4]
  wire [4:0] _T_7216; // @[Mux.scala 31:69:@2065.4]
  wire [4:0] _T_7217; // @[Mux.scala 31:69:@2066.4]
  wire [4:0] _T_7218; // @[Mux.scala 31:69:@2067.4]
  wire [4:0] _T_7219; // @[Mux.scala 31:69:@2068.4]
  wire [4:0] _T_7220; // @[Mux.scala 31:69:@2069.4]
  wire [4:0] _T_7221; // @[Mux.scala 31:69:@2070.4]
  wire [4:0] _T_7222; // @[Mux.scala 31:69:@2071.4]
  wire [4:0] _T_7223; // @[Mux.scala 31:69:@2072.4]
  wire [4:0] _T_7224; // @[Mux.scala 31:69:@2073.4]
  wire [4:0] _T_7225; // @[Mux.scala 31:69:@2074.4]
  wire [4:0] _T_7226; // @[Mux.scala 31:69:@2075.4]
  wire [4:0] _T_7227; // @[Mux.scala 31:69:@2076.4]
  wire [4:0] _T_7228; // @[Mux.scala 31:69:@2077.4]
  wire [4:0] _T_7229; // @[Mux.scala 31:69:@2078.4]
  wire [4:0] _T_7230; // @[Mux.scala 31:69:@2079.4]
  wire [4:0] select_12; // @[Mux.scala 31:69:@2080.4]
  wire [47:0] _GEN_385; // @[Switch.scala 33:19:@2082.4]
  wire [47:0] _GEN_386; // @[Switch.scala 33:19:@2082.4]
  wire [47:0] _GEN_387; // @[Switch.scala 33:19:@2082.4]
  wire [47:0] _GEN_388; // @[Switch.scala 33:19:@2082.4]
  wire [47:0] _GEN_389; // @[Switch.scala 33:19:@2082.4]
  wire [47:0] _GEN_390; // @[Switch.scala 33:19:@2082.4]
  wire [47:0] _GEN_391; // @[Switch.scala 33:19:@2082.4]
  wire [47:0] _GEN_392; // @[Switch.scala 33:19:@2082.4]
  wire [47:0] _GEN_393; // @[Switch.scala 33:19:@2082.4]
  wire [47:0] _GEN_394; // @[Switch.scala 33:19:@2082.4]
  wire [47:0] _GEN_395; // @[Switch.scala 33:19:@2082.4]
  wire [47:0] _GEN_396; // @[Switch.scala 33:19:@2082.4]
  wire [47:0] _GEN_397; // @[Switch.scala 33:19:@2082.4]
  wire [47:0] _GEN_398; // @[Switch.scala 33:19:@2082.4]
  wire [47:0] _GEN_399; // @[Switch.scala 33:19:@2082.4]
  wire [47:0] _GEN_400; // @[Switch.scala 33:19:@2082.4]
  wire [47:0] _GEN_401; // @[Switch.scala 33:19:@2082.4]
  wire [47:0] _GEN_402; // @[Switch.scala 33:19:@2082.4]
  wire [47:0] _GEN_403; // @[Switch.scala 33:19:@2082.4]
  wire [47:0] _GEN_404; // @[Switch.scala 33:19:@2082.4]
  wire [47:0] _GEN_405; // @[Switch.scala 33:19:@2082.4]
  wire [47:0] _GEN_406; // @[Switch.scala 33:19:@2082.4]
  wire [47:0] _GEN_407; // @[Switch.scala 33:19:@2082.4]
  wire [47:0] _GEN_408; // @[Switch.scala 33:19:@2082.4]
  wire [47:0] _GEN_409; // @[Switch.scala 33:19:@2082.4]
  wire [47:0] _GEN_410; // @[Switch.scala 33:19:@2082.4]
  wire [47:0] _GEN_411; // @[Switch.scala 33:19:@2082.4]
  wire [47:0] _GEN_412; // @[Switch.scala 33:19:@2082.4]
  wire [47:0] _GEN_413; // @[Switch.scala 33:19:@2082.4]
  wire [47:0] _GEN_414; // @[Switch.scala 33:19:@2082.4]
  wire [7:0] _T_7239; // @[Switch.scala 34:32:@2089.4]
  wire [15:0] _T_7247; // @[Switch.scala 34:32:@2097.4]
  wire [7:0] _T_7254; // @[Switch.scala 34:32:@2104.4]
  wire [31:0] _T_7263; // @[Switch.scala 34:32:@2113.4]
  wire  _T_7267; // @[Switch.scala 30:53:@2116.4]
  wire  valid_13_0; // @[Switch.scala 30:36:@2117.4]
  wire  _T_7270; // @[Switch.scala 30:53:@2119.4]
  wire  valid_13_1; // @[Switch.scala 30:36:@2120.4]
  wire  _T_7273; // @[Switch.scala 30:53:@2122.4]
  wire  valid_13_2; // @[Switch.scala 30:36:@2123.4]
  wire  _T_7276; // @[Switch.scala 30:53:@2125.4]
  wire  valid_13_3; // @[Switch.scala 30:36:@2126.4]
  wire  _T_7279; // @[Switch.scala 30:53:@2128.4]
  wire  valid_13_4; // @[Switch.scala 30:36:@2129.4]
  wire  _T_7282; // @[Switch.scala 30:53:@2131.4]
  wire  valid_13_5; // @[Switch.scala 30:36:@2132.4]
  wire  _T_7285; // @[Switch.scala 30:53:@2134.4]
  wire  valid_13_6; // @[Switch.scala 30:36:@2135.4]
  wire  _T_7288; // @[Switch.scala 30:53:@2137.4]
  wire  valid_13_7; // @[Switch.scala 30:36:@2138.4]
  wire  _T_7291; // @[Switch.scala 30:53:@2140.4]
  wire  valid_13_8; // @[Switch.scala 30:36:@2141.4]
  wire  _T_7294; // @[Switch.scala 30:53:@2143.4]
  wire  valid_13_9; // @[Switch.scala 30:36:@2144.4]
  wire  _T_7297; // @[Switch.scala 30:53:@2146.4]
  wire  valid_13_10; // @[Switch.scala 30:36:@2147.4]
  wire  _T_7300; // @[Switch.scala 30:53:@2149.4]
  wire  valid_13_11; // @[Switch.scala 30:36:@2150.4]
  wire  _T_7303; // @[Switch.scala 30:53:@2152.4]
  wire  valid_13_12; // @[Switch.scala 30:36:@2153.4]
  wire  _T_7306; // @[Switch.scala 30:53:@2155.4]
  wire  valid_13_13; // @[Switch.scala 30:36:@2156.4]
  wire  _T_7309; // @[Switch.scala 30:53:@2158.4]
  wire  valid_13_14; // @[Switch.scala 30:36:@2159.4]
  wire  _T_7312; // @[Switch.scala 30:53:@2161.4]
  wire  valid_13_15; // @[Switch.scala 30:36:@2162.4]
  wire  _T_7315; // @[Switch.scala 30:53:@2164.4]
  wire  valid_13_16; // @[Switch.scala 30:36:@2165.4]
  wire  _T_7318; // @[Switch.scala 30:53:@2167.4]
  wire  valid_13_17; // @[Switch.scala 30:36:@2168.4]
  wire  _T_7321; // @[Switch.scala 30:53:@2170.4]
  wire  valid_13_18; // @[Switch.scala 30:36:@2171.4]
  wire  _T_7324; // @[Switch.scala 30:53:@2173.4]
  wire  valid_13_19; // @[Switch.scala 30:36:@2174.4]
  wire  _T_7327; // @[Switch.scala 30:53:@2176.4]
  wire  valid_13_20; // @[Switch.scala 30:36:@2177.4]
  wire  _T_7330; // @[Switch.scala 30:53:@2179.4]
  wire  valid_13_21; // @[Switch.scala 30:36:@2180.4]
  wire  _T_7333; // @[Switch.scala 30:53:@2182.4]
  wire  valid_13_22; // @[Switch.scala 30:36:@2183.4]
  wire  _T_7336; // @[Switch.scala 30:53:@2185.4]
  wire  valid_13_23; // @[Switch.scala 30:36:@2186.4]
  wire  _T_7339; // @[Switch.scala 30:53:@2188.4]
  wire  valid_13_24; // @[Switch.scala 30:36:@2189.4]
  wire  _T_7342; // @[Switch.scala 30:53:@2191.4]
  wire  valid_13_25; // @[Switch.scala 30:36:@2192.4]
  wire  _T_7345; // @[Switch.scala 30:53:@2194.4]
  wire  valid_13_26; // @[Switch.scala 30:36:@2195.4]
  wire  _T_7348; // @[Switch.scala 30:53:@2197.4]
  wire  valid_13_27; // @[Switch.scala 30:36:@2198.4]
  wire  _T_7351; // @[Switch.scala 30:53:@2200.4]
  wire  valid_13_28; // @[Switch.scala 30:36:@2201.4]
  wire  _T_7354; // @[Switch.scala 30:53:@2203.4]
  wire  valid_13_29; // @[Switch.scala 30:36:@2204.4]
  wire  _T_7357; // @[Switch.scala 30:53:@2206.4]
  wire  valid_13_30; // @[Switch.scala 30:36:@2207.4]
  wire  _T_7360; // @[Switch.scala 30:53:@2209.4]
  wire  valid_13_31; // @[Switch.scala 30:36:@2210.4]
  wire [4:0] _T_7394; // @[Mux.scala 31:69:@2212.4]
  wire [4:0] _T_7395; // @[Mux.scala 31:69:@2213.4]
  wire [4:0] _T_7396; // @[Mux.scala 31:69:@2214.4]
  wire [4:0] _T_7397; // @[Mux.scala 31:69:@2215.4]
  wire [4:0] _T_7398; // @[Mux.scala 31:69:@2216.4]
  wire [4:0] _T_7399; // @[Mux.scala 31:69:@2217.4]
  wire [4:0] _T_7400; // @[Mux.scala 31:69:@2218.4]
  wire [4:0] _T_7401; // @[Mux.scala 31:69:@2219.4]
  wire [4:0] _T_7402; // @[Mux.scala 31:69:@2220.4]
  wire [4:0] _T_7403; // @[Mux.scala 31:69:@2221.4]
  wire [4:0] _T_7404; // @[Mux.scala 31:69:@2222.4]
  wire [4:0] _T_7405; // @[Mux.scala 31:69:@2223.4]
  wire [4:0] _T_7406; // @[Mux.scala 31:69:@2224.4]
  wire [4:0] _T_7407; // @[Mux.scala 31:69:@2225.4]
  wire [4:0] _T_7408; // @[Mux.scala 31:69:@2226.4]
  wire [4:0] _T_7409; // @[Mux.scala 31:69:@2227.4]
  wire [4:0] _T_7410; // @[Mux.scala 31:69:@2228.4]
  wire [4:0] _T_7411; // @[Mux.scala 31:69:@2229.4]
  wire [4:0] _T_7412; // @[Mux.scala 31:69:@2230.4]
  wire [4:0] _T_7413; // @[Mux.scala 31:69:@2231.4]
  wire [4:0] _T_7414; // @[Mux.scala 31:69:@2232.4]
  wire [4:0] _T_7415; // @[Mux.scala 31:69:@2233.4]
  wire [4:0] _T_7416; // @[Mux.scala 31:69:@2234.4]
  wire [4:0] _T_7417; // @[Mux.scala 31:69:@2235.4]
  wire [4:0] _T_7418; // @[Mux.scala 31:69:@2236.4]
  wire [4:0] _T_7419; // @[Mux.scala 31:69:@2237.4]
  wire [4:0] _T_7420; // @[Mux.scala 31:69:@2238.4]
  wire [4:0] _T_7421; // @[Mux.scala 31:69:@2239.4]
  wire [4:0] _T_7422; // @[Mux.scala 31:69:@2240.4]
  wire [4:0] _T_7423; // @[Mux.scala 31:69:@2241.4]
  wire [4:0] select_13; // @[Mux.scala 31:69:@2242.4]
  wire [47:0] _GEN_417; // @[Switch.scala 33:19:@2244.4]
  wire [47:0] _GEN_418; // @[Switch.scala 33:19:@2244.4]
  wire [47:0] _GEN_419; // @[Switch.scala 33:19:@2244.4]
  wire [47:0] _GEN_420; // @[Switch.scala 33:19:@2244.4]
  wire [47:0] _GEN_421; // @[Switch.scala 33:19:@2244.4]
  wire [47:0] _GEN_422; // @[Switch.scala 33:19:@2244.4]
  wire [47:0] _GEN_423; // @[Switch.scala 33:19:@2244.4]
  wire [47:0] _GEN_424; // @[Switch.scala 33:19:@2244.4]
  wire [47:0] _GEN_425; // @[Switch.scala 33:19:@2244.4]
  wire [47:0] _GEN_426; // @[Switch.scala 33:19:@2244.4]
  wire [47:0] _GEN_427; // @[Switch.scala 33:19:@2244.4]
  wire [47:0] _GEN_428; // @[Switch.scala 33:19:@2244.4]
  wire [47:0] _GEN_429; // @[Switch.scala 33:19:@2244.4]
  wire [47:0] _GEN_430; // @[Switch.scala 33:19:@2244.4]
  wire [47:0] _GEN_431; // @[Switch.scala 33:19:@2244.4]
  wire [47:0] _GEN_432; // @[Switch.scala 33:19:@2244.4]
  wire [47:0] _GEN_433; // @[Switch.scala 33:19:@2244.4]
  wire [47:0] _GEN_434; // @[Switch.scala 33:19:@2244.4]
  wire [47:0] _GEN_435; // @[Switch.scala 33:19:@2244.4]
  wire [47:0] _GEN_436; // @[Switch.scala 33:19:@2244.4]
  wire [47:0] _GEN_437; // @[Switch.scala 33:19:@2244.4]
  wire [47:0] _GEN_438; // @[Switch.scala 33:19:@2244.4]
  wire [47:0] _GEN_439; // @[Switch.scala 33:19:@2244.4]
  wire [47:0] _GEN_440; // @[Switch.scala 33:19:@2244.4]
  wire [47:0] _GEN_441; // @[Switch.scala 33:19:@2244.4]
  wire [47:0] _GEN_442; // @[Switch.scala 33:19:@2244.4]
  wire [47:0] _GEN_443; // @[Switch.scala 33:19:@2244.4]
  wire [47:0] _GEN_444; // @[Switch.scala 33:19:@2244.4]
  wire [47:0] _GEN_445; // @[Switch.scala 33:19:@2244.4]
  wire [47:0] _GEN_446; // @[Switch.scala 33:19:@2244.4]
  wire [7:0] _T_7432; // @[Switch.scala 34:32:@2251.4]
  wire [15:0] _T_7440; // @[Switch.scala 34:32:@2259.4]
  wire [7:0] _T_7447; // @[Switch.scala 34:32:@2266.4]
  wire [31:0] _T_7456; // @[Switch.scala 34:32:@2275.4]
  wire  _T_7460; // @[Switch.scala 30:53:@2278.4]
  wire  valid_14_0; // @[Switch.scala 30:36:@2279.4]
  wire  _T_7463; // @[Switch.scala 30:53:@2281.4]
  wire  valid_14_1; // @[Switch.scala 30:36:@2282.4]
  wire  _T_7466; // @[Switch.scala 30:53:@2284.4]
  wire  valid_14_2; // @[Switch.scala 30:36:@2285.4]
  wire  _T_7469; // @[Switch.scala 30:53:@2287.4]
  wire  valid_14_3; // @[Switch.scala 30:36:@2288.4]
  wire  _T_7472; // @[Switch.scala 30:53:@2290.4]
  wire  valid_14_4; // @[Switch.scala 30:36:@2291.4]
  wire  _T_7475; // @[Switch.scala 30:53:@2293.4]
  wire  valid_14_5; // @[Switch.scala 30:36:@2294.4]
  wire  _T_7478; // @[Switch.scala 30:53:@2296.4]
  wire  valid_14_6; // @[Switch.scala 30:36:@2297.4]
  wire  _T_7481; // @[Switch.scala 30:53:@2299.4]
  wire  valid_14_7; // @[Switch.scala 30:36:@2300.4]
  wire  _T_7484; // @[Switch.scala 30:53:@2302.4]
  wire  valid_14_8; // @[Switch.scala 30:36:@2303.4]
  wire  _T_7487; // @[Switch.scala 30:53:@2305.4]
  wire  valid_14_9; // @[Switch.scala 30:36:@2306.4]
  wire  _T_7490; // @[Switch.scala 30:53:@2308.4]
  wire  valid_14_10; // @[Switch.scala 30:36:@2309.4]
  wire  _T_7493; // @[Switch.scala 30:53:@2311.4]
  wire  valid_14_11; // @[Switch.scala 30:36:@2312.4]
  wire  _T_7496; // @[Switch.scala 30:53:@2314.4]
  wire  valid_14_12; // @[Switch.scala 30:36:@2315.4]
  wire  _T_7499; // @[Switch.scala 30:53:@2317.4]
  wire  valid_14_13; // @[Switch.scala 30:36:@2318.4]
  wire  _T_7502; // @[Switch.scala 30:53:@2320.4]
  wire  valid_14_14; // @[Switch.scala 30:36:@2321.4]
  wire  _T_7505; // @[Switch.scala 30:53:@2323.4]
  wire  valid_14_15; // @[Switch.scala 30:36:@2324.4]
  wire  _T_7508; // @[Switch.scala 30:53:@2326.4]
  wire  valid_14_16; // @[Switch.scala 30:36:@2327.4]
  wire  _T_7511; // @[Switch.scala 30:53:@2329.4]
  wire  valid_14_17; // @[Switch.scala 30:36:@2330.4]
  wire  _T_7514; // @[Switch.scala 30:53:@2332.4]
  wire  valid_14_18; // @[Switch.scala 30:36:@2333.4]
  wire  _T_7517; // @[Switch.scala 30:53:@2335.4]
  wire  valid_14_19; // @[Switch.scala 30:36:@2336.4]
  wire  _T_7520; // @[Switch.scala 30:53:@2338.4]
  wire  valid_14_20; // @[Switch.scala 30:36:@2339.4]
  wire  _T_7523; // @[Switch.scala 30:53:@2341.4]
  wire  valid_14_21; // @[Switch.scala 30:36:@2342.4]
  wire  _T_7526; // @[Switch.scala 30:53:@2344.4]
  wire  valid_14_22; // @[Switch.scala 30:36:@2345.4]
  wire  _T_7529; // @[Switch.scala 30:53:@2347.4]
  wire  valid_14_23; // @[Switch.scala 30:36:@2348.4]
  wire  _T_7532; // @[Switch.scala 30:53:@2350.4]
  wire  valid_14_24; // @[Switch.scala 30:36:@2351.4]
  wire  _T_7535; // @[Switch.scala 30:53:@2353.4]
  wire  valid_14_25; // @[Switch.scala 30:36:@2354.4]
  wire  _T_7538; // @[Switch.scala 30:53:@2356.4]
  wire  valid_14_26; // @[Switch.scala 30:36:@2357.4]
  wire  _T_7541; // @[Switch.scala 30:53:@2359.4]
  wire  valid_14_27; // @[Switch.scala 30:36:@2360.4]
  wire  _T_7544; // @[Switch.scala 30:53:@2362.4]
  wire  valid_14_28; // @[Switch.scala 30:36:@2363.4]
  wire  _T_7547; // @[Switch.scala 30:53:@2365.4]
  wire  valid_14_29; // @[Switch.scala 30:36:@2366.4]
  wire  _T_7550; // @[Switch.scala 30:53:@2368.4]
  wire  valid_14_30; // @[Switch.scala 30:36:@2369.4]
  wire  _T_7553; // @[Switch.scala 30:53:@2371.4]
  wire  valid_14_31; // @[Switch.scala 30:36:@2372.4]
  wire [4:0] _T_7587; // @[Mux.scala 31:69:@2374.4]
  wire [4:0] _T_7588; // @[Mux.scala 31:69:@2375.4]
  wire [4:0] _T_7589; // @[Mux.scala 31:69:@2376.4]
  wire [4:0] _T_7590; // @[Mux.scala 31:69:@2377.4]
  wire [4:0] _T_7591; // @[Mux.scala 31:69:@2378.4]
  wire [4:0] _T_7592; // @[Mux.scala 31:69:@2379.4]
  wire [4:0] _T_7593; // @[Mux.scala 31:69:@2380.4]
  wire [4:0] _T_7594; // @[Mux.scala 31:69:@2381.4]
  wire [4:0] _T_7595; // @[Mux.scala 31:69:@2382.4]
  wire [4:0] _T_7596; // @[Mux.scala 31:69:@2383.4]
  wire [4:0] _T_7597; // @[Mux.scala 31:69:@2384.4]
  wire [4:0] _T_7598; // @[Mux.scala 31:69:@2385.4]
  wire [4:0] _T_7599; // @[Mux.scala 31:69:@2386.4]
  wire [4:0] _T_7600; // @[Mux.scala 31:69:@2387.4]
  wire [4:0] _T_7601; // @[Mux.scala 31:69:@2388.4]
  wire [4:0] _T_7602; // @[Mux.scala 31:69:@2389.4]
  wire [4:0] _T_7603; // @[Mux.scala 31:69:@2390.4]
  wire [4:0] _T_7604; // @[Mux.scala 31:69:@2391.4]
  wire [4:0] _T_7605; // @[Mux.scala 31:69:@2392.4]
  wire [4:0] _T_7606; // @[Mux.scala 31:69:@2393.4]
  wire [4:0] _T_7607; // @[Mux.scala 31:69:@2394.4]
  wire [4:0] _T_7608; // @[Mux.scala 31:69:@2395.4]
  wire [4:0] _T_7609; // @[Mux.scala 31:69:@2396.4]
  wire [4:0] _T_7610; // @[Mux.scala 31:69:@2397.4]
  wire [4:0] _T_7611; // @[Mux.scala 31:69:@2398.4]
  wire [4:0] _T_7612; // @[Mux.scala 31:69:@2399.4]
  wire [4:0] _T_7613; // @[Mux.scala 31:69:@2400.4]
  wire [4:0] _T_7614; // @[Mux.scala 31:69:@2401.4]
  wire [4:0] _T_7615; // @[Mux.scala 31:69:@2402.4]
  wire [4:0] _T_7616; // @[Mux.scala 31:69:@2403.4]
  wire [4:0] select_14; // @[Mux.scala 31:69:@2404.4]
  wire [47:0] _GEN_449; // @[Switch.scala 33:19:@2406.4]
  wire [47:0] _GEN_450; // @[Switch.scala 33:19:@2406.4]
  wire [47:0] _GEN_451; // @[Switch.scala 33:19:@2406.4]
  wire [47:0] _GEN_452; // @[Switch.scala 33:19:@2406.4]
  wire [47:0] _GEN_453; // @[Switch.scala 33:19:@2406.4]
  wire [47:0] _GEN_454; // @[Switch.scala 33:19:@2406.4]
  wire [47:0] _GEN_455; // @[Switch.scala 33:19:@2406.4]
  wire [47:0] _GEN_456; // @[Switch.scala 33:19:@2406.4]
  wire [47:0] _GEN_457; // @[Switch.scala 33:19:@2406.4]
  wire [47:0] _GEN_458; // @[Switch.scala 33:19:@2406.4]
  wire [47:0] _GEN_459; // @[Switch.scala 33:19:@2406.4]
  wire [47:0] _GEN_460; // @[Switch.scala 33:19:@2406.4]
  wire [47:0] _GEN_461; // @[Switch.scala 33:19:@2406.4]
  wire [47:0] _GEN_462; // @[Switch.scala 33:19:@2406.4]
  wire [47:0] _GEN_463; // @[Switch.scala 33:19:@2406.4]
  wire [47:0] _GEN_464; // @[Switch.scala 33:19:@2406.4]
  wire [47:0] _GEN_465; // @[Switch.scala 33:19:@2406.4]
  wire [47:0] _GEN_466; // @[Switch.scala 33:19:@2406.4]
  wire [47:0] _GEN_467; // @[Switch.scala 33:19:@2406.4]
  wire [47:0] _GEN_468; // @[Switch.scala 33:19:@2406.4]
  wire [47:0] _GEN_469; // @[Switch.scala 33:19:@2406.4]
  wire [47:0] _GEN_470; // @[Switch.scala 33:19:@2406.4]
  wire [47:0] _GEN_471; // @[Switch.scala 33:19:@2406.4]
  wire [47:0] _GEN_472; // @[Switch.scala 33:19:@2406.4]
  wire [47:0] _GEN_473; // @[Switch.scala 33:19:@2406.4]
  wire [47:0] _GEN_474; // @[Switch.scala 33:19:@2406.4]
  wire [47:0] _GEN_475; // @[Switch.scala 33:19:@2406.4]
  wire [47:0] _GEN_476; // @[Switch.scala 33:19:@2406.4]
  wire [47:0] _GEN_477; // @[Switch.scala 33:19:@2406.4]
  wire [47:0] _GEN_478; // @[Switch.scala 33:19:@2406.4]
  wire [7:0] _T_7625; // @[Switch.scala 34:32:@2413.4]
  wire [15:0] _T_7633; // @[Switch.scala 34:32:@2421.4]
  wire [7:0] _T_7640; // @[Switch.scala 34:32:@2428.4]
  wire [31:0] _T_7649; // @[Switch.scala 34:32:@2437.4]
  wire  _T_7653; // @[Switch.scala 30:53:@2440.4]
  wire  valid_15_0; // @[Switch.scala 30:36:@2441.4]
  wire  _T_7656; // @[Switch.scala 30:53:@2443.4]
  wire  valid_15_1; // @[Switch.scala 30:36:@2444.4]
  wire  _T_7659; // @[Switch.scala 30:53:@2446.4]
  wire  valid_15_2; // @[Switch.scala 30:36:@2447.4]
  wire  _T_7662; // @[Switch.scala 30:53:@2449.4]
  wire  valid_15_3; // @[Switch.scala 30:36:@2450.4]
  wire  _T_7665; // @[Switch.scala 30:53:@2452.4]
  wire  valid_15_4; // @[Switch.scala 30:36:@2453.4]
  wire  _T_7668; // @[Switch.scala 30:53:@2455.4]
  wire  valid_15_5; // @[Switch.scala 30:36:@2456.4]
  wire  _T_7671; // @[Switch.scala 30:53:@2458.4]
  wire  valid_15_6; // @[Switch.scala 30:36:@2459.4]
  wire  _T_7674; // @[Switch.scala 30:53:@2461.4]
  wire  valid_15_7; // @[Switch.scala 30:36:@2462.4]
  wire  _T_7677; // @[Switch.scala 30:53:@2464.4]
  wire  valid_15_8; // @[Switch.scala 30:36:@2465.4]
  wire  _T_7680; // @[Switch.scala 30:53:@2467.4]
  wire  valid_15_9; // @[Switch.scala 30:36:@2468.4]
  wire  _T_7683; // @[Switch.scala 30:53:@2470.4]
  wire  valid_15_10; // @[Switch.scala 30:36:@2471.4]
  wire  _T_7686; // @[Switch.scala 30:53:@2473.4]
  wire  valid_15_11; // @[Switch.scala 30:36:@2474.4]
  wire  _T_7689; // @[Switch.scala 30:53:@2476.4]
  wire  valid_15_12; // @[Switch.scala 30:36:@2477.4]
  wire  _T_7692; // @[Switch.scala 30:53:@2479.4]
  wire  valid_15_13; // @[Switch.scala 30:36:@2480.4]
  wire  _T_7695; // @[Switch.scala 30:53:@2482.4]
  wire  valid_15_14; // @[Switch.scala 30:36:@2483.4]
  wire  _T_7698; // @[Switch.scala 30:53:@2485.4]
  wire  valid_15_15; // @[Switch.scala 30:36:@2486.4]
  wire  _T_7701; // @[Switch.scala 30:53:@2488.4]
  wire  valid_15_16; // @[Switch.scala 30:36:@2489.4]
  wire  _T_7704; // @[Switch.scala 30:53:@2491.4]
  wire  valid_15_17; // @[Switch.scala 30:36:@2492.4]
  wire  _T_7707; // @[Switch.scala 30:53:@2494.4]
  wire  valid_15_18; // @[Switch.scala 30:36:@2495.4]
  wire  _T_7710; // @[Switch.scala 30:53:@2497.4]
  wire  valid_15_19; // @[Switch.scala 30:36:@2498.4]
  wire  _T_7713; // @[Switch.scala 30:53:@2500.4]
  wire  valid_15_20; // @[Switch.scala 30:36:@2501.4]
  wire  _T_7716; // @[Switch.scala 30:53:@2503.4]
  wire  valid_15_21; // @[Switch.scala 30:36:@2504.4]
  wire  _T_7719; // @[Switch.scala 30:53:@2506.4]
  wire  valid_15_22; // @[Switch.scala 30:36:@2507.4]
  wire  _T_7722; // @[Switch.scala 30:53:@2509.4]
  wire  valid_15_23; // @[Switch.scala 30:36:@2510.4]
  wire  _T_7725; // @[Switch.scala 30:53:@2512.4]
  wire  valid_15_24; // @[Switch.scala 30:36:@2513.4]
  wire  _T_7728; // @[Switch.scala 30:53:@2515.4]
  wire  valid_15_25; // @[Switch.scala 30:36:@2516.4]
  wire  _T_7731; // @[Switch.scala 30:53:@2518.4]
  wire  valid_15_26; // @[Switch.scala 30:36:@2519.4]
  wire  _T_7734; // @[Switch.scala 30:53:@2521.4]
  wire  valid_15_27; // @[Switch.scala 30:36:@2522.4]
  wire  _T_7737; // @[Switch.scala 30:53:@2524.4]
  wire  valid_15_28; // @[Switch.scala 30:36:@2525.4]
  wire  _T_7740; // @[Switch.scala 30:53:@2527.4]
  wire  valid_15_29; // @[Switch.scala 30:36:@2528.4]
  wire  _T_7743; // @[Switch.scala 30:53:@2530.4]
  wire  valid_15_30; // @[Switch.scala 30:36:@2531.4]
  wire  _T_7746; // @[Switch.scala 30:53:@2533.4]
  wire  valid_15_31; // @[Switch.scala 30:36:@2534.4]
  wire [4:0] _T_7780; // @[Mux.scala 31:69:@2536.4]
  wire [4:0] _T_7781; // @[Mux.scala 31:69:@2537.4]
  wire [4:0] _T_7782; // @[Mux.scala 31:69:@2538.4]
  wire [4:0] _T_7783; // @[Mux.scala 31:69:@2539.4]
  wire [4:0] _T_7784; // @[Mux.scala 31:69:@2540.4]
  wire [4:0] _T_7785; // @[Mux.scala 31:69:@2541.4]
  wire [4:0] _T_7786; // @[Mux.scala 31:69:@2542.4]
  wire [4:0] _T_7787; // @[Mux.scala 31:69:@2543.4]
  wire [4:0] _T_7788; // @[Mux.scala 31:69:@2544.4]
  wire [4:0] _T_7789; // @[Mux.scala 31:69:@2545.4]
  wire [4:0] _T_7790; // @[Mux.scala 31:69:@2546.4]
  wire [4:0] _T_7791; // @[Mux.scala 31:69:@2547.4]
  wire [4:0] _T_7792; // @[Mux.scala 31:69:@2548.4]
  wire [4:0] _T_7793; // @[Mux.scala 31:69:@2549.4]
  wire [4:0] _T_7794; // @[Mux.scala 31:69:@2550.4]
  wire [4:0] _T_7795; // @[Mux.scala 31:69:@2551.4]
  wire [4:0] _T_7796; // @[Mux.scala 31:69:@2552.4]
  wire [4:0] _T_7797; // @[Mux.scala 31:69:@2553.4]
  wire [4:0] _T_7798; // @[Mux.scala 31:69:@2554.4]
  wire [4:0] _T_7799; // @[Mux.scala 31:69:@2555.4]
  wire [4:0] _T_7800; // @[Mux.scala 31:69:@2556.4]
  wire [4:0] _T_7801; // @[Mux.scala 31:69:@2557.4]
  wire [4:0] _T_7802; // @[Mux.scala 31:69:@2558.4]
  wire [4:0] _T_7803; // @[Mux.scala 31:69:@2559.4]
  wire [4:0] _T_7804; // @[Mux.scala 31:69:@2560.4]
  wire [4:0] _T_7805; // @[Mux.scala 31:69:@2561.4]
  wire [4:0] _T_7806; // @[Mux.scala 31:69:@2562.4]
  wire [4:0] _T_7807; // @[Mux.scala 31:69:@2563.4]
  wire [4:0] _T_7808; // @[Mux.scala 31:69:@2564.4]
  wire [4:0] _T_7809; // @[Mux.scala 31:69:@2565.4]
  wire [4:0] select_15; // @[Mux.scala 31:69:@2566.4]
  wire [47:0] _GEN_481; // @[Switch.scala 33:19:@2568.4]
  wire [47:0] _GEN_482; // @[Switch.scala 33:19:@2568.4]
  wire [47:0] _GEN_483; // @[Switch.scala 33:19:@2568.4]
  wire [47:0] _GEN_484; // @[Switch.scala 33:19:@2568.4]
  wire [47:0] _GEN_485; // @[Switch.scala 33:19:@2568.4]
  wire [47:0] _GEN_486; // @[Switch.scala 33:19:@2568.4]
  wire [47:0] _GEN_487; // @[Switch.scala 33:19:@2568.4]
  wire [47:0] _GEN_488; // @[Switch.scala 33:19:@2568.4]
  wire [47:0] _GEN_489; // @[Switch.scala 33:19:@2568.4]
  wire [47:0] _GEN_490; // @[Switch.scala 33:19:@2568.4]
  wire [47:0] _GEN_491; // @[Switch.scala 33:19:@2568.4]
  wire [47:0] _GEN_492; // @[Switch.scala 33:19:@2568.4]
  wire [47:0] _GEN_493; // @[Switch.scala 33:19:@2568.4]
  wire [47:0] _GEN_494; // @[Switch.scala 33:19:@2568.4]
  wire [47:0] _GEN_495; // @[Switch.scala 33:19:@2568.4]
  wire [47:0] _GEN_496; // @[Switch.scala 33:19:@2568.4]
  wire [47:0] _GEN_497; // @[Switch.scala 33:19:@2568.4]
  wire [47:0] _GEN_498; // @[Switch.scala 33:19:@2568.4]
  wire [47:0] _GEN_499; // @[Switch.scala 33:19:@2568.4]
  wire [47:0] _GEN_500; // @[Switch.scala 33:19:@2568.4]
  wire [47:0] _GEN_501; // @[Switch.scala 33:19:@2568.4]
  wire [47:0] _GEN_502; // @[Switch.scala 33:19:@2568.4]
  wire [47:0] _GEN_503; // @[Switch.scala 33:19:@2568.4]
  wire [47:0] _GEN_504; // @[Switch.scala 33:19:@2568.4]
  wire [47:0] _GEN_505; // @[Switch.scala 33:19:@2568.4]
  wire [47:0] _GEN_506; // @[Switch.scala 33:19:@2568.4]
  wire [47:0] _GEN_507; // @[Switch.scala 33:19:@2568.4]
  wire [47:0] _GEN_508; // @[Switch.scala 33:19:@2568.4]
  wire [47:0] _GEN_509; // @[Switch.scala 33:19:@2568.4]
  wire [47:0] _GEN_510; // @[Switch.scala 33:19:@2568.4]
  wire [7:0] _T_7818; // @[Switch.scala 34:32:@2575.4]
  wire [15:0] _T_7826; // @[Switch.scala 34:32:@2583.4]
  wire [7:0] _T_7833; // @[Switch.scala 34:32:@2590.4]
  wire [31:0] _T_7842; // @[Switch.scala 34:32:@2599.4]
  wire  _T_7846; // @[Switch.scala 30:53:@2602.4]
  wire  valid_16_0; // @[Switch.scala 30:36:@2603.4]
  wire  _T_7849; // @[Switch.scala 30:53:@2605.4]
  wire  valid_16_1; // @[Switch.scala 30:36:@2606.4]
  wire  _T_7852; // @[Switch.scala 30:53:@2608.4]
  wire  valid_16_2; // @[Switch.scala 30:36:@2609.4]
  wire  _T_7855; // @[Switch.scala 30:53:@2611.4]
  wire  valid_16_3; // @[Switch.scala 30:36:@2612.4]
  wire  _T_7858; // @[Switch.scala 30:53:@2614.4]
  wire  valid_16_4; // @[Switch.scala 30:36:@2615.4]
  wire  _T_7861; // @[Switch.scala 30:53:@2617.4]
  wire  valid_16_5; // @[Switch.scala 30:36:@2618.4]
  wire  _T_7864; // @[Switch.scala 30:53:@2620.4]
  wire  valid_16_6; // @[Switch.scala 30:36:@2621.4]
  wire  _T_7867; // @[Switch.scala 30:53:@2623.4]
  wire  valid_16_7; // @[Switch.scala 30:36:@2624.4]
  wire  _T_7870; // @[Switch.scala 30:53:@2626.4]
  wire  valid_16_8; // @[Switch.scala 30:36:@2627.4]
  wire  _T_7873; // @[Switch.scala 30:53:@2629.4]
  wire  valid_16_9; // @[Switch.scala 30:36:@2630.4]
  wire  _T_7876; // @[Switch.scala 30:53:@2632.4]
  wire  valid_16_10; // @[Switch.scala 30:36:@2633.4]
  wire  _T_7879; // @[Switch.scala 30:53:@2635.4]
  wire  valid_16_11; // @[Switch.scala 30:36:@2636.4]
  wire  _T_7882; // @[Switch.scala 30:53:@2638.4]
  wire  valid_16_12; // @[Switch.scala 30:36:@2639.4]
  wire  _T_7885; // @[Switch.scala 30:53:@2641.4]
  wire  valid_16_13; // @[Switch.scala 30:36:@2642.4]
  wire  _T_7888; // @[Switch.scala 30:53:@2644.4]
  wire  valid_16_14; // @[Switch.scala 30:36:@2645.4]
  wire  _T_7891; // @[Switch.scala 30:53:@2647.4]
  wire  valid_16_15; // @[Switch.scala 30:36:@2648.4]
  wire  _T_7894; // @[Switch.scala 30:53:@2650.4]
  wire  valid_16_16; // @[Switch.scala 30:36:@2651.4]
  wire  _T_7897; // @[Switch.scala 30:53:@2653.4]
  wire  valid_16_17; // @[Switch.scala 30:36:@2654.4]
  wire  _T_7900; // @[Switch.scala 30:53:@2656.4]
  wire  valid_16_18; // @[Switch.scala 30:36:@2657.4]
  wire  _T_7903; // @[Switch.scala 30:53:@2659.4]
  wire  valid_16_19; // @[Switch.scala 30:36:@2660.4]
  wire  _T_7906; // @[Switch.scala 30:53:@2662.4]
  wire  valid_16_20; // @[Switch.scala 30:36:@2663.4]
  wire  _T_7909; // @[Switch.scala 30:53:@2665.4]
  wire  valid_16_21; // @[Switch.scala 30:36:@2666.4]
  wire  _T_7912; // @[Switch.scala 30:53:@2668.4]
  wire  valid_16_22; // @[Switch.scala 30:36:@2669.4]
  wire  _T_7915; // @[Switch.scala 30:53:@2671.4]
  wire  valid_16_23; // @[Switch.scala 30:36:@2672.4]
  wire  _T_7918; // @[Switch.scala 30:53:@2674.4]
  wire  valid_16_24; // @[Switch.scala 30:36:@2675.4]
  wire  _T_7921; // @[Switch.scala 30:53:@2677.4]
  wire  valid_16_25; // @[Switch.scala 30:36:@2678.4]
  wire  _T_7924; // @[Switch.scala 30:53:@2680.4]
  wire  valid_16_26; // @[Switch.scala 30:36:@2681.4]
  wire  _T_7927; // @[Switch.scala 30:53:@2683.4]
  wire  valid_16_27; // @[Switch.scala 30:36:@2684.4]
  wire  _T_7930; // @[Switch.scala 30:53:@2686.4]
  wire  valid_16_28; // @[Switch.scala 30:36:@2687.4]
  wire  _T_7933; // @[Switch.scala 30:53:@2689.4]
  wire  valid_16_29; // @[Switch.scala 30:36:@2690.4]
  wire  _T_7936; // @[Switch.scala 30:53:@2692.4]
  wire  valid_16_30; // @[Switch.scala 30:36:@2693.4]
  wire  _T_7939; // @[Switch.scala 30:53:@2695.4]
  wire  valid_16_31; // @[Switch.scala 30:36:@2696.4]
  wire [4:0] _T_7973; // @[Mux.scala 31:69:@2698.4]
  wire [4:0] _T_7974; // @[Mux.scala 31:69:@2699.4]
  wire [4:0] _T_7975; // @[Mux.scala 31:69:@2700.4]
  wire [4:0] _T_7976; // @[Mux.scala 31:69:@2701.4]
  wire [4:0] _T_7977; // @[Mux.scala 31:69:@2702.4]
  wire [4:0] _T_7978; // @[Mux.scala 31:69:@2703.4]
  wire [4:0] _T_7979; // @[Mux.scala 31:69:@2704.4]
  wire [4:0] _T_7980; // @[Mux.scala 31:69:@2705.4]
  wire [4:0] _T_7981; // @[Mux.scala 31:69:@2706.4]
  wire [4:0] _T_7982; // @[Mux.scala 31:69:@2707.4]
  wire [4:0] _T_7983; // @[Mux.scala 31:69:@2708.4]
  wire [4:0] _T_7984; // @[Mux.scala 31:69:@2709.4]
  wire [4:0] _T_7985; // @[Mux.scala 31:69:@2710.4]
  wire [4:0] _T_7986; // @[Mux.scala 31:69:@2711.4]
  wire [4:0] _T_7987; // @[Mux.scala 31:69:@2712.4]
  wire [4:0] _T_7988; // @[Mux.scala 31:69:@2713.4]
  wire [4:0] _T_7989; // @[Mux.scala 31:69:@2714.4]
  wire [4:0] _T_7990; // @[Mux.scala 31:69:@2715.4]
  wire [4:0] _T_7991; // @[Mux.scala 31:69:@2716.4]
  wire [4:0] _T_7992; // @[Mux.scala 31:69:@2717.4]
  wire [4:0] _T_7993; // @[Mux.scala 31:69:@2718.4]
  wire [4:0] _T_7994; // @[Mux.scala 31:69:@2719.4]
  wire [4:0] _T_7995; // @[Mux.scala 31:69:@2720.4]
  wire [4:0] _T_7996; // @[Mux.scala 31:69:@2721.4]
  wire [4:0] _T_7997; // @[Mux.scala 31:69:@2722.4]
  wire [4:0] _T_7998; // @[Mux.scala 31:69:@2723.4]
  wire [4:0] _T_7999; // @[Mux.scala 31:69:@2724.4]
  wire [4:0] _T_8000; // @[Mux.scala 31:69:@2725.4]
  wire [4:0] _T_8001; // @[Mux.scala 31:69:@2726.4]
  wire [4:0] _T_8002; // @[Mux.scala 31:69:@2727.4]
  wire [4:0] select_16; // @[Mux.scala 31:69:@2728.4]
  wire [47:0] _GEN_513; // @[Switch.scala 33:19:@2730.4]
  wire [47:0] _GEN_514; // @[Switch.scala 33:19:@2730.4]
  wire [47:0] _GEN_515; // @[Switch.scala 33:19:@2730.4]
  wire [47:0] _GEN_516; // @[Switch.scala 33:19:@2730.4]
  wire [47:0] _GEN_517; // @[Switch.scala 33:19:@2730.4]
  wire [47:0] _GEN_518; // @[Switch.scala 33:19:@2730.4]
  wire [47:0] _GEN_519; // @[Switch.scala 33:19:@2730.4]
  wire [47:0] _GEN_520; // @[Switch.scala 33:19:@2730.4]
  wire [47:0] _GEN_521; // @[Switch.scala 33:19:@2730.4]
  wire [47:0] _GEN_522; // @[Switch.scala 33:19:@2730.4]
  wire [47:0] _GEN_523; // @[Switch.scala 33:19:@2730.4]
  wire [47:0] _GEN_524; // @[Switch.scala 33:19:@2730.4]
  wire [47:0] _GEN_525; // @[Switch.scala 33:19:@2730.4]
  wire [47:0] _GEN_526; // @[Switch.scala 33:19:@2730.4]
  wire [47:0] _GEN_527; // @[Switch.scala 33:19:@2730.4]
  wire [47:0] _GEN_528; // @[Switch.scala 33:19:@2730.4]
  wire [47:0] _GEN_529; // @[Switch.scala 33:19:@2730.4]
  wire [47:0] _GEN_530; // @[Switch.scala 33:19:@2730.4]
  wire [47:0] _GEN_531; // @[Switch.scala 33:19:@2730.4]
  wire [47:0] _GEN_532; // @[Switch.scala 33:19:@2730.4]
  wire [47:0] _GEN_533; // @[Switch.scala 33:19:@2730.4]
  wire [47:0] _GEN_534; // @[Switch.scala 33:19:@2730.4]
  wire [47:0] _GEN_535; // @[Switch.scala 33:19:@2730.4]
  wire [47:0] _GEN_536; // @[Switch.scala 33:19:@2730.4]
  wire [47:0] _GEN_537; // @[Switch.scala 33:19:@2730.4]
  wire [47:0] _GEN_538; // @[Switch.scala 33:19:@2730.4]
  wire [47:0] _GEN_539; // @[Switch.scala 33:19:@2730.4]
  wire [47:0] _GEN_540; // @[Switch.scala 33:19:@2730.4]
  wire [47:0] _GEN_541; // @[Switch.scala 33:19:@2730.4]
  wire [47:0] _GEN_542; // @[Switch.scala 33:19:@2730.4]
  wire [7:0] _T_8011; // @[Switch.scala 34:32:@2737.4]
  wire [15:0] _T_8019; // @[Switch.scala 34:32:@2745.4]
  wire [7:0] _T_8026; // @[Switch.scala 34:32:@2752.4]
  wire [31:0] _T_8035; // @[Switch.scala 34:32:@2761.4]
  wire  _T_8039; // @[Switch.scala 30:53:@2764.4]
  wire  valid_17_0; // @[Switch.scala 30:36:@2765.4]
  wire  _T_8042; // @[Switch.scala 30:53:@2767.4]
  wire  valid_17_1; // @[Switch.scala 30:36:@2768.4]
  wire  _T_8045; // @[Switch.scala 30:53:@2770.4]
  wire  valid_17_2; // @[Switch.scala 30:36:@2771.4]
  wire  _T_8048; // @[Switch.scala 30:53:@2773.4]
  wire  valid_17_3; // @[Switch.scala 30:36:@2774.4]
  wire  _T_8051; // @[Switch.scala 30:53:@2776.4]
  wire  valid_17_4; // @[Switch.scala 30:36:@2777.4]
  wire  _T_8054; // @[Switch.scala 30:53:@2779.4]
  wire  valid_17_5; // @[Switch.scala 30:36:@2780.4]
  wire  _T_8057; // @[Switch.scala 30:53:@2782.4]
  wire  valid_17_6; // @[Switch.scala 30:36:@2783.4]
  wire  _T_8060; // @[Switch.scala 30:53:@2785.4]
  wire  valid_17_7; // @[Switch.scala 30:36:@2786.4]
  wire  _T_8063; // @[Switch.scala 30:53:@2788.4]
  wire  valid_17_8; // @[Switch.scala 30:36:@2789.4]
  wire  _T_8066; // @[Switch.scala 30:53:@2791.4]
  wire  valid_17_9; // @[Switch.scala 30:36:@2792.4]
  wire  _T_8069; // @[Switch.scala 30:53:@2794.4]
  wire  valid_17_10; // @[Switch.scala 30:36:@2795.4]
  wire  _T_8072; // @[Switch.scala 30:53:@2797.4]
  wire  valid_17_11; // @[Switch.scala 30:36:@2798.4]
  wire  _T_8075; // @[Switch.scala 30:53:@2800.4]
  wire  valid_17_12; // @[Switch.scala 30:36:@2801.4]
  wire  _T_8078; // @[Switch.scala 30:53:@2803.4]
  wire  valid_17_13; // @[Switch.scala 30:36:@2804.4]
  wire  _T_8081; // @[Switch.scala 30:53:@2806.4]
  wire  valid_17_14; // @[Switch.scala 30:36:@2807.4]
  wire  _T_8084; // @[Switch.scala 30:53:@2809.4]
  wire  valid_17_15; // @[Switch.scala 30:36:@2810.4]
  wire  _T_8087; // @[Switch.scala 30:53:@2812.4]
  wire  valid_17_16; // @[Switch.scala 30:36:@2813.4]
  wire  _T_8090; // @[Switch.scala 30:53:@2815.4]
  wire  valid_17_17; // @[Switch.scala 30:36:@2816.4]
  wire  _T_8093; // @[Switch.scala 30:53:@2818.4]
  wire  valid_17_18; // @[Switch.scala 30:36:@2819.4]
  wire  _T_8096; // @[Switch.scala 30:53:@2821.4]
  wire  valid_17_19; // @[Switch.scala 30:36:@2822.4]
  wire  _T_8099; // @[Switch.scala 30:53:@2824.4]
  wire  valid_17_20; // @[Switch.scala 30:36:@2825.4]
  wire  _T_8102; // @[Switch.scala 30:53:@2827.4]
  wire  valid_17_21; // @[Switch.scala 30:36:@2828.4]
  wire  _T_8105; // @[Switch.scala 30:53:@2830.4]
  wire  valid_17_22; // @[Switch.scala 30:36:@2831.4]
  wire  _T_8108; // @[Switch.scala 30:53:@2833.4]
  wire  valid_17_23; // @[Switch.scala 30:36:@2834.4]
  wire  _T_8111; // @[Switch.scala 30:53:@2836.4]
  wire  valid_17_24; // @[Switch.scala 30:36:@2837.4]
  wire  _T_8114; // @[Switch.scala 30:53:@2839.4]
  wire  valid_17_25; // @[Switch.scala 30:36:@2840.4]
  wire  _T_8117; // @[Switch.scala 30:53:@2842.4]
  wire  valid_17_26; // @[Switch.scala 30:36:@2843.4]
  wire  _T_8120; // @[Switch.scala 30:53:@2845.4]
  wire  valid_17_27; // @[Switch.scala 30:36:@2846.4]
  wire  _T_8123; // @[Switch.scala 30:53:@2848.4]
  wire  valid_17_28; // @[Switch.scala 30:36:@2849.4]
  wire  _T_8126; // @[Switch.scala 30:53:@2851.4]
  wire  valid_17_29; // @[Switch.scala 30:36:@2852.4]
  wire  _T_8129; // @[Switch.scala 30:53:@2854.4]
  wire  valid_17_30; // @[Switch.scala 30:36:@2855.4]
  wire  _T_8132; // @[Switch.scala 30:53:@2857.4]
  wire  valid_17_31; // @[Switch.scala 30:36:@2858.4]
  wire [4:0] _T_8166; // @[Mux.scala 31:69:@2860.4]
  wire [4:0] _T_8167; // @[Mux.scala 31:69:@2861.4]
  wire [4:0] _T_8168; // @[Mux.scala 31:69:@2862.4]
  wire [4:0] _T_8169; // @[Mux.scala 31:69:@2863.4]
  wire [4:0] _T_8170; // @[Mux.scala 31:69:@2864.4]
  wire [4:0] _T_8171; // @[Mux.scala 31:69:@2865.4]
  wire [4:0] _T_8172; // @[Mux.scala 31:69:@2866.4]
  wire [4:0] _T_8173; // @[Mux.scala 31:69:@2867.4]
  wire [4:0] _T_8174; // @[Mux.scala 31:69:@2868.4]
  wire [4:0] _T_8175; // @[Mux.scala 31:69:@2869.4]
  wire [4:0] _T_8176; // @[Mux.scala 31:69:@2870.4]
  wire [4:0] _T_8177; // @[Mux.scala 31:69:@2871.4]
  wire [4:0] _T_8178; // @[Mux.scala 31:69:@2872.4]
  wire [4:0] _T_8179; // @[Mux.scala 31:69:@2873.4]
  wire [4:0] _T_8180; // @[Mux.scala 31:69:@2874.4]
  wire [4:0] _T_8181; // @[Mux.scala 31:69:@2875.4]
  wire [4:0] _T_8182; // @[Mux.scala 31:69:@2876.4]
  wire [4:0] _T_8183; // @[Mux.scala 31:69:@2877.4]
  wire [4:0] _T_8184; // @[Mux.scala 31:69:@2878.4]
  wire [4:0] _T_8185; // @[Mux.scala 31:69:@2879.4]
  wire [4:0] _T_8186; // @[Mux.scala 31:69:@2880.4]
  wire [4:0] _T_8187; // @[Mux.scala 31:69:@2881.4]
  wire [4:0] _T_8188; // @[Mux.scala 31:69:@2882.4]
  wire [4:0] _T_8189; // @[Mux.scala 31:69:@2883.4]
  wire [4:0] _T_8190; // @[Mux.scala 31:69:@2884.4]
  wire [4:0] _T_8191; // @[Mux.scala 31:69:@2885.4]
  wire [4:0] _T_8192; // @[Mux.scala 31:69:@2886.4]
  wire [4:0] _T_8193; // @[Mux.scala 31:69:@2887.4]
  wire [4:0] _T_8194; // @[Mux.scala 31:69:@2888.4]
  wire [4:0] _T_8195; // @[Mux.scala 31:69:@2889.4]
  wire [4:0] select_17; // @[Mux.scala 31:69:@2890.4]
  wire [47:0] _GEN_545; // @[Switch.scala 33:19:@2892.4]
  wire [47:0] _GEN_546; // @[Switch.scala 33:19:@2892.4]
  wire [47:0] _GEN_547; // @[Switch.scala 33:19:@2892.4]
  wire [47:0] _GEN_548; // @[Switch.scala 33:19:@2892.4]
  wire [47:0] _GEN_549; // @[Switch.scala 33:19:@2892.4]
  wire [47:0] _GEN_550; // @[Switch.scala 33:19:@2892.4]
  wire [47:0] _GEN_551; // @[Switch.scala 33:19:@2892.4]
  wire [47:0] _GEN_552; // @[Switch.scala 33:19:@2892.4]
  wire [47:0] _GEN_553; // @[Switch.scala 33:19:@2892.4]
  wire [47:0] _GEN_554; // @[Switch.scala 33:19:@2892.4]
  wire [47:0] _GEN_555; // @[Switch.scala 33:19:@2892.4]
  wire [47:0] _GEN_556; // @[Switch.scala 33:19:@2892.4]
  wire [47:0] _GEN_557; // @[Switch.scala 33:19:@2892.4]
  wire [47:0] _GEN_558; // @[Switch.scala 33:19:@2892.4]
  wire [47:0] _GEN_559; // @[Switch.scala 33:19:@2892.4]
  wire [47:0] _GEN_560; // @[Switch.scala 33:19:@2892.4]
  wire [47:0] _GEN_561; // @[Switch.scala 33:19:@2892.4]
  wire [47:0] _GEN_562; // @[Switch.scala 33:19:@2892.4]
  wire [47:0] _GEN_563; // @[Switch.scala 33:19:@2892.4]
  wire [47:0] _GEN_564; // @[Switch.scala 33:19:@2892.4]
  wire [47:0] _GEN_565; // @[Switch.scala 33:19:@2892.4]
  wire [47:0] _GEN_566; // @[Switch.scala 33:19:@2892.4]
  wire [47:0] _GEN_567; // @[Switch.scala 33:19:@2892.4]
  wire [47:0] _GEN_568; // @[Switch.scala 33:19:@2892.4]
  wire [47:0] _GEN_569; // @[Switch.scala 33:19:@2892.4]
  wire [47:0] _GEN_570; // @[Switch.scala 33:19:@2892.4]
  wire [47:0] _GEN_571; // @[Switch.scala 33:19:@2892.4]
  wire [47:0] _GEN_572; // @[Switch.scala 33:19:@2892.4]
  wire [47:0] _GEN_573; // @[Switch.scala 33:19:@2892.4]
  wire [47:0] _GEN_574; // @[Switch.scala 33:19:@2892.4]
  wire [7:0] _T_8204; // @[Switch.scala 34:32:@2899.4]
  wire [15:0] _T_8212; // @[Switch.scala 34:32:@2907.4]
  wire [7:0] _T_8219; // @[Switch.scala 34:32:@2914.4]
  wire [31:0] _T_8228; // @[Switch.scala 34:32:@2923.4]
  wire  _T_8232; // @[Switch.scala 30:53:@2926.4]
  wire  valid_18_0; // @[Switch.scala 30:36:@2927.4]
  wire  _T_8235; // @[Switch.scala 30:53:@2929.4]
  wire  valid_18_1; // @[Switch.scala 30:36:@2930.4]
  wire  _T_8238; // @[Switch.scala 30:53:@2932.4]
  wire  valid_18_2; // @[Switch.scala 30:36:@2933.4]
  wire  _T_8241; // @[Switch.scala 30:53:@2935.4]
  wire  valid_18_3; // @[Switch.scala 30:36:@2936.4]
  wire  _T_8244; // @[Switch.scala 30:53:@2938.4]
  wire  valid_18_4; // @[Switch.scala 30:36:@2939.4]
  wire  _T_8247; // @[Switch.scala 30:53:@2941.4]
  wire  valid_18_5; // @[Switch.scala 30:36:@2942.4]
  wire  _T_8250; // @[Switch.scala 30:53:@2944.4]
  wire  valid_18_6; // @[Switch.scala 30:36:@2945.4]
  wire  _T_8253; // @[Switch.scala 30:53:@2947.4]
  wire  valid_18_7; // @[Switch.scala 30:36:@2948.4]
  wire  _T_8256; // @[Switch.scala 30:53:@2950.4]
  wire  valid_18_8; // @[Switch.scala 30:36:@2951.4]
  wire  _T_8259; // @[Switch.scala 30:53:@2953.4]
  wire  valid_18_9; // @[Switch.scala 30:36:@2954.4]
  wire  _T_8262; // @[Switch.scala 30:53:@2956.4]
  wire  valid_18_10; // @[Switch.scala 30:36:@2957.4]
  wire  _T_8265; // @[Switch.scala 30:53:@2959.4]
  wire  valid_18_11; // @[Switch.scala 30:36:@2960.4]
  wire  _T_8268; // @[Switch.scala 30:53:@2962.4]
  wire  valid_18_12; // @[Switch.scala 30:36:@2963.4]
  wire  _T_8271; // @[Switch.scala 30:53:@2965.4]
  wire  valid_18_13; // @[Switch.scala 30:36:@2966.4]
  wire  _T_8274; // @[Switch.scala 30:53:@2968.4]
  wire  valid_18_14; // @[Switch.scala 30:36:@2969.4]
  wire  _T_8277; // @[Switch.scala 30:53:@2971.4]
  wire  valid_18_15; // @[Switch.scala 30:36:@2972.4]
  wire  _T_8280; // @[Switch.scala 30:53:@2974.4]
  wire  valid_18_16; // @[Switch.scala 30:36:@2975.4]
  wire  _T_8283; // @[Switch.scala 30:53:@2977.4]
  wire  valid_18_17; // @[Switch.scala 30:36:@2978.4]
  wire  _T_8286; // @[Switch.scala 30:53:@2980.4]
  wire  valid_18_18; // @[Switch.scala 30:36:@2981.4]
  wire  _T_8289; // @[Switch.scala 30:53:@2983.4]
  wire  valid_18_19; // @[Switch.scala 30:36:@2984.4]
  wire  _T_8292; // @[Switch.scala 30:53:@2986.4]
  wire  valid_18_20; // @[Switch.scala 30:36:@2987.4]
  wire  _T_8295; // @[Switch.scala 30:53:@2989.4]
  wire  valid_18_21; // @[Switch.scala 30:36:@2990.4]
  wire  _T_8298; // @[Switch.scala 30:53:@2992.4]
  wire  valid_18_22; // @[Switch.scala 30:36:@2993.4]
  wire  _T_8301; // @[Switch.scala 30:53:@2995.4]
  wire  valid_18_23; // @[Switch.scala 30:36:@2996.4]
  wire  _T_8304; // @[Switch.scala 30:53:@2998.4]
  wire  valid_18_24; // @[Switch.scala 30:36:@2999.4]
  wire  _T_8307; // @[Switch.scala 30:53:@3001.4]
  wire  valid_18_25; // @[Switch.scala 30:36:@3002.4]
  wire  _T_8310; // @[Switch.scala 30:53:@3004.4]
  wire  valid_18_26; // @[Switch.scala 30:36:@3005.4]
  wire  _T_8313; // @[Switch.scala 30:53:@3007.4]
  wire  valid_18_27; // @[Switch.scala 30:36:@3008.4]
  wire  _T_8316; // @[Switch.scala 30:53:@3010.4]
  wire  valid_18_28; // @[Switch.scala 30:36:@3011.4]
  wire  _T_8319; // @[Switch.scala 30:53:@3013.4]
  wire  valid_18_29; // @[Switch.scala 30:36:@3014.4]
  wire  _T_8322; // @[Switch.scala 30:53:@3016.4]
  wire  valid_18_30; // @[Switch.scala 30:36:@3017.4]
  wire  _T_8325; // @[Switch.scala 30:53:@3019.4]
  wire  valid_18_31; // @[Switch.scala 30:36:@3020.4]
  wire [4:0] _T_8359; // @[Mux.scala 31:69:@3022.4]
  wire [4:0] _T_8360; // @[Mux.scala 31:69:@3023.4]
  wire [4:0] _T_8361; // @[Mux.scala 31:69:@3024.4]
  wire [4:0] _T_8362; // @[Mux.scala 31:69:@3025.4]
  wire [4:0] _T_8363; // @[Mux.scala 31:69:@3026.4]
  wire [4:0] _T_8364; // @[Mux.scala 31:69:@3027.4]
  wire [4:0] _T_8365; // @[Mux.scala 31:69:@3028.4]
  wire [4:0] _T_8366; // @[Mux.scala 31:69:@3029.4]
  wire [4:0] _T_8367; // @[Mux.scala 31:69:@3030.4]
  wire [4:0] _T_8368; // @[Mux.scala 31:69:@3031.4]
  wire [4:0] _T_8369; // @[Mux.scala 31:69:@3032.4]
  wire [4:0] _T_8370; // @[Mux.scala 31:69:@3033.4]
  wire [4:0] _T_8371; // @[Mux.scala 31:69:@3034.4]
  wire [4:0] _T_8372; // @[Mux.scala 31:69:@3035.4]
  wire [4:0] _T_8373; // @[Mux.scala 31:69:@3036.4]
  wire [4:0] _T_8374; // @[Mux.scala 31:69:@3037.4]
  wire [4:0] _T_8375; // @[Mux.scala 31:69:@3038.4]
  wire [4:0] _T_8376; // @[Mux.scala 31:69:@3039.4]
  wire [4:0] _T_8377; // @[Mux.scala 31:69:@3040.4]
  wire [4:0] _T_8378; // @[Mux.scala 31:69:@3041.4]
  wire [4:0] _T_8379; // @[Mux.scala 31:69:@3042.4]
  wire [4:0] _T_8380; // @[Mux.scala 31:69:@3043.4]
  wire [4:0] _T_8381; // @[Mux.scala 31:69:@3044.4]
  wire [4:0] _T_8382; // @[Mux.scala 31:69:@3045.4]
  wire [4:0] _T_8383; // @[Mux.scala 31:69:@3046.4]
  wire [4:0] _T_8384; // @[Mux.scala 31:69:@3047.4]
  wire [4:0] _T_8385; // @[Mux.scala 31:69:@3048.4]
  wire [4:0] _T_8386; // @[Mux.scala 31:69:@3049.4]
  wire [4:0] _T_8387; // @[Mux.scala 31:69:@3050.4]
  wire [4:0] _T_8388; // @[Mux.scala 31:69:@3051.4]
  wire [4:0] select_18; // @[Mux.scala 31:69:@3052.4]
  wire [47:0] _GEN_577; // @[Switch.scala 33:19:@3054.4]
  wire [47:0] _GEN_578; // @[Switch.scala 33:19:@3054.4]
  wire [47:0] _GEN_579; // @[Switch.scala 33:19:@3054.4]
  wire [47:0] _GEN_580; // @[Switch.scala 33:19:@3054.4]
  wire [47:0] _GEN_581; // @[Switch.scala 33:19:@3054.4]
  wire [47:0] _GEN_582; // @[Switch.scala 33:19:@3054.4]
  wire [47:0] _GEN_583; // @[Switch.scala 33:19:@3054.4]
  wire [47:0] _GEN_584; // @[Switch.scala 33:19:@3054.4]
  wire [47:0] _GEN_585; // @[Switch.scala 33:19:@3054.4]
  wire [47:0] _GEN_586; // @[Switch.scala 33:19:@3054.4]
  wire [47:0] _GEN_587; // @[Switch.scala 33:19:@3054.4]
  wire [47:0] _GEN_588; // @[Switch.scala 33:19:@3054.4]
  wire [47:0] _GEN_589; // @[Switch.scala 33:19:@3054.4]
  wire [47:0] _GEN_590; // @[Switch.scala 33:19:@3054.4]
  wire [47:0] _GEN_591; // @[Switch.scala 33:19:@3054.4]
  wire [47:0] _GEN_592; // @[Switch.scala 33:19:@3054.4]
  wire [47:0] _GEN_593; // @[Switch.scala 33:19:@3054.4]
  wire [47:0] _GEN_594; // @[Switch.scala 33:19:@3054.4]
  wire [47:0] _GEN_595; // @[Switch.scala 33:19:@3054.4]
  wire [47:0] _GEN_596; // @[Switch.scala 33:19:@3054.4]
  wire [47:0] _GEN_597; // @[Switch.scala 33:19:@3054.4]
  wire [47:0] _GEN_598; // @[Switch.scala 33:19:@3054.4]
  wire [47:0] _GEN_599; // @[Switch.scala 33:19:@3054.4]
  wire [47:0] _GEN_600; // @[Switch.scala 33:19:@3054.4]
  wire [47:0] _GEN_601; // @[Switch.scala 33:19:@3054.4]
  wire [47:0] _GEN_602; // @[Switch.scala 33:19:@3054.4]
  wire [47:0] _GEN_603; // @[Switch.scala 33:19:@3054.4]
  wire [47:0] _GEN_604; // @[Switch.scala 33:19:@3054.4]
  wire [47:0] _GEN_605; // @[Switch.scala 33:19:@3054.4]
  wire [47:0] _GEN_606; // @[Switch.scala 33:19:@3054.4]
  wire [7:0] _T_8397; // @[Switch.scala 34:32:@3061.4]
  wire [15:0] _T_8405; // @[Switch.scala 34:32:@3069.4]
  wire [7:0] _T_8412; // @[Switch.scala 34:32:@3076.4]
  wire [31:0] _T_8421; // @[Switch.scala 34:32:@3085.4]
  wire  _T_8425; // @[Switch.scala 30:53:@3088.4]
  wire  valid_19_0; // @[Switch.scala 30:36:@3089.4]
  wire  _T_8428; // @[Switch.scala 30:53:@3091.4]
  wire  valid_19_1; // @[Switch.scala 30:36:@3092.4]
  wire  _T_8431; // @[Switch.scala 30:53:@3094.4]
  wire  valid_19_2; // @[Switch.scala 30:36:@3095.4]
  wire  _T_8434; // @[Switch.scala 30:53:@3097.4]
  wire  valid_19_3; // @[Switch.scala 30:36:@3098.4]
  wire  _T_8437; // @[Switch.scala 30:53:@3100.4]
  wire  valid_19_4; // @[Switch.scala 30:36:@3101.4]
  wire  _T_8440; // @[Switch.scala 30:53:@3103.4]
  wire  valid_19_5; // @[Switch.scala 30:36:@3104.4]
  wire  _T_8443; // @[Switch.scala 30:53:@3106.4]
  wire  valid_19_6; // @[Switch.scala 30:36:@3107.4]
  wire  _T_8446; // @[Switch.scala 30:53:@3109.4]
  wire  valid_19_7; // @[Switch.scala 30:36:@3110.4]
  wire  _T_8449; // @[Switch.scala 30:53:@3112.4]
  wire  valid_19_8; // @[Switch.scala 30:36:@3113.4]
  wire  _T_8452; // @[Switch.scala 30:53:@3115.4]
  wire  valid_19_9; // @[Switch.scala 30:36:@3116.4]
  wire  _T_8455; // @[Switch.scala 30:53:@3118.4]
  wire  valid_19_10; // @[Switch.scala 30:36:@3119.4]
  wire  _T_8458; // @[Switch.scala 30:53:@3121.4]
  wire  valid_19_11; // @[Switch.scala 30:36:@3122.4]
  wire  _T_8461; // @[Switch.scala 30:53:@3124.4]
  wire  valid_19_12; // @[Switch.scala 30:36:@3125.4]
  wire  _T_8464; // @[Switch.scala 30:53:@3127.4]
  wire  valid_19_13; // @[Switch.scala 30:36:@3128.4]
  wire  _T_8467; // @[Switch.scala 30:53:@3130.4]
  wire  valid_19_14; // @[Switch.scala 30:36:@3131.4]
  wire  _T_8470; // @[Switch.scala 30:53:@3133.4]
  wire  valid_19_15; // @[Switch.scala 30:36:@3134.4]
  wire  _T_8473; // @[Switch.scala 30:53:@3136.4]
  wire  valid_19_16; // @[Switch.scala 30:36:@3137.4]
  wire  _T_8476; // @[Switch.scala 30:53:@3139.4]
  wire  valid_19_17; // @[Switch.scala 30:36:@3140.4]
  wire  _T_8479; // @[Switch.scala 30:53:@3142.4]
  wire  valid_19_18; // @[Switch.scala 30:36:@3143.4]
  wire  _T_8482; // @[Switch.scala 30:53:@3145.4]
  wire  valid_19_19; // @[Switch.scala 30:36:@3146.4]
  wire  _T_8485; // @[Switch.scala 30:53:@3148.4]
  wire  valid_19_20; // @[Switch.scala 30:36:@3149.4]
  wire  _T_8488; // @[Switch.scala 30:53:@3151.4]
  wire  valid_19_21; // @[Switch.scala 30:36:@3152.4]
  wire  _T_8491; // @[Switch.scala 30:53:@3154.4]
  wire  valid_19_22; // @[Switch.scala 30:36:@3155.4]
  wire  _T_8494; // @[Switch.scala 30:53:@3157.4]
  wire  valid_19_23; // @[Switch.scala 30:36:@3158.4]
  wire  _T_8497; // @[Switch.scala 30:53:@3160.4]
  wire  valid_19_24; // @[Switch.scala 30:36:@3161.4]
  wire  _T_8500; // @[Switch.scala 30:53:@3163.4]
  wire  valid_19_25; // @[Switch.scala 30:36:@3164.4]
  wire  _T_8503; // @[Switch.scala 30:53:@3166.4]
  wire  valid_19_26; // @[Switch.scala 30:36:@3167.4]
  wire  _T_8506; // @[Switch.scala 30:53:@3169.4]
  wire  valid_19_27; // @[Switch.scala 30:36:@3170.4]
  wire  _T_8509; // @[Switch.scala 30:53:@3172.4]
  wire  valid_19_28; // @[Switch.scala 30:36:@3173.4]
  wire  _T_8512; // @[Switch.scala 30:53:@3175.4]
  wire  valid_19_29; // @[Switch.scala 30:36:@3176.4]
  wire  _T_8515; // @[Switch.scala 30:53:@3178.4]
  wire  valid_19_30; // @[Switch.scala 30:36:@3179.4]
  wire  _T_8518; // @[Switch.scala 30:53:@3181.4]
  wire  valid_19_31; // @[Switch.scala 30:36:@3182.4]
  wire [4:0] _T_8552; // @[Mux.scala 31:69:@3184.4]
  wire [4:0] _T_8553; // @[Mux.scala 31:69:@3185.4]
  wire [4:0] _T_8554; // @[Mux.scala 31:69:@3186.4]
  wire [4:0] _T_8555; // @[Mux.scala 31:69:@3187.4]
  wire [4:0] _T_8556; // @[Mux.scala 31:69:@3188.4]
  wire [4:0] _T_8557; // @[Mux.scala 31:69:@3189.4]
  wire [4:0] _T_8558; // @[Mux.scala 31:69:@3190.4]
  wire [4:0] _T_8559; // @[Mux.scala 31:69:@3191.4]
  wire [4:0] _T_8560; // @[Mux.scala 31:69:@3192.4]
  wire [4:0] _T_8561; // @[Mux.scala 31:69:@3193.4]
  wire [4:0] _T_8562; // @[Mux.scala 31:69:@3194.4]
  wire [4:0] _T_8563; // @[Mux.scala 31:69:@3195.4]
  wire [4:0] _T_8564; // @[Mux.scala 31:69:@3196.4]
  wire [4:0] _T_8565; // @[Mux.scala 31:69:@3197.4]
  wire [4:0] _T_8566; // @[Mux.scala 31:69:@3198.4]
  wire [4:0] _T_8567; // @[Mux.scala 31:69:@3199.4]
  wire [4:0] _T_8568; // @[Mux.scala 31:69:@3200.4]
  wire [4:0] _T_8569; // @[Mux.scala 31:69:@3201.4]
  wire [4:0] _T_8570; // @[Mux.scala 31:69:@3202.4]
  wire [4:0] _T_8571; // @[Mux.scala 31:69:@3203.4]
  wire [4:0] _T_8572; // @[Mux.scala 31:69:@3204.4]
  wire [4:0] _T_8573; // @[Mux.scala 31:69:@3205.4]
  wire [4:0] _T_8574; // @[Mux.scala 31:69:@3206.4]
  wire [4:0] _T_8575; // @[Mux.scala 31:69:@3207.4]
  wire [4:0] _T_8576; // @[Mux.scala 31:69:@3208.4]
  wire [4:0] _T_8577; // @[Mux.scala 31:69:@3209.4]
  wire [4:0] _T_8578; // @[Mux.scala 31:69:@3210.4]
  wire [4:0] _T_8579; // @[Mux.scala 31:69:@3211.4]
  wire [4:0] _T_8580; // @[Mux.scala 31:69:@3212.4]
  wire [4:0] _T_8581; // @[Mux.scala 31:69:@3213.4]
  wire [4:0] select_19; // @[Mux.scala 31:69:@3214.4]
  wire [47:0] _GEN_609; // @[Switch.scala 33:19:@3216.4]
  wire [47:0] _GEN_610; // @[Switch.scala 33:19:@3216.4]
  wire [47:0] _GEN_611; // @[Switch.scala 33:19:@3216.4]
  wire [47:0] _GEN_612; // @[Switch.scala 33:19:@3216.4]
  wire [47:0] _GEN_613; // @[Switch.scala 33:19:@3216.4]
  wire [47:0] _GEN_614; // @[Switch.scala 33:19:@3216.4]
  wire [47:0] _GEN_615; // @[Switch.scala 33:19:@3216.4]
  wire [47:0] _GEN_616; // @[Switch.scala 33:19:@3216.4]
  wire [47:0] _GEN_617; // @[Switch.scala 33:19:@3216.4]
  wire [47:0] _GEN_618; // @[Switch.scala 33:19:@3216.4]
  wire [47:0] _GEN_619; // @[Switch.scala 33:19:@3216.4]
  wire [47:0] _GEN_620; // @[Switch.scala 33:19:@3216.4]
  wire [47:0] _GEN_621; // @[Switch.scala 33:19:@3216.4]
  wire [47:0] _GEN_622; // @[Switch.scala 33:19:@3216.4]
  wire [47:0] _GEN_623; // @[Switch.scala 33:19:@3216.4]
  wire [47:0] _GEN_624; // @[Switch.scala 33:19:@3216.4]
  wire [47:0] _GEN_625; // @[Switch.scala 33:19:@3216.4]
  wire [47:0] _GEN_626; // @[Switch.scala 33:19:@3216.4]
  wire [47:0] _GEN_627; // @[Switch.scala 33:19:@3216.4]
  wire [47:0] _GEN_628; // @[Switch.scala 33:19:@3216.4]
  wire [47:0] _GEN_629; // @[Switch.scala 33:19:@3216.4]
  wire [47:0] _GEN_630; // @[Switch.scala 33:19:@3216.4]
  wire [47:0] _GEN_631; // @[Switch.scala 33:19:@3216.4]
  wire [47:0] _GEN_632; // @[Switch.scala 33:19:@3216.4]
  wire [47:0] _GEN_633; // @[Switch.scala 33:19:@3216.4]
  wire [47:0] _GEN_634; // @[Switch.scala 33:19:@3216.4]
  wire [47:0] _GEN_635; // @[Switch.scala 33:19:@3216.4]
  wire [47:0] _GEN_636; // @[Switch.scala 33:19:@3216.4]
  wire [47:0] _GEN_637; // @[Switch.scala 33:19:@3216.4]
  wire [47:0] _GEN_638; // @[Switch.scala 33:19:@3216.4]
  wire [7:0] _T_8590; // @[Switch.scala 34:32:@3223.4]
  wire [15:0] _T_8598; // @[Switch.scala 34:32:@3231.4]
  wire [7:0] _T_8605; // @[Switch.scala 34:32:@3238.4]
  wire [31:0] _T_8614; // @[Switch.scala 34:32:@3247.4]
  wire  _T_8618; // @[Switch.scala 30:53:@3250.4]
  wire  valid_20_0; // @[Switch.scala 30:36:@3251.4]
  wire  _T_8621; // @[Switch.scala 30:53:@3253.4]
  wire  valid_20_1; // @[Switch.scala 30:36:@3254.4]
  wire  _T_8624; // @[Switch.scala 30:53:@3256.4]
  wire  valid_20_2; // @[Switch.scala 30:36:@3257.4]
  wire  _T_8627; // @[Switch.scala 30:53:@3259.4]
  wire  valid_20_3; // @[Switch.scala 30:36:@3260.4]
  wire  _T_8630; // @[Switch.scala 30:53:@3262.4]
  wire  valid_20_4; // @[Switch.scala 30:36:@3263.4]
  wire  _T_8633; // @[Switch.scala 30:53:@3265.4]
  wire  valid_20_5; // @[Switch.scala 30:36:@3266.4]
  wire  _T_8636; // @[Switch.scala 30:53:@3268.4]
  wire  valid_20_6; // @[Switch.scala 30:36:@3269.4]
  wire  _T_8639; // @[Switch.scala 30:53:@3271.4]
  wire  valid_20_7; // @[Switch.scala 30:36:@3272.4]
  wire  _T_8642; // @[Switch.scala 30:53:@3274.4]
  wire  valid_20_8; // @[Switch.scala 30:36:@3275.4]
  wire  _T_8645; // @[Switch.scala 30:53:@3277.4]
  wire  valid_20_9; // @[Switch.scala 30:36:@3278.4]
  wire  _T_8648; // @[Switch.scala 30:53:@3280.4]
  wire  valid_20_10; // @[Switch.scala 30:36:@3281.4]
  wire  _T_8651; // @[Switch.scala 30:53:@3283.4]
  wire  valid_20_11; // @[Switch.scala 30:36:@3284.4]
  wire  _T_8654; // @[Switch.scala 30:53:@3286.4]
  wire  valid_20_12; // @[Switch.scala 30:36:@3287.4]
  wire  _T_8657; // @[Switch.scala 30:53:@3289.4]
  wire  valid_20_13; // @[Switch.scala 30:36:@3290.4]
  wire  _T_8660; // @[Switch.scala 30:53:@3292.4]
  wire  valid_20_14; // @[Switch.scala 30:36:@3293.4]
  wire  _T_8663; // @[Switch.scala 30:53:@3295.4]
  wire  valid_20_15; // @[Switch.scala 30:36:@3296.4]
  wire  _T_8666; // @[Switch.scala 30:53:@3298.4]
  wire  valid_20_16; // @[Switch.scala 30:36:@3299.4]
  wire  _T_8669; // @[Switch.scala 30:53:@3301.4]
  wire  valid_20_17; // @[Switch.scala 30:36:@3302.4]
  wire  _T_8672; // @[Switch.scala 30:53:@3304.4]
  wire  valid_20_18; // @[Switch.scala 30:36:@3305.4]
  wire  _T_8675; // @[Switch.scala 30:53:@3307.4]
  wire  valid_20_19; // @[Switch.scala 30:36:@3308.4]
  wire  _T_8678; // @[Switch.scala 30:53:@3310.4]
  wire  valid_20_20; // @[Switch.scala 30:36:@3311.4]
  wire  _T_8681; // @[Switch.scala 30:53:@3313.4]
  wire  valid_20_21; // @[Switch.scala 30:36:@3314.4]
  wire  _T_8684; // @[Switch.scala 30:53:@3316.4]
  wire  valid_20_22; // @[Switch.scala 30:36:@3317.4]
  wire  _T_8687; // @[Switch.scala 30:53:@3319.4]
  wire  valid_20_23; // @[Switch.scala 30:36:@3320.4]
  wire  _T_8690; // @[Switch.scala 30:53:@3322.4]
  wire  valid_20_24; // @[Switch.scala 30:36:@3323.4]
  wire  _T_8693; // @[Switch.scala 30:53:@3325.4]
  wire  valid_20_25; // @[Switch.scala 30:36:@3326.4]
  wire  _T_8696; // @[Switch.scala 30:53:@3328.4]
  wire  valid_20_26; // @[Switch.scala 30:36:@3329.4]
  wire  _T_8699; // @[Switch.scala 30:53:@3331.4]
  wire  valid_20_27; // @[Switch.scala 30:36:@3332.4]
  wire  _T_8702; // @[Switch.scala 30:53:@3334.4]
  wire  valid_20_28; // @[Switch.scala 30:36:@3335.4]
  wire  _T_8705; // @[Switch.scala 30:53:@3337.4]
  wire  valid_20_29; // @[Switch.scala 30:36:@3338.4]
  wire  _T_8708; // @[Switch.scala 30:53:@3340.4]
  wire  valid_20_30; // @[Switch.scala 30:36:@3341.4]
  wire  _T_8711; // @[Switch.scala 30:53:@3343.4]
  wire  valid_20_31; // @[Switch.scala 30:36:@3344.4]
  wire [4:0] _T_8745; // @[Mux.scala 31:69:@3346.4]
  wire [4:0] _T_8746; // @[Mux.scala 31:69:@3347.4]
  wire [4:0] _T_8747; // @[Mux.scala 31:69:@3348.4]
  wire [4:0] _T_8748; // @[Mux.scala 31:69:@3349.4]
  wire [4:0] _T_8749; // @[Mux.scala 31:69:@3350.4]
  wire [4:0] _T_8750; // @[Mux.scala 31:69:@3351.4]
  wire [4:0] _T_8751; // @[Mux.scala 31:69:@3352.4]
  wire [4:0] _T_8752; // @[Mux.scala 31:69:@3353.4]
  wire [4:0] _T_8753; // @[Mux.scala 31:69:@3354.4]
  wire [4:0] _T_8754; // @[Mux.scala 31:69:@3355.4]
  wire [4:0] _T_8755; // @[Mux.scala 31:69:@3356.4]
  wire [4:0] _T_8756; // @[Mux.scala 31:69:@3357.4]
  wire [4:0] _T_8757; // @[Mux.scala 31:69:@3358.4]
  wire [4:0] _T_8758; // @[Mux.scala 31:69:@3359.4]
  wire [4:0] _T_8759; // @[Mux.scala 31:69:@3360.4]
  wire [4:0] _T_8760; // @[Mux.scala 31:69:@3361.4]
  wire [4:0] _T_8761; // @[Mux.scala 31:69:@3362.4]
  wire [4:0] _T_8762; // @[Mux.scala 31:69:@3363.4]
  wire [4:0] _T_8763; // @[Mux.scala 31:69:@3364.4]
  wire [4:0] _T_8764; // @[Mux.scala 31:69:@3365.4]
  wire [4:0] _T_8765; // @[Mux.scala 31:69:@3366.4]
  wire [4:0] _T_8766; // @[Mux.scala 31:69:@3367.4]
  wire [4:0] _T_8767; // @[Mux.scala 31:69:@3368.4]
  wire [4:0] _T_8768; // @[Mux.scala 31:69:@3369.4]
  wire [4:0] _T_8769; // @[Mux.scala 31:69:@3370.4]
  wire [4:0] _T_8770; // @[Mux.scala 31:69:@3371.4]
  wire [4:0] _T_8771; // @[Mux.scala 31:69:@3372.4]
  wire [4:0] _T_8772; // @[Mux.scala 31:69:@3373.4]
  wire [4:0] _T_8773; // @[Mux.scala 31:69:@3374.4]
  wire [4:0] _T_8774; // @[Mux.scala 31:69:@3375.4]
  wire [4:0] select_20; // @[Mux.scala 31:69:@3376.4]
  wire [47:0] _GEN_641; // @[Switch.scala 33:19:@3378.4]
  wire [47:0] _GEN_642; // @[Switch.scala 33:19:@3378.4]
  wire [47:0] _GEN_643; // @[Switch.scala 33:19:@3378.4]
  wire [47:0] _GEN_644; // @[Switch.scala 33:19:@3378.4]
  wire [47:0] _GEN_645; // @[Switch.scala 33:19:@3378.4]
  wire [47:0] _GEN_646; // @[Switch.scala 33:19:@3378.4]
  wire [47:0] _GEN_647; // @[Switch.scala 33:19:@3378.4]
  wire [47:0] _GEN_648; // @[Switch.scala 33:19:@3378.4]
  wire [47:0] _GEN_649; // @[Switch.scala 33:19:@3378.4]
  wire [47:0] _GEN_650; // @[Switch.scala 33:19:@3378.4]
  wire [47:0] _GEN_651; // @[Switch.scala 33:19:@3378.4]
  wire [47:0] _GEN_652; // @[Switch.scala 33:19:@3378.4]
  wire [47:0] _GEN_653; // @[Switch.scala 33:19:@3378.4]
  wire [47:0] _GEN_654; // @[Switch.scala 33:19:@3378.4]
  wire [47:0] _GEN_655; // @[Switch.scala 33:19:@3378.4]
  wire [47:0] _GEN_656; // @[Switch.scala 33:19:@3378.4]
  wire [47:0] _GEN_657; // @[Switch.scala 33:19:@3378.4]
  wire [47:0] _GEN_658; // @[Switch.scala 33:19:@3378.4]
  wire [47:0] _GEN_659; // @[Switch.scala 33:19:@3378.4]
  wire [47:0] _GEN_660; // @[Switch.scala 33:19:@3378.4]
  wire [47:0] _GEN_661; // @[Switch.scala 33:19:@3378.4]
  wire [47:0] _GEN_662; // @[Switch.scala 33:19:@3378.4]
  wire [47:0] _GEN_663; // @[Switch.scala 33:19:@3378.4]
  wire [47:0] _GEN_664; // @[Switch.scala 33:19:@3378.4]
  wire [47:0] _GEN_665; // @[Switch.scala 33:19:@3378.4]
  wire [47:0] _GEN_666; // @[Switch.scala 33:19:@3378.4]
  wire [47:0] _GEN_667; // @[Switch.scala 33:19:@3378.4]
  wire [47:0] _GEN_668; // @[Switch.scala 33:19:@3378.4]
  wire [47:0] _GEN_669; // @[Switch.scala 33:19:@3378.4]
  wire [47:0] _GEN_670; // @[Switch.scala 33:19:@3378.4]
  wire [7:0] _T_8783; // @[Switch.scala 34:32:@3385.4]
  wire [15:0] _T_8791; // @[Switch.scala 34:32:@3393.4]
  wire [7:0] _T_8798; // @[Switch.scala 34:32:@3400.4]
  wire [31:0] _T_8807; // @[Switch.scala 34:32:@3409.4]
  wire  _T_8811; // @[Switch.scala 30:53:@3412.4]
  wire  valid_21_0; // @[Switch.scala 30:36:@3413.4]
  wire  _T_8814; // @[Switch.scala 30:53:@3415.4]
  wire  valid_21_1; // @[Switch.scala 30:36:@3416.4]
  wire  _T_8817; // @[Switch.scala 30:53:@3418.4]
  wire  valid_21_2; // @[Switch.scala 30:36:@3419.4]
  wire  _T_8820; // @[Switch.scala 30:53:@3421.4]
  wire  valid_21_3; // @[Switch.scala 30:36:@3422.4]
  wire  _T_8823; // @[Switch.scala 30:53:@3424.4]
  wire  valid_21_4; // @[Switch.scala 30:36:@3425.4]
  wire  _T_8826; // @[Switch.scala 30:53:@3427.4]
  wire  valid_21_5; // @[Switch.scala 30:36:@3428.4]
  wire  _T_8829; // @[Switch.scala 30:53:@3430.4]
  wire  valid_21_6; // @[Switch.scala 30:36:@3431.4]
  wire  _T_8832; // @[Switch.scala 30:53:@3433.4]
  wire  valid_21_7; // @[Switch.scala 30:36:@3434.4]
  wire  _T_8835; // @[Switch.scala 30:53:@3436.4]
  wire  valid_21_8; // @[Switch.scala 30:36:@3437.4]
  wire  _T_8838; // @[Switch.scala 30:53:@3439.4]
  wire  valid_21_9; // @[Switch.scala 30:36:@3440.4]
  wire  _T_8841; // @[Switch.scala 30:53:@3442.4]
  wire  valid_21_10; // @[Switch.scala 30:36:@3443.4]
  wire  _T_8844; // @[Switch.scala 30:53:@3445.4]
  wire  valid_21_11; // @[Switch.scala 30:36:@3446.4]
  wire  _T_8847; // @[Switch.scala 30:53:@3448.4]
  wire  valid_21_12; // @[Switch.scala 30:36:@3449.4]
  wire  _T_8850; // @[Switch.scala 30:53:@3451.4]
  wire  valid_21_13; // @[Switch.scala 30:36:@3452.4]
  wire  _T_8853; // @[Switch.scala 30:53:@3454.4]
  wire  valid_21_14; // @[Switch.scala 30:36:@3455.4]
  wire  _T_8856; // @[Switch.scala 30:53:@3457.4]
  wire  valid_21_15; // @[Switch.scala 30:36:@3458.4]
  wire  _T_8859; // @[Switch.scala 30:53:@3460.4]
  wire  valid_21_16; // @[Switch.scala 30:36:@3461.4]
  wire  _T_8862; // @[Switch.scala 30:53:@3463.4]
  wire  valid_21_17; // @[Switch.scala 30:36:@3464.4]
  wire  _T_8865; // @[Switch.scala 30:53:@3466.4]
  wire  valid_21_18; // @[Switch.scala 30:36:@3467.4]
  wire  _T_8868; // @[Switch.scala 30:53:@3469.4]
  wire  valid_21_19; // @[Switch.scala 30:36:@3470.4]
  wire  _T_8871; // @[Switch.scala 30:53:@3472.4]
  wire  valid_21_20; // @[Switch.scala 30:36:@3473.4]
  wire  _T_8874; // @[Switch.scala 30:53:@3475.4]
  wire  valid_21_21; // @[Switch.scala 30:36:@3476.4]
  wire  _T_8877; // @[Switch.scala 30:53:@3478.4]
  wire  valid_21_22; // @[Switch.scala 30:36:@3479.4]
  wire  _T_8880; // @[Switch.scala 30:53:@3481.4]
  wire  valid_21_23; // @[Switch.scala 30:36:@3482.4]
  wire  _T_8883; // @[Switch.scala 30:53:@3484.4]
  wire  valid_21_24; // @[Switch.scala 30:36:@3485.4]
  wire  _T_8886; // @[Switch.scala 30:53:@3487.4]
  wire  valid_21_25; // @[Switch.scala 30:36:@3488.4]
  wire  _T_8889; // @[Switch.scala 30:53:@3490.4]
  wire  valid_21_26; // @[Switch.scala 30:36:@3491.4]
  wire  _T_8892; // @[Switch.scala 30:53:@3493.4]
  wire  valid_21_27; // @[Switch.scala 30:36:@3494.4]
  wire  _T_8895; // @[Switch.scala 30:53:@3496.4]
  wire  valid_21_28; // @[Switch.scala 30:36:@3497.4]
  wire  _T_8898; // @[Switch.scala 30:53:@3499.4]
  wire  valid_21_29; // @[Switch.scala 30:36:@3500.4]
  wire  _T_8901; // @[Switch.scala 30:53:@3502.4]
  wire  valid_21_30; // @[Switch.scala 30:36:@3503.4]
  wire  _T_8904; // @[Switch.scala 30:53:@3505.4]
  wire  valid_21_31; // @[Switch.scala 30:36:@3506.4]
  wire [4:0] _T_8938; // @[Mux.scala 31:69:@3508.4]
  wire [4:0] _T_8939; // @[Mux.scala 31:69:@3509.4]
  wire [4:0] _T_8940; // @[Mux.scala 31:69:@3510.4]
  wire [4:0] _T_8941; // @[Mux.scala 31:69:@3511.4]
  wire [4:0] _T_8942; // @[Mux.scala 31:69:@3512.4]
  wire [4:0] _T_8943; // @[Mux.scala 31:69:@3513.4]
  wire [4:0] _T_8944; // @[Mux.scala 31:69:@3514.4]
  wire [4:0] _T_8945; // @[Mux.scala 31:69:@3515.4]
  wire [4:0] _T_8946; // @[Mux.scala 31:69:@3516.4]
  wire [4:0] _T_8947; // @[Mux.scala 31:69:@3517.4]
  wire [4:0] _T_8948; // @[Mux.scala 31:69:@3518.4]
  wire [4:0] _T_8949; // @[Mux.scala 31:69:@3519.4]
  wire [4:0] _T_8950; // @[Mux.scala 31:69:@3520.4]
  wire [4:0] _T_8951; // @[Mux.scala 31:69:@3521.4]
  wire [4:0] _T_8952; // @[Mux.scala 31:69:@3522.4]
  wire [4:0] _T_8953; // @[Mux.scala 31:69:@3523.4]
  wire [4:0] _T_8954; // @[Mux.scala 31:69:@3524.4]
  wire [4:0] _T_8955; // @[Mux.scala 31:69:@3525.4]
  wire [4:0] _T_8956; // @[Mux.scala 31:69:@3526.4]
  wire [4:0] _T_8957; // @[Mux.scala 31:69:@3527.4]
  wire [4:0] _T_8958; // @[Mux.scala 31:69:@3528.4]
  wire [4:0] _T_8959; // @[Mux.scala 31:69:@3529.4]
  wire [4:0] _T_8960; // @[Mux.scala 31:69:@3530.4]
  wire [4:0] _T_8961; // @[Mux.scala 31:69:@3531.4]
  wire [4:0] _T_8962; // @[Mux.scala 31:69:@3532.4]
  wire [4:0] _T_8963; // @[Mux.scala 31:69:@3533.4]
  wire [4:0] _T_8964; // @[Mux.scala 31:69:@3534.4]
  wire [4:0] _T_8965; // @[Mux.scala 31:69:@3535.4]
  wire [4:0] _T_8966; // @[Mux.scala 31:69:@3536.4]
  wire [4:0] _T_8967; // @[Mux.scala 31:69:@3537.4]
  wire [4:0] select_21; // @[Mux.scala 31:69:@3538.4]
  wire [47:0] _GEN_673; // @[Switch.scala 33:19:@3540.4]
  wire [47:0] _GEN_674; // @[Switch.scala 33:19:@3540.4]
  wire [47:0] _GEN_675; // @[Switch.scala 33:19:@3540.4]
  wire [47:0] _GEN_676; // @[Switch.scala 33:19:@3540.4]
  wire [47:0] _GEN_677; // @[Switch.scala 33:19:@3540.4]
  wire [47:0] _GEN_678; // @[Switch.scala 33:19:@3540.4]
  wire [47:0] _GEN_679; // @[Switch.scala 33:19:@3540.4]
  wire [47:0] _GEN_680; // @[Switch.scala 33:19:@3540.4]
  wire [47:0] _GEN_681; // @[Switch.scala 33:19:@3540.4]
  wire [47:0] _GEN_682; // @[Switch.scala 33:19:@3540.4]
  wire [47:0] _GEN_683; // @[Switch.scala 33:19:@3540.4]
  wire [47:0] _GEN_684; // @[Switch.scala 33:19:@3540.4]
  wire [47:0] _GEN_685; // @[Switch.scala 33:19:@3540.4]
  wire [47:0] _GEN_686; // @[Switch.scala 33:19:@3540.4]
  wire [47:0] _GEN_687; // @[Switch.scala 33:19:@3540.4]
  wire [47:0] _GEN_688; // @[Switch.scala 33:19:@3540.4]
  wire [47:0] _GEN_689; // @[Switch.scala 33:19:@3540.4]
  wire [47:0] _GEN_690; // @[Switch.scala 33:19:@3540.4]
  wire [47:0] _GEN_691; // @[Switch.scala 33:19:@3540.4]
  wire [47:0] _GEN_692; // @[Switch.scala 33:19:@3540.4]
  wire [47:0] _GEN_693; // @[Switch.scala 33:19:@3540.4]
  wire [47:0] _GEN_694; // @[Switch.scala 33:19:@3540.4]
  wire [47:0] _GEN_695; // @[Switch.scala 33:19:@3540.4]
  wire [47:0] _GEN_696; // @[Switch.scala 33:19:@3540.4]
  wire [47:0] _GEN_697; // @[Switch.scala 33:19:@3540.4]
  wire [47:0] _GEN_698; // @[Switch.scala 33:19:@3540.4]
  wire [47:0] _GEN_699; // @[Switch.scala 33:19:@3540.4]
  wire [47:0] _GEN_700; // @[Switch.scala 33:19:@3540.4]
  wire [47:0] _GEN_701; // @[Switch.scala 33:19:@3540.4]
  wire [47:0] _GEN_702; // @[Switch.scala 33:19:@3540.4]
  wire [7:0] _T_8976; // @[Switch.scala 34:32:@3547.4]
  wire [15:0] _T_8984; // @[Switch.scala 34:32:@3555.4]
  wire [7:0] _T_8991; // @[Switch.scala 34:32:@3562.4]
  wire [31:0] _T_9000; // @[Switch.scala 34:32:@3571.4]
  wire  _T_9004; // @[Switch.scala 30:53:@3574.4]
  wire  valid_22_0; // @[Switch.scala 30:36:@3575.4]
  wire  _T_9007; // @[Switch.scala 30:53:@3577.4]
  wire  valid_22_1; // @[Switch.scala 30:36:@3578.4]
  wire  _T_9010; // @[Switch.scala 30:53:@3580.4]
  wire  valid_22_2; // @[Switch.scala 30:36:@3581.4]
  wire  _T_9013; // @[Switch.scala 30:53:@3583.4]
  wire  valid_22_3; // @[Switch.scala 30:36:@3584.4]
  wire  _T_9016; // @[Switch.scala 30:53:@3586.4]
  wire  valid_22_4; // @[Switch.scala 30:36:@3587.4]
  wire  _T_9019; // @[Switch.scala 30:53:@3589.4]
  wire  valid_22_5; // @[Switch.scala 30:36:@3590.4]
  wire  _T_9022; // @[Switch.scala 30:53:@3592.4]
  wire  valid_22_6; // @[Switch.scala 30:36:@3593.4]
  wire  _T_9025; // @[Switch.scala 30:53:@3595.4]
  wire  valid_22_7; // @[Switch.scala 30:36:@3596.4]
  wire  _T_9028; // @[Switch.scala 30:53:@3598.4]
  wire  valid_22_8; // @[Switch.scala 30:36:@3599.4]
  wire  _T_9031; // @[Switch.scala 30:53:@3601.4]
  wire  valid_22_9; // @[Switch.scala 30:36:@3602.4]
  wire  _T_9034; // @[Switch.scala 30:53:@3604.4]
  wire  valid_22_10; // @[Switch.scala 30:36:@3605.4]
  wire  _T_9037; // @[Switch.scala 30:53:@3607.4]
  wire  valid_22_11; // @[Switch.scala 30:36:@3608.4]
  wire  _T_9040; // @[Switch.scala 30:53:@3610.4]
  wire  valid_22_12; // @[Switch.scala 30:36:@3611.4]
  wire  _T_9043; // @[Switch.scala 30:53:@3613.4]
  wire  valid_22_13; // @[Switch.scala 30:36:@3614.4]
  wire  _T_9046; // @[Switch.scala 30:53:@3616.4]
  wire  valid_22_14; // @[Switch.scala 30:36:@3617.4]
  wire  _T_9049; // @[Switch.scala 30:53:@3619.4]
  wire  valid_22_15; // @[Switch.scala 30:36:@3620.4]
  wire  _T_9052; // @[Switch.scala 30:53:@3622.4]
  wire  valid_22_16; // @[Switch.scala 30:36:@3623.4]
  wire  _T_9055; // @[Switch.scala 30:53:@3625.4]
  wire  valid_22_17; // @[Switch.scala 30:36:@3626.4]
  wire  _T_9058; // @[Switch.scala 30:53:@3628.4]
  wire  valid_22_18; // @[Switch.scala 30:36:@3629.4]
  wire  _T_9061; // @[Switch.scala 30:53:@3631.4]
  wire  valid_22_19; // @[Switch.scala 30:36:@3632.4]
  wire  _T_9064; // @[Switch.scala 30:53:@3634.4]
  wire  valid_22_20; // @[Switch.scala 30:36:@3635.4]
  wire  _T_9067; // @[Switch.scala 30:53:@3637.4]
  wire  valid_22_21; // @[Switch.scala 30:36:@3638.4]
  wire  _T_9070; // @[Switch.scala 30:53:@3640.4]
  wire  valid_22_22; // @[Switch.scala 30:36:@3641.4]
  wire  _T_9073; // @[Switch.scala 30:53:@3643.4]
  wire  valid_22_23; // @[Switch.scala 30:36:@3644.4]
  wire  _T_9076; // @[Switch.scala 30:53:@3646.4]
  wire  valid_22_24; // @[Switch.scala 30:36:@3647.4]
  wire  _T_9079; // @[Switch.scala 30:53:@3649.4]
  wire  valid_22_25; // @[Switch.scala 30:36:@3650.4]
  wire  _T_9082; // @[Switch.scala 30:53:@3652.4]
  wire  valid_22_26; // @[Switch.scala 30:36:@3653.4]
  wire  _T_9085; // @[Switch.scala 30:53:@3655.4]
  wire  valid_22_27; // @[Switch.scala 30:36:@3656.4]
  wire  _T_9088; // @[Switch.scala 30:53:@3658.4]
  wire  valid_22_28; // @[Switch.scala 30:36:@3659.4]
  wire  _T_9091; // @[Switch.scala 30:53:@3661.4]
  wire  valid_22_29; // @[Switch.scala 30:36:@3662.4]
  wire  _T_9094; // @[Switch.scala 30:53:@3664.4]
  wire  valid_22_30; // @[Switch.scala 30:36:@3665.4]
  wire  _T_9097; // @[Switch.scala 30:53:@3667.4]
  wire  valid_22_31; // @[Switch.scala 30:36:@3668.4]
  wire [4:0] _T_9131; // @[Mux.scala 31:69:@3670.4]
  wire [4:0] _T_9132; // @[Mux.scala 31:69:@3671.4]
  wire [4:0] _T_9133; // @[Mux.scala 31:69:@3672.4]
  wire [4:0] _T_9134; // @[Mux.scala 31:69:@3673.4]
  wire [4:0] _T_9135; // @[Mux.scala 31:69:@3674.4]
  wire [4:0] _T_9136; // @[Mux.scala 31:69:@3675.4]
  wire [4:0] _T_9137; // @[Mux.scala 31:69:@3676.4]
  wire [4:0] _T_9138; // @[Mux.scala 31:69:@3677.4]
  wire [4:0] _T_9139; // @[Mux.scala 31:69:@3678.4]
  wire [4:0] _T_9140; // @[Mux.scala 31:69:@3679.4]
  wire [4:0] _T_9141; // @[Mux.scala 31:69:@3680.4]
  wire [4:0] _T_9142; // @[Mux.scala 31:69:@3681.4]
  wire [4:0] _T_9143; // @[Mux.scala 31:69:@3682.4]
  wire [4:0] _T_9144; // @[Mux.scala 31:69:@3683.4]
  wire [4:0] _T_9145; // @[Mux.scala 31:69:@3684.4]
  wire [4:0] _T_9146; // @[Mux.scala 31:69:@3685.4]
  wire [4:0] _T_9147; // @[Mux.scala 31:69:@3686.4]
  wire [4:0] _T_9148; // @[Mux.scala 31:69:@3687.4]
  wire [4:0] _T_9149; // @[Mux.scala 31:69:@3688.4]
  wire [4:0] _T_9150; // @[Mux.scala 31:69:@3689.4]
  wire [4:0] _T_9151; // @[Mux.scala 31:69:@3690.4]
  wire [4:0] _T_9152; // @[Mux.scala 31:69:@3691.4]
  wire [4:0] _T_9153; // @[Mux.scala 31:69:@3692.4]
  wire [4:0] _T_9154; // @[Mux.scala 31:69:@3693.4]
  wire [4:0] _T_9155; // @[Mux.scala 31:69:@3694.4]
  wire [4:0] _T_9156; // @[Mux.scala 31:69:@3695.4]
  wire [4:0] _T_9157; // @[Mux.scala 31:69:@3696.4]
  wire [4:0] _T_9158; // @[Mux.scala 31:69:@3697.4]
  wire [4:0] _T_9159; // @[Mux.scala 31:69:@3698.4]
  wire [4:0] _T_9160; // @[Mux.scala 31:69:@3699.4]
  wire [4:0] select_22; // @[Mux.scala 31:69:@3700.4]
  wire [47:0] _GEN_705; // @[Switch.scala 33:19:@3702.4]
  wire [47:0] _GEN_706; // @[Switch.scala 33:19:@3702.4]
  wire [47:0] _GEN_707; // @[Switch.scala 33:19:@3702.4]
  wire [47:0] _GEN_708; // @[Switch.scala 33:19:@3702.4]
  wire [47:0] _GEN_709; // @[Switch.scala 33:19:@3702.4]
  wire [47:0] _GEN_710; // @[Switch.scala 33:19:@3702.4]
  wire [47:0] _GEN_711; // @[Switch.scala 33:19:@3702.4]
  wire [47:0] _GEN_712; // @[Switch.scala 33:19:@3702.4]
  wire [47:0] _GEN_713; // @[Switch.scala 33:19:@3702.4]
  wire [47:0] _GEN_714; // @[Switch.scala 33:19:@3702.4]
  wire [47:0] _GEN_715; // @[Switch.scala 33:19:@3702.4]
  wire [47:0] _GEN_716; // @[Switch.scala 33:19:@3702.4]
  wire [47:0] _GEN_717; // @[Switch.scala 33:19:@3702.4]
  wire [47:0] _GEN_718; // @[Switch.scala 33:19:@3702.4]
  wire [47:0] _GEN_719; // @[Switch.scala 33:19:@3702.4]
  wire [47:0] _GEN_720; // @[Switch.scala 33:19:@3702.4]
  wire [47:0] _GEN_721; // @[Switch.scala 33:19:@3702.4]
  wire [47:0] _GEN_722; // @[Switch.scala 33:19:@3702.4]
  wire [47:0] _GEN_723; // @[Switch.scala 33:19:@3702.4]
  wire [47:0] _GEN_724; // @[Switch.scala 33:19:@3702.4]
  wire [47:0] _GEN_725; // @[Switch.scala 33:19:@3702.4]
  wire [47:0] _GEN_726; // @[Switch.scala 33:19:@3702.4]
  wire [47:0] _GEN_727; // @[Switch.scala 33:19:@3702.4]
  wire [47:0] _GEN_728; // @[Switch.scala 33:19:@3702.4]
  wire [47:0] _GEN_729; // @[Switch.scala 33:19:@3702.4]
  wire [47:0] _GEN_730; // @[Switch.scala 33:19:@3702.4]
  wire [47:0] _GEN_731; // @[Switch.scala 33:19:@3702.4]
  wire [47:0] _GEN_732; // @[Switch.scala 33:19:@3702.4]
  wire [47:0] _GEN_733; // @[Switch.scala 33:19:@3702.4]
  wire [47:0] _GEN_734; // @[Switch.scala 33:19:@3702.4]
  wire [7:0] _T_9169; // @[Switch.scala 34:32:@3709.4]
  wire [15:0] _T_9177; // @[Switch.scala 34:32:@3717.4]
  wire [7:0] _T_9184; // @[Switch.scala 34:32:@3724.4]
  wire [31:0] _T_9193; // @[Switch.scala 34:32:@3733.4]
  wire  _T_9197; // @[Switch.scala 30:53:@3736.4]
  wire  valid_23_0; // @[Switch.scala 30:36:@3737.4]
  wire  _T_9200; // @[Switch.scala 30:53:@3739.4]
  wire  valid_23_1; // @[Switch.scala 30:36:@3740.4]
  wire  _T_9203; // @[Switch.scala 30:53:@3742.4]
  wire  valid_23_2; // @[Switch.scala 30:36:@3743.4]
  wire  _T_9206; // @[Switch.scala 30:53:@3745.4]
  wire  valid_23_3; // @[Switch.scala 30:36:@3746.4]
  wire  _T_9209; // @[Switch.scala 30:53:@3748.4]
  wire  valid_23_4; // @[Switch.scala 30:36:@3749.4]
  wire  _T_9212; // @[Switch.scala 30:53:@3751.4]
  wire  valid_23_5; // @[Switch.scala 30:36:@3752.4]
  wire  _T_9215; // @[Switch.scala 30:53:@3754.4]
  wire  valid_23_6; // @[Switch.scala 30:36:@3755.4]
  wire  _T_9218; // @[Switch.scala 30:53:@3757.4]
  wire  valid_23_7; // @[Switch.scala 30:36:@3758.4]
  wire  _T_9221; // @[Switch.scala 30:53:@3760.4]
  wire  valid_23_8; // @[Switch.scala 30:36:@3761.4]
  wire  _T_9224; // @[Switch.scala 30:53:@3763.4]
  wire  valid_23_9; // @[Switch.scala 30:36:@3764.4]
  wire  _T_9227; // @[Switch.scala 30:53:@3766.4]
  wire  valid_23_10; // @[Switch.scala 30:36:@3767.4]
  wire  _T_9230; // @[Switch.scala 30:53:@3769.4]
  wire  valid_23_11; // @[Switch.scala 30:36:@3770.4]
  wire  _T_9233; // @[Switch.scala 30:53:@3772.4]
  wire  valid_23_12; // @[Switch.scala 30:36:@3773.4]
  wire  _T_9236; // @[Switch.scala 30:53:@3775.4]
  wire  valid_23_13; // @[Switch.scala 30:36:@3776.4]
  wire  _T_9239; // @[Switch.scala 30:53:@3778.4]
  wire  valid_23_14; // @[Switch.scala 30:36:@3779.4]
  wire  _T_9242; // @[Switch.scala 30:53:@3781.4]
  wire  valid_23_15; // @[Switch.scala 30:36:@3782.4]
  wire  _T_9245; // @[Switch.scala 30:53:@3784.4]
  wire  valid_23_16; // @[Switch.scala 30:36:@3785.4]
  wire  _T_9248; // @[Switch.scala 30:53:@3787.4]
  wire  valid_23_17; // @[Switch.scala 30:36:@3788.4]
  wire  _T_9251; // @[Switch.scala 30:53:@3790.4]
  wire  valid_23_18; // @[Switch.scala 30:36:@3791.4]
  wire  _T_9254; // @[Switch.scala 30:53:@3793.4]
  wire  valid_23_19; // @[Switch.scala 30:36:@3794.4]
  wire  _T_9257; // @[Switch.scala 30:53:@3796.4]
  wire  valid_23_20; // @[Switch.scala 30:36:@3797.4]
  wire  _T_9260; // @[Switch.scala 30:53:@3799.4]
  wire  valid_23_21; // @[Switch.scala 30:36:@3800.4]
  wire  _T_9263; // @[Switch.scala 30:53:@3802.4]
  wire  valid_23_22; // @[Switch.scala 30:36:@3803.4]
  wire  _T_9266; // @[Switch.scala 30:53:@3805.4]
  wire  valid_23_23; // @[Switch.scala 30:36:@3806.4]
  wire  _T_9269; // @[Switch.scala 30:53:@3808.4]
  wire  valid_23_24; // @[Switch.scala 30:36:@3809.4]
  wire  _T_9272; // @[Switch.scala 30:53:@3811.4]
  wire  valid_23_25; // @[Switch.scala 30:36:@3812.4]
  wire  _T_9275; // @[Switch.scala 30:53:@3814.4]
  wire  valid_23_26; // @[Switch.scala 30:36:@3815.4]
  wire  _T_9278; // @[Switch.scala 30:53:@3817.4]
  wire  valid_23_27; // @[Switch.scala 30:36:@3818.4]
  wire  _T_9281; // @[Switch.scala 30:53:@3820.4]
  wire  valid_23_28; // @[Switch.scala 30:36:@3821.4]
  wire  _T_9284; // @[Switch.scala 30:53:@3823.4]
  wire  valid_23_29; // @[Switch.scala 30:36:@3824.4]
  wire  _T_9287; // @[Switch.scala 30:53:@3826.4]
  wire  valid_23_30; // @[Switch.scala 30:36:@3827.4]
  wire  _T_9290; // @[Switch.scala 30:53:@3829.4]
  wire  valid_23_31; // @[Switch.scala 30:36:@3830.4]
  wire [4:0] _T_9324; // @[Mux.scala 31:69:@3832.4]
  wire [4:0] _T_9325; // @[Mux.scala 31:69:@3833.4]
  wire [4:0] _T_9326; // @[Mux.scala 31:69:@3834.4]
  wire [4:0] _T_9327; // @[Mux.scala 31:69:@3835.4]
  wire [4:0] _T_9328; // @[Mux.scala 31:69:@3836.4]
  wire [4:0] _T_9329; // @[Mux.scala 31:69:@3837.4]
  wire [4:0] _T_9330; // @[Mux.scala 31:69:@3838.4]
  wire [4:0] _T_9331; // @[Mux.scala 31:69:@3839.4]
  wire [4:0] _T_9332; // @[Mux.scala 31:69:@3840.4]
  wire [4:0] _T_9333; // @[Mux.scala 31:69:@3841.4]
  wire [4:0] _T_9334; // @[Mux.scala 31:69:@3842.4]
  wire [4:0] _T_9335; // @[Mux.scala 31:69:@3843.4]
  wire [4:0] _T_9336; // @[Mux.scala 31:69:@3844.4]
  wire [4:0] _T_9337; // @[Mux.scala 31:69:@3845.4]
  wire [4:0] _T_9338; // @[Mux.scala 31:69:@3846.4]
  wire [4:0] _T_9339; // @[Mux.scala 31:69:@3847.4]
  wire [4:0] _T_9340; // @[Mux.scala 31:69:@3848.4]
  wire [4:0] _T_9341; // @[Mux.scala 31:69:@3849.4]
  wire [4:0] _T_9342; // @[Mux.scala 31:69:@3850.4]
  wire [4:0] _T_9343; // @[Mux.scala 31:69:@3851.4]
  wire [4:0] _T_9344; // @[Mux.scala 31:69:@3852.4]
  wire [4:0] _T_9345; // @[Mux.scala 31:69:@3853.4]
  wire [4:0] _T_9346; // @[Mux.scala 31:69:@3854.4]
  wire [4:0] _T_9347; // @[Mux.scala 31:69:@3855.4]
  wire [4:0] _T_9348; // @[Mux.scala 31:69:@3856.4]
  wire [4:0] _T_9349; // @[Mux.scala 31:69:@3857.4]
  wire [4:0] _T_9350; // @[Mux.scala 31:69:@3858.4]
  wire [4:0] _T_9351; // @[Mux.scala 31:69:@3859.4]
  wire [4:0] _T_9352; // @[Mux.scala 31:69:@3860.4]
  wire [4:0] _T_9353; // @[Mux.scala 31:69:@3861.4]
  wire [4:0] select_23; // @[Mux.scala 31:69:@3862.4]
  wire [47:0] _GEN_737; // @[Switch.scala 33:19:@3864.4]
  wire [47:0] _GEN_738; // @[Switch.scala 33:19:@3864.4]
  wire [47:0] _GEN_739; // @[Switch.scala 33:19:@3864.4]
  wire [47:0] _GEN_740; // @[Switch.scala 33:19:@3864.4]
  wire [47:0] _GEN_741; // @[Switch.scala 33:19:@3864.4]
  wire [47:0] _GEN_742; // @[Switch.scala 33:19:@3864.4]
  wire [47:0] _GEN_743; // @[Switch.scala 33:19:@3864.4]
  wire [47:0] _GEN_744; // @[Switch.scala 33:19:@3864.4]
  wire [47:0] _GEN_745; // @[Switch.scala 33:19:@3864.4]
  wire [47:0] _GEN_746; // @[Switch.scala 33:19:@3864.4]
  wire [47:0] _GEN_747; // @[Switch.scala 33:19:@3864.4]
  wire [47:0] _GEN_748; // @[Switch.scala 33:19:@3864.4]
  wire [47:0] _GEN_749; // @[Switch.scala 33:19:@3864.4]
  wire [47:0] _GEN_750; // @[Switch.scala 33:19:@3864.4]
  wire [47:0] _GEN_751; // @[Switch.scala 33:19:@3864.4]
  wire [47:0] _GEN_752; // @[Switch.scala 33:19:@3864.4]
  wire [47:0] _GEN_753; // @[Switch.scala 33:19:@3864.4]
  wire [47:0] _GEN_754; // @[Switch.scala 33:19:@3864.4]
  wire [47:0] _GEN_755; // @[Switch.scala 33:19:@3864.4]
  wire [47:0] _GEN_756; // @[Switch.scala 33:19:@3864.4]
  wire [47:0] _GEN_757; // @[Switch.scala 33:19:@3864.4]
  wire [47:0] _GEN_758; // @[Switch.scala 33:19:@3864.4]
  wire [47:0] _GEN_759; // @[Switch.scala 33:19:@3864.4]
  wire [47:0] _GEN_760; // @[Switch.scala 33:19:@3864.4]
  wire [47:0] _GEN_761; // @[Switch.scala 33:19:@3864.4]
  wire [47:0] _GEN_762; // @[Switch.scala 33:19:@3864.4]
  wire [47:0] _GEN_763; // @[Switch.scala 33:19:@3864.4]
  wire [47:0] _GEN_764; // @[Switch.scala 33:19:@3864.4]
  wire [47:0] _GEN_765; // @[Switch.scala 33:19:@3864.4]
  wire [47:0] _GEN_766; // @[Switch.scala 33:19:@3864.4]
  wire [7:0] _T_9362; // @[Switch.scala 34:32:@3871.4]
  wire [15:0] _T_9370; // @[Switch.scala 34:32:@3879.4]
  wire [7:0] _T_9377; // @[Switch.scala 34:32:@3886.4]
  wire [31:0] _T_9386; // @[Switch.scala 34:32:@3895.4]
  wire  _T_9390; // @[Switch.scala 30:53:@3898.4]
  wire  valid_24_0; // @[Switch.scala 30:36:@3899.4]
  wire  _T_9393; // @[Switch.scala 30:53:@3901.4]
  wire  valid_24_1; // @[Switch.scala 30:36:@3902.4]
  wire  _T_9396; // @[Switch.scala 30:53:@3904.4]
  wire  valid_24_2; // @[Switch.scala 30:36:@3905.4]
  wire  _T_9399; // @[Switch.scala 30:53:@3907.4]
  wire  valid_24_3; // @[Switch.scala 30:36:@3908.4]
  wire  _T_9402; // @[Switch.scala 30:53:@3910.4]
  wire  valid_24_4; // @[Switch.scala 30:36:@3911.4]
  wire  _T_9405; // @[Switch.scala 30:53:@3913.4]
  wire  valid_24_5; // @[Switch.scala 30:36:@3914.4]
  wire  _T_9408; // @[Switch.scala 30:53:@3916.4]
  wire  valid_24_6; // @[Switch.scala 30:36:@3917.4]
  wire  _T_9411; // @[Switch.scala 30:53:@3919.4]
  wire  valid_24_7; // @[Switch.scala 30:36:@3920.4]
  wire  _T_9414; // @[Switch.scala 30:53:@3922.4]
  wire  valid_24_8; // @[Switch.scala 30:36:@3923.4]
  wire  _T_9417; // @[Switch.scala 30:53:@3925.4]
  wire  valid_24_9; // @[Switch.scala 30:36:@3926.4]
  wire  _T_9420; // @[Switch.scala 30:53:@3928.4]
  wire  valid_24_10; // @[Switch.scala 30:36:@3929.4]
  wire  _T_9423; // @[Switch.scala 30:53:@3931.4]
  wire  valid_24_11; // @[Switch.scala 30:36:@3932.4]
  wire  _T_9426; // @[Switch.scala 30:53:@3934.4]
  wire  valid_24_12; // @[Switch.scala 30:36:@3935.4]
  wire  _T_9429; // @[Switch.scala 30:53:@3937.4]
  wire  valid_24_13; // @[Switch.scala 30:36:@3938.4]
  wire  _T_9432; // @[Switch.scala 30:53:@3940.4]
  wire  valid_24_14; // @[Switch.scala 30:36:@3941.4]
  wire  _T_9435; // @[Switch.scala 30:53:@3943.4]
  wire  valid_24_15; // @[Switch.scala 30:36:@3944.4]
  wire  _T_9438; // @[Switch.scala 30:53:@3946.4]
  wire  valid_24_16; // @[Switch.scala 30:36:@3947.4]
  wire  _T_9441; // @[Switch.scala 30:53:@3949.4]
  wire  valid_24_17; // @[Switch.scala 30:36:@3950.4]
  wire  _T_9444; // @[Switch.scala 30:53:@3952.4]
  wire  valid_24_18; // @[Switch.scala 30:36:@3953.4]
  wire  _T_9447; // @[Switch.scala 30:53:@3955.4]
  wire  valid_24_19; // @[Switch.scala 30:36:@3956.4]
  wire  _T_9450; // @[Switch.scala 30:53:@3958.4]
  wire  valid_24_20; // @[Switch.scala 30:36:@3959.4]
  wire  _T_9453; // @[Switch.scala 30:53:@3961.4]
  wire  valid_24_21; // @[Switch.scala 30:36:@3962.4]
  wire  _T_9456; // @[Switch.scala 30:53:@3964.4]
  wire  valid_24_22; // @[Switch.scala 30:36:@3965.4]
  wire  _T_9459; // @[Switch.scala 30:53:@3967.4]
  wire  valid_24_23; // @[Switch.scala 30:36:@3968.4]
  wire  _T_9462; // @[Switch.scala 30:53:@3970.4]
  wire  valid_24_24; // @[Switch.scala 30:36:@3971.4]
  wire  _T_9465; // @[Switch.scala 30:53:@3973.4]
  wire  valid_24_25; // @[Switch.scala 30:36:@3974.4]
  wire  _T_9468; // @[Switch.scala 30:53:@3976.4]
  wire  valid_24_26; // @[Switch.scala 30:36:@3977.4]
  wire  _T_9471; // @[Switch.scala 30:53:@3979.4]
  wire  valid_24_27; // @[Switch.scala 30:36:@3980.4]
  wire  _T_9474; // @[Switch.scala 30:53:@3982.4]
  wire  valid_24_28; // @[Switch.scala 30:36:@3983.4]
  wire  _T_9477; // @[Switch.scala 30:53:@3985.4]
  wire  valid_24_29; // @[Switch.scala 30:36:@3986.4]
  wire  _T_9480; // @[Switch.scala 30:53:@3988.4]
  wire  valid_24_30; // @[Switch.scala 30:36:@3989.4]
  wire  _T_9483; // @[Switch.scala 30:53:@3991.4]
  wire  valid_24_31; // @[Switch.scala 30:36:@3992.4]
  wire [4:0] _T_9517; // @[Mux.scala 31:69:@3994.4]
  wire [4:0] _T_9518; // @[Mux.scala 31:69:@3995.4]
  wire [4:0] _T_9519; // @[Mux.scala 31:69:@3996.4]
  wire [4:0] _T_9520; // @[Mux.scala 31:69:@3997.4]
  wire [4:0] _T_9521; // @[Mux.scala 31:69:@3998.4]
  wire [4:0] _T_9522; // @[Mux.scala 31:69:@3999.4]
  wire [4:0] _T_9523; // @[Mux.scala 31:69:@4000.4]
  wire [4:0] _T_9524; // @[Mux.scala 31:69:@4001.4]
  wire [4:0] _T_9525; // @[Mux.scala 31:69:@4002.4]
  wire [4:0] _T_9526; // @[Mux.scala 31:69:@4003.4]
  wire [4:0] _T_9527; // @[Mux.scala 31:69:@4004.4]
  wire [4:0] _T_9528; // @[Mux.scala 31:69:@4005.4]
  wire [4:0] _T_9529; // @[Mux.scala 31:69:@4006.4]
  wire [4:0] _T_9530; // @[Mux.scala 31:69:@4007.4]
  wire [4:0] _T_9531; // @[Mux.scala 31:69:@4008.4]
  wire [4:0] _T_9532; // @[Mux.scala 31:69:@4009.4]
  wire [4:0] _T_9533; // @[Mux.scala 31:69:@4010.4]
  wire [4:0] _T_9534; // @[Mux.scala 31:69:@4011.4]
  wire [4:0] _T_9535; // @[Mux.scala 31:69:@4012.4]
  wire [4:0] _T_9536; // @[Mux.scala 31:69:@4013.4]
  wire [4:0] _T_9537; // @[Mux.scala 31:69:@4014.4]
  wire [4:0] _T_9538; // @[Mux.scala 31:69:@4015.4]
  wire [4:0] _T_9539; // @[Mux.scala 31:69:@4016.4]
  wire [4:0] _T_9540; // @[Mux.scala 31:69:@4017.4]
  wire [4:0] _T_9541; // @[Mux.scala 31:69:@4018.4]
  wire [4:0] _T_9542; // @[Mux.scala 31:69:@4019.4]
  wire [4:0] _T_9543; // @[Mux.scala 31:69:@4020.4]
  wire [4:0] _T_9544; // @[Mux.scala 31:69:@4021.4]
  wire [4:0] _T_9545; // @[Mux.scala 31:69:@4022.4]
  wire [4:0] _T_9546; // @[Mux.scala 31:69:@4023.4]
  wire [4:0] select_24; // @[Mux.scala 31:69:@4024.4]
  wire [47:0] _GEN_769; // @[Switch.scala 33:19:@4026.4]
  wire [47:0] _GEN_770; // @[Switch.scala 33:19:@4026.4]
  wire [47:0] _GEN_771; // @[Switch.scala 33:19:@4026.4]
  wire [47:0] _GEN_772; // @[Switch.scala 33:19:@4026.4]
  wire [47:0] _GEN_773; // @[Switch.scala 33:19:@4026.4]
  wire [47:0] _GEN_774; // @[Switch.scala 33:19:@4026.4]
  wire [47:0] _GEN_775; // @[Switch.scala 33:19:@4026.4]
  wire [47:0] _GEN_776; // @[Switch.scala 33:19:@4026.4]
  wire [47:0] _GEN_777; // @[Switch.scala 33:19:@4026.4]
  wire [47:0] _GEN_778; // @[Switch.scala 33:19:@4026.4]
  wire [47:0] _GEN_779; // @[Switch.scala 33:19:@4026.4]
  wire [47:0] _GEN_780; // @[Switch.scala 33:19:@4026.4]
  wire [47:0] _GEN_781; // @[Switch.scala 33:19:@4026.4]
  wire [47:0] _GEN_782; // @[Switch.scala 33:19:@4026.4]
  wire [47:0] _GEN_783; // @[Switch.scala 33:19:@4026.4]
  wire [47:0] _GEN_784; // @[Switch.scala 33:19:@4026.4]
  wire [47:0] _GEN_785; // @[Switch.scala 33:19:@4026.4]
  wire [47:0] _GEN_786; // @[Switch.scala 33:19:@4026.4]
  wire [47:0] _GEN_787; // @[Switch.scala 33:19:@4026.4]
  wire [47:0] _GEN_788; // @[Switch.scala 33:19:@4026.4]
  wire [47:0] _GEN_789; // @[Switch.scala 33:19:@4026.4]
  wire [47:0] _GEN_790; // @[Switch.scala 33:19:@4026.4]
  wire [47:0] _GEN_791; // @[Switch.scala 33:19:@4026.4]
  wire [47:0] _GEN_792; // @[Switch.scala 33:19:@4026.4]
  wire [47:0] _GEN_793; // @[Switch.scala 33:19:@4026.4]
  wire [47:0] _GEN_794; // @[Switch.scala 33:19:@4026.4]
  wire [47:0] _GEN_795; // @[Switch.scala 33:19:@4026.4]
  wire [47:0] _GEN_796; // @[Switch.scala 33:19:@4026.4]
  wire [47:0] _GEN_797; // @[Switch.scala 33:19:@4026.4]
  wire [47:0] _GEN_798; // @[Switch.scala 33:19:@4026.4]
  wire [7:0] _T_9555; // @[Switch.scala 34:32:@4033.4]
  wire [15:0] _T_9563; // @[Switch.scala 34:32:@4041.4]
  wire [7:0] _T_9570; // @[Switch.scala 34:32:@4048.4]
  wire [31:0] _T_9579; // @[Switch.scala 34:32:@4057.4]
  wire  _T_9583; // @[Switch.scala 30:53:@4060.4]
  wire  valid_25_0; // @[Switch.scala 30:36:@4061.4]
  wire  _T_9586; // @[Switch.scala 30:53:@4063.4]
  wire  valid_25_1; // @[Switch.scala 30:36:@4064.4]
  wire  _T_9589; // @[Switch.scala 30:53:@4066.4]
  wire  valid_25_2; // @[Switch.scala 30:36:@4067.4]
  wire  _T_9592; // @[Switch.scala 30:53:@4069.4]
  wire  valid_25_3; // @[Switch.scala 30:36:@4070.4]
  wire  _T_9595; // @[Switch.scala 30:53:@4072.4]
  wire  valid_25_4; // @[Switch.scala 30:36:@4073.4]
  wire  _T_9598; // @[Switch.scala 30:53:@4075.4]
  wire  valid_25_5; // @[Switch.scala 30:36:@4076.4]
  wire  _T_9601; // @[Switch.scala 30:53:@4078.4]
  wire  valid_25_6; // @[Switch.scala 30:36:@4079.4]
  wire  _T_9604; // @[Switch.scala 30:53:@4081.4]
  wire  valid_25_7; // @[Switch.scala 30:36:@4082.4]
  wire  _T_9607; // @[Switch.scala 30:53:@4084.4]
  wire  valid_25_8; // @[Switch.scala 30:36:@4085.4]
  wire  _T_9610; // @[Switch.scala 30:53:@4087.4]
  wire  valid_25_9; // @[Switch.scala 30:36:@4088.4]
  wire  _T_9613; // @[Switch.scala 30:53:@4090.4]
  wire  valid_25_10; // @[Switch.scala 30:36:@4091.4]
  wire  _T_9616; // @[Switch.scala 30:53:@4093.4]
  wire  valid_25_11; // @[Switch.scala 30:36:@4094.4]
  wire  _T_9619; // @[Switch.scala 30:53:@4096.4]
  wire  valid_25_12; // @[Switch.scala 30:36:@4097.4]
  wire  _T_9622; // @[Switch.scala 30:53:@4099.4]
  wire  valid_25_13; // @[Switch.scala 30:36:@4100.4]
  wire  _T_9625; // @[Switch.scala 30:53:@4102.4]
  wire  valid_25_14; // @[Switch.scala 30:36:@4103.4]
  wire  _T_9628; // @[Switch.scala 30:53:@4105.4]
  wire  valid_25_15; // @[Switch.scala 30:36:@4106.4]
  wire  _T_9631; // @[Switch.scala 30:53:@4108.4]
  wire  valid_25_16; // @[Switch.scala 30:36:@4109.4]
  wire  _T_9634; // @[Switch.scala 30:53:@4111.4]
  wire  valid_25_17; // @[Switch.scala 30:36:@4112.4]
  wire  _T_9637; // @[Switch.scala 30:53:@4114.4]
  wire  valid_25_18; // @[Switch.scala 30:36:@4115.4]
  wire  _T_9640; // @[Switch.scala 30:53:@4117.4]
  wire  valid_25_19; // @[Switch.scala 30:36:@4118.4]
  wire  _T_9643; // @[Switch.scala 30:53:@4120.4]
  wire  valid_25_20; // @[Switch.scala 30:36:@4121.4]
  wire  _T_9646; // @[Switch.scala 30:53:@4123.4]
  wire  valid_25_21; // @[Switch.scala 30:36:@4124.4]
  wire  _T_9649; // @[Switch.scala 30:53:@4126.4]
  wire  valid_25_22; // @[Switch.scala 30:36:@4127.4]
  wire  _T_9652; // @[Switch.scala 30:53:@4129.4]
  wire  valid_25_23; // @[Switch.scala 30:36:@4130.4]
  wire  _T_9655; // @[Switch.scala 30:53:@4132.4]
  wire  valid_25_24; // @[Switch.scala 30:36:@4133.4]
  wire  _T_9658; // @[Switch.scala 30:53:@4135.4]
  wire  valid_25_25; // @[Switch.scala 30:36:@4136.4]
  wire  _T_9661; // @[Switch.scala 30:53:@4138.4]
  wire  valid_25_26; // @[Switch.scala 30:36:@4139.4]
  wire  _T_9664; // @[Switch.scala 30:53:@4141.4]
  wire  valid_25_27; // @[Switch.scala 30:36:@4142.4]
  wire  _T_9667; // @[Switch.scala 30:53:@4144.4]
  wire  valid_25_28; // @[Switch.scala 30:36:@4145.4]
  wire  _T_9670; // @[Switch.scala 30:53:@4147.4]
  wire  valid_25_29; // @[Switch.scala 30:36:@4148.4]
  wire  _T_9673; // @[Switch.scala 30:53:@4150.4]
  wire  valid_25_30; // @[Switch.scala 30:36:@4151.4]
  wire  _T_9676; // @[Switch.scala 30:53:@4153.4]
  wire  valid_25_31; // @[Switch.scala 30:36:@4154.4]
  wire [4:0] _T_9710; // @[Mux.scala 31:69:@4156.4]
  wire [4:0] _T_9711; // @[Mux.scala 31:69:@4157.4]
  wire [4:0] _T_9712; // @[Mux.scala 31:69:@4158.4]
  wire [4:0] _T_9713; // @[Mux.scala 31:69:@4159.4]
  wire [4:0] _T_9714; // @[Mux.scala 31:69:@4160.4]
  wire [4:0] _T_9715; // @[Mux.scala 31:69:@4161.4]
  wire [4:0] _T_9716; // @[Mux.scala 31:69:@4162.4]
  wire [4:0] _T_9717; // @[Mux.scala 31:69:@4163.4]
  wire [4:0] _T_9718; // @[Mux.scala 31:69:@4164.4]
  wire [4:0] _T_9719; // @[Mux.scala 31:69:@4165.4]
  wire [4:0] _T_9720; // @[Mux.scala 31:69:@4166.4]
  wire [4:0] _T_9721; // @[Mux.scala 31:69:@4167.4]
  wire [4:0] _T_9722; // @[Mux.scala 31:69:@4168.4]
  wire [4:0] _T_9723; // @[Mux.scala 31:69:@4169.4]
  wire [4:0] _T_9724; // @[Mux.scala 31:69:@4170.4]
  wire [4:0] _T_9725; // @[Mux.scala 31:69:@4171.4]
  wire [4:0] _T_9726; // @[Mux.scala 31:69:@4172.4]
  wire [4:0] _T_9727; // @[Mux.scala 31:69:@4173.4]
  wire [4:0] _T_9728; // @[Mux.scala 31:69:@4174.4]
  wire [4:0] _T_9729; // @[Mux.scala 31:69:@4175.4]
  wire [4:0] _T_9730; // @[Mux.scala 31:69:@4176.4]
  wire [4:0] _T_9731; // @[Mux.scala 31:69:@4177.4]
  wire [4:0] _T_9732; // @[Mux.scala 31:69:@4178.4]
  wire [4:0] _T_9733; // @[Mux.scala 31:69:@4179.4]
  wire [4:0] _T_9734; // @[Mux.scala 31:69:@4180.4]
  wire [4:0] _T_9735; // @[Mux.scala 31:69:@4181.4]
  wire [4:0] _T_9736; // @[Mux.scala 31:69:@4182.4]
  wire [4:0] _T_9737; // @[Mux.scala 31:69:@4183.4]
  wire [4:0] _T_9738; // @[Mux.scala 31:69:@4184.4]
  wire [4:0] _T_9739; // @[Mux.scala 31:69:@4185.4]
  wire [4:0] select_25; // @[Mux.scala 31:69:@4186.4]
  wire [47:0] _GEN_801; // @[Switch.scala 33:19:@4188.4]
  wire [47:0] _GEN_802; // @[Switch.scala 33:19:@4188.4]
  wire [47:0] _GEN_803; // @[Switch.scala 33:19:@4188.4]
  wire [47:0] _GEN_804; // @[Switch.scala 33:19:@4188.4]
  wire [47:0] _GEN_805; // @[Switch.scala 33:19:@4188.4]
  wire [47:0] _GEN_806; // @[Switch.scala 33:19:@4188.4]
  wire [47:0] _GEN_807; // @[Switch.scala 33:19:@4188.4]
  wire [47:0] _GEN_808; // @[Switch.scala 33:19:@4188.4]
  wire [47:0] _GEN_809; // @[Switch.scala 33:19:@4188.4]
  wire [47:0] _GEN_810; // @[Switch.scala 33:19:@4188.4]
  wire [47:0] _GEN_811; // @[Switch.scala 33:19:@4188.4]
  wire [47:0] _GEN_812; // @[Switch.scala 33:19:@4188.4]
  wire [47:0] _GEN_813; // @[Switch.scala 33:19:@4188.4]
  wire [47:0] _GEN_814; // @[Switch.scala 33:19:@4188.4]
  wire [47:0] _GEN_815; // @[Switch.scala 33:19:@4188.4]
  wire [47:0] _GEN_816; // @[Switch.scala 33:19:@4188.4]
  wire [47:0] _GEN_817; // @[Switch.scala 33:19:@4188.4]
  wire [47:0] _GEN_818; // @[Switch.scala 33:19:@4188.4]
  wire [47:0] _GEN_819; // @[Switch.scala 33:19:@4188.4]
  wire [47:0] _GEN_820; // @[Switch.scala 33:19:@4188.4]
  wire [47:0] _GEN_821; // @[Switch.scala 33:19:@4188.4]
  wire [47:0] _GEN_822; // @[Switch.scala 33:19:@4188.4]
  wire [47:0] _GEN_823; // @[Switch.scala 33:19:@4188.4]
  wire [47:0] _GEN_824; // @[Switch.scala 33:19:@4188.4]
  wire [47:0] _GEN_825; // @[Switch.scala 33:19:@4188.4]
  wire [47:0] _GEN_826; // @[Switch.scala 33:19:@4188.4]
  wire [47:0] _GEN_827; // @[Switch.scala 33:19:@4188.4]
  wire [47:0] _GEN_828; // @[Switch.scala 33:19:@4188.4]
  wire [47:0] _GEN_829; // @[Switch.scala 33:19:@4188.4]
  wire [47:0] _GEN_830; // @[Switch.scala 33:19:@4188.4]
  wire [7:0] _T_9748; // @[Switch.scala 34:32:@4195.4]
  wire [15:0] _T_9756; // @[Switch.scala 34:32:@4203.4]
  wire [7:0] _T_9763; // @[Switch.scala 34:32:@4210.4]
  wire [31:0] _T_9772; // @[Switch.scala 34:32:@4219.4]
  wire  _T_9776; // @[Switch.scala 30:53:@4222.4]
  wire  valid_26_0; // @[Switch.scala 30:36:@4223.4]
  wire  _T_9779; // @[Switch.scala 30:53:@4225.4]
  wire  valid_26_1; // @[Switch.scala 30:36:@4226.4]
  wire  _T_9782; // @[Switch.scala 30:53:@4228.4]
  wire  valid_26_2; // @[Switch.scala 30:36:@4229.4]
  wire  _T_9785; // @[Switch.scala 30:53:@4231.4]
  wire  valid_26_3; // @[Switch.scala 30:36:@4232.4]
  wire  _T_9788; // @[Switch.scala 30:53:@4234.4]
  wire  valid_26_4; // @[Switch.scala 30:36:@4235.4]
  wire  _T_9791; // @[Switch.scala 30:53:@4237.4]
  wire  valid_26_5; // @[Switch.scala 30:36:@4238.4]
  wire  _T_9794; // @[Switch.scala 30:53:@4240.4]
  wire  valid_26_6; // @[Switch.scala 30:36:@4241.4]
  wire  _T_9797; // @[Switch.scala 30:53:@4243.4]
  wire  valid_26_7; // @[Switch.scala 30:36:@4244.4]
  wire  _T_9800; // @[Switch.scala 30:53:@4246.4]
  wire  valid_26_8; // @[Switch.scala 30:36:@4247.4]
  wire  _T_9803; // @[Switch.scala 30:53:@4249.4]
  wire  valid_26_9; // @[Switch.scala 30:36:@4250.4]
  wire  _T_9806; // @[Switch.scala 30:53:@4252.4]
  wire  valid_26_10; // @[Switch.scala 30:36:@4253.4]
  wire  _T_9809; // @[Switch.scala 30:53:@4255.4]
  wire  valid_26_11; // @[Switch.scala 30:36:@4256.4]
  wire  _T_9812; // @[Switch.scala 30:53:@4258.4]
  wire  valid_26_12; // @[Switch.scala 30:36:@4259.4]
  wire  _T_9815; // @[Switch.scala 30:53:@4261.4]
  wire  valid_26_13; // @[Switch.scala 30:36:@4262.4]
  wire  _T_9818; // @[Switch.scala 30:53:@4264.4]
  wire  valid_26_14; // @[Switch.scala 30:36:@4265.4]
  wire  _T_9821; // @[Switch.scala 30:53:@4267.4]
  wire  valid_26_15; // @[Switch.scala 30:36:@4268.4]
  wire  _T_9824; // @[Switch.scala 30:53:@4270.4]
  wire  valid_26_16; // @[Switch.scala 30:36:@4271.4]
  wire  _T_9827; // @[Switch.scala 30:53:@4273.4]
  wire  valid_26_17; // @[Switch.scala 30:36:@4274.4]
  wire  _T_9830; // @[Switch.scala 30:53:@4276.4]
  wire  valid_26_18; // @[Switch.scala 30:36:@4277.4]
  wire  _T_9833; // @[Switch.scala 30:53:@4279.4]
  wire  valid_26_19; // @[Switch.scala 30:36:@4280.4]
  wire  _T_9836; // @[Switch.scala 30:53:@4282.4]
  wire  valid_26_20; // @[Switch.scala 30:36:@4283.4]
  wire  _T_9839; // @[Switch.scala 30:53:@4285.4]
  wire  valid_26_21; // @[Switch.scala 30:36:@4286.4]
  wire  _T_9842; // @[Switch.scala 30:53:@4288.4]
  wire  valid_26_22; // @[Switch.scala 30:36:@4289.4]
  wire  _T_9845; // @[Switch.scala 30:53:@4291.4]
  wire  valid_26_23; // @[Switch.scala 30:36:@4292.4]
  wire  _T_9848; // @[Switch.scala 30:53:@4294.4]
  wire  valid_26_24; // @[Switch.scala 30:36:@4295.4]
  wire  _T_9851; // @[Switch.scala 30:53:@4297.4]
  wire  valid_26_25; // @[Switch.scala 30:36:@4298.4]
  wire  _T_9854; // @[Switch.scala 30:53:@4300.4]
  wire  valid_26_26; // @[Switch.scala 30:36:@4301.4]
  wire  _T_9857; // @[Switch.scala 30:53:@4303.4]
  wire  valid_26_27; // @[Switch.scala 30:36:@4304.4]
  wire  _T_9860; // @[Switch.scala 30:53:@4306.4]
  wire  valid_26_28; // @[Switch.scala 30:36:@4307.4]
  wire  _T_9863; // @[Switch.scala 30:53:@4309.4]
  wire  valid_26_29; // @[Switch.scala 30:36:@4310.4]
  wire  _T_9866; // @[Switch.scala 30:53:@4312.4]
  wire  valid_26_30; // @[Switch.scala 30:36:@4313.4]
  wire  _T_9869; // @[Switch.scala 30:53:@4315.4]
  wire  valid_26_31; // @[Switch.scala 30:36:@4316.4]
  wire [4:0] _T_9903; // @[Mux.scala 31:69:@4318.4]
  wire [4:0] _T_9904; // @[Mux.scala 31:69:@4319.4]
  wire [4:0] _T_9905; // @[Mux.scala 31:69:@4320.4]
  wire [4:0] _T_9906; // @[Mux.scala 31:69:@4321.4]
  wire [4:0] _T_9907; // @[Mux.scala 31:69:@4322.4]
  wire [4:0] _T_9908; // @[Mux.scala 31:69:@4323.4]
  wire [4:0] _T_9909; // @[Mux.scala 31:69:@4324.4]
  wire [4:0] _T_9910; // @[Mux.scala 31:69:@4325.4]
  wire [4:0] _T_9911; // @[Mux.scala 31:69:@4326.4]
  wire [4:0] _T_9912; // @[Mux.scala 31:69:@4327.4]
  wire [4:0] _T_9913; // @[Mux.scala 31:69:@4328.4]
  wire [4:0] _T_9914; // @[Mux.scala 31:69:@4329.4]
  wire [4:0] _T_9915; // @[Mux.scala 31:69:@4330.4]
  wire [4:0] _T_9916; // @[Mux.scala 31:69:@4331.4]
  wire [4:0] _T_9917; // @[Mux.scala 31:69:@4332.4]
  wire [4:0] _T_9918; // @[Mux.scala 31:69:@4333.4]
  wire [4:0] _T_9919; // @[Mux.scala 31:69:@4334.4]
  wire [4:0] _T_9920; // @[Mux.scala 31:69:@4335.4]
  wire [4:0] _T_9921; // @[Mux.scala 31:69:@4336.4]
  wire [4:0] _T_9922; // @[Mux.scala 31:69:@4337.4]
  wire [4:0] _T_9923; // @[Mux.scala 31:69:@4338.4]
  wire [4:0] _T_9924; // @[Mux.scala 31:69:@4339.4]
  wire [4:0] _T_9925; // @[Mux.scala 31:69:@4340.4]
  wire [4:0] _T_9926; // @[Mux.scala 31:69:@4341.4]
  wire [4:0] _T_9927; // @[Mux.scala 31:69:@4342.4]
  wire [4:0] _T_9928; // @[Mux.scala 31:69:@4343.4]
  wire [4:0] _T_9929; // @[Mux.scala 31:69:@4344.4]
  wire [4:0] _T_9930; // @[Mux.scala 31:69:@4345.4]
  wire [4:0] _T_9931; // @[Mux.scala 31:69:@4346.4]
  wire [4:0] _T_9932; // @[Mux.scala 31:69:@4347.4]
  wire [4:0] select_26; // @[Mux.scala 31:69:@4348.4]
  wire [47:0] _GEN_833; // @[Switch.scala 33:19:@4350.4]
  wire [47:0] _GEN_834; // @[Switch.scala 33:19:@4350.4]
  wire [47:0] _GEN_835; // @[Switch.scala 33:19:@4350.4]
  wire [47:0] _GEN_836; // @[Switch.scala 33:19:@4350.4]
  wire [47:0] _GEN_837; // @[Switch.scala 33:19:@4350.4]
  wire [47:0] _GEN_838; // @[Switch.scala 33:19:@4350.4]
  wire [47:0] _GEN_839; // @[Switch.scala 33:19:@4350.4]
  wire [47:0] _GEN_840; // @[Switch.scala 33:19:@4350.4]
  wire [47:0] _GEN_841; // @[Switch.scala 33:19:@4350.4]
  wire [47:0] _GEN_842; // @[Switch.scala 33:19:@4350.4]
  wire [47:0] _GEN_843; // @[Switch.scala 33:19:@4350.4]
  wire [47:0] _GEN_844; // @[Switch.scala 33:19:@4350.4]
  wire [47:0] _GEN_845; // @[Switch.scala 33:19:@4350.4]
  wire [47:0] _GEN_846; // @[Switch.scala 33:19:@4350.4]
  wire [47:0] _GEN_847; // @[Switch.scala 33:19:@4350.4]
  wire [47:0] _GEN_848; // @[Switch.scala 33:19:@4350.4]
  wire [47:0] _GEN_849; // @[Switch.scala 33:19:@4350.4]
  wire [47:0] _GEN_850; // @[Switch.scala 33:19:@4350.4]
  wire [47:0] _GEN_851; // @[Switch.scala 33:19:@4350.4]
  wire [47:0] _GEN_852; // @[Switch.scala 33:19:@4350.4]
  wire [47:0] _GEN_853; // @[Switch.scala 33:19:@4350.4]
  wire [47:0] _GEN_854; // @[Switch.scala 33:19:@4350.4]
  wire [47:0] _GEN_855; // @[Switch.scala 33:19:@4350.4]
  wire [47:0] _GEN_856; // @[Switch.scala 33:19:@4350.4]
  wire [47:0] _GEN_857; // @[Switch.scala 33:19:@4350.4]
  wire [47:0] _GEN_858; // @[Switch.scala 33:19:@4350.4]
  wire [47:0] _GEN_859; // @[Switch.scala 33:19:@4350.4]
  wire [47:0] _GEN_860; // @[Switch.scala 33:19:@4350.4]
  wire [47:0] _GEN_861; // @[Switch.scala 33:19:@4350.4]
  wire [47:0] _GEN_862; // @[Switch.scala 33:19:@4350.4]
  wire [7:0] _T_9941; // @[Switch.scala 34:32:@4357.4]
  wire [15:0] _T_9949; // @[Switch.scala 34:32:@4365.4]
  wire [7:0] _T_9956; // @[Switch.scala 34:32:@4372.4]
  wire [31:0] _T_9965; // @[Switch.scala 34:32:@4381.4]
  wire  _T_9969; // @[Switch.scala 30:53:@4384.4]
  wire  valid_27_0; // @[Switch.scala 30:36:@4385.4]
  wire  _T_9972; // @[Switch.scala 30:53:@4387.4]
  wire  valid_27_1; // @[Switch.scala 30:36:@4388.4]
  wire  _T_9975; // @[Switch.scala 30:53:@4390.4]
  wire  valid_27_2; // @[Switch.scala 30:36:@4391.4]
  wire  _T_9978; // @[Switch.scala 30:53:@4393.4]
  wire  valid_27_3; // @[Switch.scala 30:36:@4394.4]
  wire  _T_9981; // @[Switch.scala 30:53:@4396.4]
  wire  valid_27_4; // @[Switch.scala 30:36:@4397.4]
  wire  _T_9984; // @[Switch.scala 30:53:@4399.4]
  wire  valid_27_5; // @[Switch.scala 30:36:@4400.4]
  wire  _T_9987; // @[Switch.scala 30:53:@4402.4]
  wire  valid_27_6; // @[Switch.scala 30:36:@4403.4]
  wire  _T_9990; // @[Switch.scala 30:53:@4405.4]
  wire  valid_27_7; // @[Switch.scala 30:36:@4406.4]
  wire  _T_9993; // @[Switch.scala 30:53:@4408.4]
  wire  valid_27_8; // @[Switch.scala 30:36:@4409.4]
  wire  _T_9996; // @[Switch.scala 30:53:@4411.4]
  wire  valid_27_9; // @[Switch.scala 30:36:@4412.4]
  wire  _T_9999; // @[Switch.scala 30:53:@4414.4]
  wire  valid_27_10; // @[Switch.scala 30:36:@4415.4]
  wire  _T_10002; // @[Switch.scala 30:53:@4417.4]
  wire  valid_27_11; // @[Switch.scala 30:36:@4418.4]
  wire  _T_10005; // @[Switch.scala 30:53:@4420.4]
  wire  valid_27_12; // @[Switch.scala 30:36:@4421.4]
  wire  _T_10008; // @[Switch.scala 30:53:@4423.4]
  wire  valid_27_13; // @[Switch.scala 30:36:@4424.4]
  wire  _T_10011; // @[Switch.scala 30:53:@4426.4]
  wire  valid_27_14; // @[Switch.scala 30:36:@4427.4]
  wire  _T_10014; // @[Switch.scala 30:53:@4429.4]
  wire  valid_27_15; // @[Switch.scala 30:36:@4430.4]
  wire  _T_10017; // @[Switch.scala 30:53:@4432.4]
  wire  valid_27_16; // @[Switch.scala 30:36:@4433.4]
  wire  _T_10020; // @[Switch.scala 30:53:@4435.4]
  wire  valid_27_17; // @[Switch.scala 30:36:@4436.4]
  wire  _T_10023; // @[Switch.scala 30:53:@4438.4]
  wire  valid_27_18; // @[Switch.scala 30:36:@4439.4]
  wire  _T_10026; // @[Switch.scala 30:53:@4441.4]
  wire  valid_27_19; // @[Switch.scala 30:36:@4442.4]
  wire  _T_10029; // @[Switch.scala 30:53:@4444.4]
  wire  valid_27_20; // @[Switch.scala 30:36:@4445.4]
  wire  _T_10032; // @[Switch.scala 30:53:@4447.4]
  wire  valid_27_21; // @[Switch.scala 30:36:@4448.4]
  wire  _T_10035; // @[Switch.scala 30:53:@4450.4]
  wire  valid_27_22; // @[Switch.scala 30:36:@4451.4]
  wire  _T_10038; // @[Switch.scala 30:53:@4453.4]
  wire  valid_27_23; // @[Switch.scala 30:36:@4454.4]
  wire  _T_10041; // @[Switch.scala 30:53:@4456.4]
  wire  valid_27_24; // @[Switch.scala 30:36:@4457.4]
  wire  _T_10044; // @[Switch.scala 30:53:@4459.4]
  wire  valid_27_25; // @[Switch.scala 30:36:@4460.4]
  wire  _T_10047; // @[Switch.scala 30:53:@4462.4]
  wire  valid_27_26; // @[Switch.scala 30:36:@4463.4]
  wire  _T_10050; // @[Switch.scala 30:53:@4465.4]
  wire  valid_27_27; // @[Switch.scala 30:36:@4466.4]
  wire  _T_10053; // @[Switch.scala 30:53:@4468.4]
  wire  valid_27_28; // @[Switch.scala 30:36:@4469.4]
  wire  _T_10056; // @[Switch.scala 30:53:@4471.4]
  wire  valid_27_29; // @[Switch.scala 30:36:@4472.4]
  wire  _T_10059; // @[Switch.scala 30:53:@4474.4]
  wire  valid_27_30; // @[Switch.scala 30:36:@4475.4]
  wire  _T_10062; // @[Switch.scala 30:53:@4477.4]
  wire  valid_27_31; // @[Switch.scala 30:36:@4478.4]
  wire [4:0] _T_10096; // @[Mux.scala 31:69:@4480.4]
  wire [4:0] _T_10097; // @[Mux.scala 31:69:@4481.4]
  wire [4:0] _T_10098; // @[Mux.scala 31:69:@4482.4]
  wire [4:0] _T_10099; // @[Mux.scala 31:69:@4483.4]
  wire [4:0] _T_10100; // @[Mux.scala 31:69:@4484.4]
  wire [4:0] _T_10101; // @[Mux.scala 31:69:@4485.4]
  wire [4:0] _T_10102; // @[Mux.scala 31:69:@4486.4]
  wire [4:0] _T_10103; // @[Mux.scala 31:69:@4487.4]
  wire [4:0] _T_10104; // @[Mux.scala 31:69:@4488.4]
  wire [4:0] _T_10105; // @[Mux.scala 31:69:@4489.4]
  wire [4:0] _T_10106; // @[Mux.scala 31:69:@4490.4]
  wire [4:0] _T_10107; // @[Mux.scala 31:69:@4491.4]
  wire [4:0] _T_10108; // @[Mux.scala 31:69:@4492.4]
  wire [4:0] _T_10109; // @[Mux.scala 31:69:@4493.4]
  wire [4:0] _T_10110; // @[Mux.scala 31:69:@4494.4]
  wire [4:0] _T_10111; // @[Mux.scala 31:69:@4495.4]
  wire [4:0] _T_10112; // @[Mux.scala 31:69:@4496.4]
  wire [4:0] _T_10113; // @[Mux.scala 31:69:@4497.4]
  wire [4:0] _T_10114; // @[Mux.scala 31:69:@4498.4]
  wire [4:0] _T_10115; // @[Mux.scala 31:69:@4499.4]
  wire [4:0] _T_10116; // @[Mux.scala 31:69:@4500.4]
  wire [4:0] _T_10117; // @[Mux.scala 31:69:@4501.4]
  wire [4:0] _T_10118; // @[Mux.scala 31:69:@4502.4]
  wire [4:0] _T_10119; // @[Mux.scala 31:69:@4503.4]
  wire [4:0] _T_10120; // @[Mux.scala 31:69:@4504.4]
  wire [4:0] _T_10121; // @[Mux.scala 31:69:@4505.4]
  wire [4:0] _T_10122; // @[Mux.scala 31:69:@4506.4]
  wire [4:0] _T_10123; // @[Mux.scala 31:69:@4507.4]
  wire [4:0] _T_10124; // @[Mux.scala 31:69:@4508.4]
  wire [4:0] _T_10125; // @[Mux.scala 31:69:@4509.4]
  wire [4:0] select_27; // @[Mux.scala 31:69:@4510.4]
  wire [47:0] _GEN_865; // @[Switch.scala 33:19:@4512.4]
  wire [47:0] _GEN_866; // @[Switch.scala 33:19:@4512.4]
  wire [47:0] _GEN_867; // @[Switch.scala 33:19:@4512.4]
  wire [47:0] _GEN_868; // @[Switch.scala 33:19:@4512.4]
  wire [47:0] _GEN_869; // @[Switch.scala 33:19:@4512.4]
  wire [47:0] _GEN_870; // @[Switch.scala 33:19:@4512.4]
  wire [47:0] _GEN_871; // @[Switch.scala 33:19:@4512.4]
  wire [47:0] _GEN_872; // @[Switch.scala 33:19:@4512.4]
  wire [47:0] _GEN_873; // @[Switch.scala 33:19:@4512.4]
  wire [47:0] _GEN_874; // @[Switch.scala 33:19:@4512.4]
  wire [47:0] _GEN_875; // @[Switch.scala 33:19:@4512.4]
  wire [47:0] _GEN_876; // @[Switch.scala 33:19:@4512.4]
  wire [47:0] _GEN_877; // @[Switch.scala 33:19:@4512.4]
  wire [47:0] _GEN_878; // @[Switch.scala 33:19:@4512.4]
  wire [47:0] _GEN_879; // @[Switch.scala 33:19:@4512.4]
  wire [47:0] _GEN_880; // @[Switch.scala 33:19:@4512.4]
  wire [47:0] _GEN_881; // @[Switch.scala 33:19:@4512.4]
  wire [47:0] _GEN_882; // @[Switch.scala 33:19:@4512.4]
  wire [47:0] _GEN_883; // @[Switch.scala 33:19:@4512.4]
  wire [47:0] _GEN_884; // @[Switch.scala 33:19:@4512.4]
  wire [47:0] _GEN_885; // @[Switch.scala 33:19:@4512.4]
  wire [47:0] _GEN_886; // @[Switch.scala 33:19:@4512.4]
  wire [47:0] _GEN_887; // @[Switch.scala 33:19:@4512.4]
  wire [47:0] _GEN_888; // @[Switch.scala 33:19:@4512.4]
  wire [47:0] _GEN_889; // @[Switch.scala 33:19:@4512.4]
  wire [47:0] _GEN_890; // @[Switch.scala 33:19:@4512.4]
  wire [47:0] _GEN_891; // @[Switch.scala 33:19:@4512.4]
  wire [47:0] _GEN_892; // @[Switch.scala 33:19:@4512.4]
  wire [47:0] _GEN_893; // @[Switch.scala 33:19:@4512.4]
  wire [47:0] _GEN_894; // @[Switch.scala 33:19:@4512.4]
  wire [7:0] _T_10134; // @[Switch.scala 34:32:@4519.4]
  wire [15:0] _T_10142; // @[Switch.scala 34:32:@4527.4]
  wire [7:0] _T_10149; // @[Switch.scala 34:32:@4534.4]
  wire [31:0] _T_10158; // @[Switch.scala 34:32:@4543.4]
  wire  _T_10162; // @[Switch.scala 30:53:@4546.4]
  wire  valid_28_0; // @[Switch.scala 30:36:@4547.4]
  wire  _T_10165; // @[Switch.scala 30:53:@4549.4]
  wire  valid_28_1; // @[Switch.scala 30:36:@4550.4]
  wire  _T_10168; // @[Switch.scala 30:53:@4552.4]
  wire  valid_28_2; // @[Switch.scala 30:36:@4553.4]
  wire  _T_10171; // @[Switch.scala 30:53:@4555.4]
  wire  valid_28_3; // @[Switch.scala 30:36:@4556.4]
  wire  _T_10174; // @[Switch.scala 30:53:@4558.4]
  wire  valid_28_4; // @[Switch.scala 30:36:@4559.4]
  wire  _T_10177; // @[Switch.scala 30:53:@4561.4]
  wire  valid_28_5; // @[Switch.scala 30:36:@4562.4]
  wire  _T_10180; // @[Switch.scala 30:53:@4564.4]
  wire  valid_28_6; // @[Switch.scala 30:36:@4565.4]
  wire  _T_10183; // @[Switch.scala 30:53:@4567.4]
  wire  valid_28_7; // @[Switch.scala 30:36:@4568.4]
  wire  _T_10186; // @[Switch.scala 30:53:@4570.4]
  wire  valid_28_8; // @[Switch.scala 30:36:@4571.4]
  wire  _T_10189; // @[Switch.scala 30:53:@4573.4]
  wire  valid_28_9; // @[Switch.scala 30:36:@4574.4]
  wire  _T_10192; // @[Switch.scala 30:53:@4576.4]
  wire  valid_28_10; // @[Switch.scala 30:36:@4577.4]
  wire  _T_10195; // @[Switch.scala 30:53:@4579.4]
  wire  valid_28_11; // @[Switch.scala 30:36:@4580.4]
  wire  _T_10198; // @[Switch.scala 30:53:@4582.4]
  wire  valid_28_12; // @[Switch.scala 30:36:@4583.4]
  wire  _T_10201; // @[Switch.scala 30:53:@4585.4]
  wire  valid_28_13; // @[Switch.scala 30:36:@4586.4]
  wire  _T_10204; // @[Switch.scala 30:53:@4588.4]
  wire  valid_28_14; // @[Switch.scala 30:36:@4589.4]
  wire  _T_10207; // @[Switch.scala 30:53:@4591.4]
  wire  valid_28_15; // @[Switch.scala 30:36:@4592.4]
  wire  _T_10210; // @[Switch.scala 30:53:@4594.4]
  wire  valid_28_16; // @[Switch.scala 30:36:@4595.4]
  wire  _T_10213; // @[Switch.scala 30:53:@4597.4]
  wire  valid_28_17; // @[Switch.scala 30:36:@4598.4]
  wire  _T_10216; // @[Switch.scala 30:53:@4600.4]
  wire  valid_28_18; // @[Switch.scala 30:36:@4601.4]
  wire  _T_10219; // @[Switch.scala 30:53:@4603.4]
  wire  valid_28_19; // @[Switch.scala 30:36:@4604.4]
  wire  _T_10222; // @[Switch.scala 30:53:@4606.4]
  wire  valid_28_20; // @[Switch.scala 30:36:@4607.4]
  wire  _T_10225; // @[Switch.scala 30:53:@4609.4]
  wire  valid_28_21; // @[Switch.scala 30:36:@4610.4]
  wire  _T_10228; // @[Switch.scala 30:53:@4612.4]
  wire  valid_28_22; // @[Switch.scala 30:36:@4613.4]
  wire  _T_10231; // @[Switch.scala 30:53:@4615.4]
  wire  valid_28_23; // @[Switch.scala 30:36:@4616.4]
  wire  _T_10234; // @[Switch.scala 30:53:@4618.4]
  wire  valid_28_24; // @[Switch.scala 30:36:@4619.4]
  wire  _T_10237; // @[Switch.scala 30:53:@4621.4]
  wire  valid_28_25; // @[Switch.scala 30:36:@4622.4]
  wire  _T_10240; // @[Switch.scala 30:53:@4624.4]
  wire  valid_28_26; // @[Switch.scala 30:36:@4625.4]
  wire  _T_10243; // @[Switch.scala 30:53:@4627.4]
  wire  valid_28_27; // @[Switch.scala 30:36:@4628.4]
  wire  _T_10246; // @[Switch.scala 30:53:@4630.4]
  wire  valid_28_28; // @[Switch.scala 30:36:@4631.4]
  wire  _T_10249; // @[Switch.scala 30:53:@4633.4]
  wire  valid_28_29; // @[Switch.scala 30:36:@4634.4]
  wire  _T_10252; // @[Switch.scala 30:53:@4636.4]
  wire  valid_28_30; // @[Switch.scala 30:36:@4637.4]
  wire  _T_10255; // @[Switch.scala 30:53:@4639.4]
  wire  valid_28_31; // @[Switch.scala 30:36:@4640.4]
  wire [4:0] _T_10289; // @[Mux.scala 31:69:@4642.4]
  wire [4:0] _T_10290; // @[Mux.scala 31:69:@4643.4]
  wire [4:0] _T_10291; // @[Mux.scala 31:69:@4644.4]
  wire [4:0] _T_10292; // @[Mux.scala 31:69:@4645.4]
  wire [4:0] _T_10293; // @[Mux.scala 31:69:@4646.4]
  wire [4:0] _T_10294; // @[Mux.scala 31:69:@4647.4]
  wire [4:0] _T_10295; // @[Mux.scala 31:69:@4648.4]
  wire [4:0] _T_10296; // @[Mux.scala 31:69:@4649.4]
  wire [4:0] _T_10297; // @[Mux.scala 31:69:@4650.4]
  wire [4:0] _T_10298; // @[Mux.scala 31:69:@4651.4]
  wire [4:0] _T_10299; // @[Mux.scala 31:69:@4652.4]
  wire [4:0] _T_10300; // @[Mux.scala 31:69:@4653.4]
  wire [4:0] _T_10301; // @[Mux.scala 31:69:@4654.4]
  wire [4:0] _T_10302; // @[Mux.scala 31:69:@4655.4]
  wire [4:0] _T_10303; // @[Mux.scala 31:69:@4656.4]
  wire [4:0] _T_10304; // @[Mux.scala 31:69:@4657.4]
  wire [4:0] _T_10305; // @[Mux.scala 31:69:@4658.4]
  wire [4:0] _T_10306; // @[Mux.scala 31:69:@4659.4]
  wire [4:0] _T_10307; // @[Mux.scala 31:69:@4660.4]
  wire [4:0] _T_10308; // @[Mux.scala 31:69:@4661.4]
  wire [4:0] _T_10309; // @[Mux.scala 31:69:@4662.4]
  wire [4:0] _T_10310; // @[Mux.scala 31:69:@4663.4]
  wire [4:0] _T_10311; // @[Mux.scala 31:69:@4664.4]
  wire [4:0] _T_10312; // @[Mux.scala 31:69:@4665.4]
  wire [4:0] _T_10313; // @[Mux.scala 31:69:@4666.4]
  wire [4:0] _T_10314; // @[Mux.scala 31:69:@4667.4]
  wire [4:0] _T_10315; // @[Mux.scala 31:69:@4668.4]
  wire [4:0] _T_10316; // @[Mux.scala 31:69:@4669.4]
  wire [4:0] _T_10317; // @[Mux.scala 31:69:@4670.4]
  wire [4:0] _T_10318; // @[Mux.scala 31:69:@4671.4]
  wire [4:0] select_28; // @[Mux.scala 31:69:@4672.4]
  wire [47:0] _GEN_897; // @[Switch.scala 33:19:@4674.4]
  wire [47:0] _GEN_898; // @[Switch.scala 33:19:@4674.4]
  wire [47:0] _GEN_899; // @[Switch.scala 33:19:@4674.4]
  wire [47:0] _GEN_900; // @[Switch.scala 33:19:@4674.4]
  wire [47:0] _GEN_901; // @[Switch.scala 33:19:@4674.4]
  wire [47:0] _GEN_902; // @[Switch.scala 33:19:@4674.4]
  wire [47:0] _GEN_903; // @[Switch.scala 33:19:@4674.4]
  wire [47:0] _GEN_904; // @[Switch.scala 33:19:@4674.4]
  wire [47:0] _GEN_905; // @[Switch.scala 33:19:@4674.4]
  wire [47:0] _GEN_906; // @[Switch.scala 33:19:@4674.4]
  wire [47:0] _GEN_907; // @[Switch.scala 33:19:@4674.4]
  wire [47:0] _GEN_908; // @[Switch.scala 33:19:@4674.4]
  wire [47:0] _GEN_909; // @[Switch.scala 33:19:@4674.4]
  wire [47:0] _GEN_910; // @[Switch.scala 33:19:@4674.4]
  wire [47:0] _GEN_911; // @[Switch.scala 33:19:@4674.4]
  wire [47:0] _GEN_912; // @[Switch.scala 33:19:@4674.4]
  wire [47:0] _GEN_913; // @[Switch.scala 33:19:@4674.4]
  wire [47:0] _GEN_914; // @[Switch.scala 33:19:@4674.4]
  wire [47:0] _GEN_915; // @[Switch.scala 33:19:@4674.4]
  wire [47:0] _GEN_916; // @[Switch.scala 33:19:@4674.4]
  wire [47:0] _GEN_917; // @[Switch.scala 33:19:@4674.4]
  wire [47:0] _GEN_918; // @[Switch.scala 33:19:@4674.4]
  wire [47:0] _GEN_919; // @[Switch.scala 33:19:@4674.4]
  wire [47:0] _GEN_920; // @[Switch.scala 33:19:@4674.4]
  wire [47:0] _GEN_921; // @[Switch.scala 33:19:@4674.4]
  wire [47:0] _GEN_922; // @[Switch.scala 33:19:@4674.4]
  wire [47:0] _GEN_923; // @[Switch.scala 33:19:@4674.4]
  wire [47:0] _GEN_924; // @[Switch.scala 33:19:@4674.4]
  wire [47:0] _GEN_925; // @[Switch.scala 33:19:@4674.4]
  wire [47:0] _GEN_926; // @[Switch.scala 33:19:@4674.4]
  wire [7:0] _T_10327; // @[Switch.scala 34:32:@4681.4]
  wire [15:0] _T_10335; // @[Switch.scala 34:32:@4689.4]
  wire [7:0] _T_10342; // @[Switch.scala 34:32:@4696.4]
  wire [31:0] _T_10351; // @[Switch.scala 34:32:@4705.4]
  wire  _T_10355; // @[Switch.scala 30:53:@4708.4]
  wire  valid_29_0; // @[Switch.scala 30:36:@4709.4]
  wire  _T_10358; // @[Switch.scala 30:53:@4711.4]
  wire  valid_29_1; // @[Switch.scala 30:36:@4712.4]
  wire  _T_10361; // @[Switch.scala 30:53:@4714.4]
  wire  valid_29_2; // @[Switch.scala 30:36:@4715.4]
  wire  _T_10364; // @[Switch.scala 30:53:@4717.4]
  wire  valid_29_3; // @[Switch.scala 30:36:@4718.4]
  wire  _T_10367; // @[Switch.scala 30:53:@4720.4]
  wire  valid_29_4; // @[Switch.scala 30:36:@4721.4]
  wire  _T_10370; // @[Switch.scala 30:53:@4723.4]
  wire  valid_29_5; // @[Switch.scala 30:36:@4724.4]
  wire  _T_10373; // @[Switch.scala 30:53:@4726.4]
  wire  valid_29_6; // @[Switch.scala 30:36:@4727.4]
  wire  _T_10376; // @[Switch.scala 30:53:@4729.4]
  wire  valid_29_7; // @[Switch.scala 30:36:@4730.4]
  wire  _T_10379; // @[Switch.scala 30:53:@4732.4]
  wire  valid_29_8; // @[Switch.scala 30:36:@4733.4]
  wire  _T_10382; // @[Switch.scala 30:53:@4735.4]
  wire  valid_29_9; // @[Switch.scala 30:36:@4736.4]
  wire  _T_10385; // @[Switch.scala 30:53:@4738.4]
  wire  valid_29_10; // @[Switch.scala 30:36:@4739.4]
  wire  _T_10388; // @[Switch.scala 30:53:@4741.4]
  wire  valid_29_11; // @[Switch.scala 30:36:@4742.4]
  wire  _T_10391; // @[Switch.scala 30:53:@4744.4]
  wire  valid_29_12; // @[Switch.scala 30:36:@4745.4]
  wire  _T_10394; // @[Switch.scala 30:53:@4747.4]
  wire  valid_29_13; // @[Switch.scala 30:36:@4748.4]
  wire  _T_10397; // @[Switch.scala 30:53:@4750.4]
  wire  valid_29_14; // @[Switch.scala 30:36:@4751.4]
  wire  _T_10400; // @[Switch.scala 30:53:@4753.4]
  wire  valid_29_15; // @[Switch.scala 30:36:@4754.4]
  wire  _T_10403; // @[Switch.scala 30:53:@4756.4]
  wire  valid_29_16; // @[Switch.scala 30:36:@4757.4]
  wire  _T_10406; // @[Switch.scala 30:53:@4759.4]
  wire  valid_29_17; // @[Switch.scala 30:36:@4760.4]
  wire  _T_10409; // @[Switch.scala 30:53:@4762.4]
  wire  valid_29_18; // @[Switch.scala 30:36:@4763.4]
  wire  _T_10412; // @[Switch.scala 30:53:@4765.4]
  wire  valid_29_19; // @[Switch.scala 30:36:@4766.4]
  wire  _T_10415; // @[Switch.scala 30:53:@4768.4]
  wire  valid_29_20; // @[Switch.scala 30:36:@4769.4]
  wire  _T_10418; // @[Switch.scala 30:53:@4771.4]
  wire  valid_29_21; // @[Switch.scala 30:36:@4772.4]
  wire  _T_10421; // @[Switch.scala 30:53:@4774.4]
  wire  valid_29_22; // @[Switch.scala 30:36:@4775.4]
  wire  _T_10424; // @[Switch.scala 30:53:@4777.4]
  wire  valid_29_23; // @[Switch.scala 30:36:@4778.4]
  wire  _T_10427; // @[Switch.scala 30:53:@4780.4]
  wire  valid_29_24; // @[Switch.scala 30:36:@4781.4]
  wire  _T_10430; // @[Switch.scala 30:53:@4783.4]
  wire  valid_29_25; // @[Switch.scala 30:36:@4784.4]
  wire  _T_10433; // @[Switch.scala 30:53:@4786.4]
  wire  valid_29_26; // @[Switch.scala 30:36:@4787.4]
  wire  _T_10436; // @[Switch.scala 30:53:@4789.4]
  wire  valid_29_27; // @[Switch.scala 30:36:@4790.4]
  wire  _T_10439; // @[Switch.scala 30:53:@4792.4]
  wire  valid_29_28; // @[Switch.scala 30:36:@4793.4]
  wire  _T_10442; // @[Switch.scala 30:53:@4795.4]
  wire  valid_29_29; // @[Switch.scala 30:36:@4796.4]
  wire  _T_10445; // @[Switch.scala 30:53:@4798.4]
  wire  valid_29_30; // @[Switch.scala 30:36:@4799.4]
  wire  _T_10448; // @[Switch.scala 30:53:@4801.4]
  wire  valid_29_31; // @[Switch.scala 30:36:@4802.4]
  wire [4:0] _T_10482; // @[Mux.scala 31:69:@4804.4]
  wire [4:0] _T_10483; // @[Mux.scala 31:69:@4805.4]
  wire [4:0] _T_10484; // @[Mux.scala 31:69:@4806.4]
  wire [4:0] _T_10485; // @[Mux.scala 31:69:@4807.4]
  wire [4:0] _T_10486; // @[Mux.scala 31:69:@4808.4]
  wire [4:0] _T_10487; // @[Mux.scala 31:69:@4809.4]
  wire [4:0] _T_10488; // @[Mux.scala 31:69:@4810.4]
  wire [4:0] _T_10489; // @[Mux.scala 31:69:@4811.4]
  wire [4:0] _T_10490; // @[Mux.scala 31:69:@4812.4]
  wire [4:0] _T_10491; // @[Mux.scala 31:69:@4813.4]
  wire [4:0] _T_10492; // @[Mux.scala 31:69:@4814.4]
  wire [4:0] _T_10493; // @[Mux.scala 31:69:@4815.4]
  wire [4:0] _T_10494; // @[Mux.scala 31:69:@4816.4]
  wire [4:0] _T_10495; // @[Mux.scala 31:69:@4817.4]
  wire [4:0] _T_10496; // @[Mux.scala 31:69:@4818.4]
  wire [4:0] _T_10497; // @[Mux.scala 31:69:@4819.4]
  wire [4:0] _T_10498; // @[Mux.scala 31:69:@4820.4]
  wire [4:0] _T_10499; // @[Mux.scala 31:69:@4821.4]
  wire [4:0] _T_10500; // @[Mux.scala 31:69:@4822.4]
  wire [4:0] _T_10501; // @[Mux.scala 31:69:@4823.4]
  wire [4:0] _T_10502; // @[Mux.scala 31:69:@4824.4]
  wire [4:0] _T_10503; // @[Mux.scala 31:69:@4825.4]
  wire [4:0] _T_10504; // @[Mux.scala 31:69:@4826.4]
  wire [4:0] _T_10505; // @[Mux.scala 31:69:@4827.4]
  wire [4:0] _T_10506; // @[Mux.scala 31:69:@4828.4]
  wire [4:0] _T_10507; // @[Mux.scala 31:69:@4829.4]
  wire [4:0] _T_10508; // @[Mux.scala 31:69:@4830.4]
  wire [4:0] _T_10509; // @[Mux.scala 31:69:@4831.4]
  wire [4:0] _T_10510; // @[Mux.scala 31:69:@4832.4]
  wire [4:0] _T_10511; // @[Mux.scala 31:69:@4833.4]
  wire [4:0] select_29; // @[Mux.scala 31:69:@4834.4]
  wire [47:0] _GEN_929; // @[Switch.scala 33:19:@4836.4]
  wire [47:0] _GEN_930; // @[Switch.scala 33:19:@4836.4]
  wire [47:0] _GEN_931; // @[Switch.scala 33:19:@4836.4]
  wire [47:0] _GEN_932; // @[Switch.scala 33:19:@4836.4]
  wire [47:0] _GEN_933; // @[Switch.scala 33:19:@4836.4]
  wire [47:0] _GEN_934; // @[Switch.scala 33:19:@4836.4]
  wire [47:0] _GEN_935; // @[Switch.scala 33:19:@4836.4]
  wire [47:0] _GEN_936; // @[Switch.scala 33:19:@4836.4]
  wire [47:0] _GEN_937; // @[Switch.scala 33:19:@4836.4]
  wire [47:0] _GEN_938; // @[Switch.scala 33:19:@4836.4]
  wire [47:0] _GEN_939; // @[Switch.scala 33:19:@4836.4]
  wire [47:0] _GEN_940; // @[Switch.scala 33:19:@4836.4]
  wire [47:0] _GEN_941; // @[Switch.scala 33:19:@4836.4]
  wire [47:0] _GEN_942; // @[Switch.scala 33:19:@4836.4]
  wire [47:0] _GEN_943; // @[Switch.scala 33:19:@4836.4]
  wire [47:0] _GEN_944; // @[Switch.scala 33:19:@4836.4]
  wire [47:0] _GEN_945; // @[Switch.scala 33:19:@4836.4]
  wire [47:0] _GEN_946; // @[Switch.scala 33:19:@4836.4]
  wire [47:0] _GEN_947; // @[Switch.scala 33:19:@4836.4]
  wire [47:0] _GEN_948; // @[Switch.scala 33:19:@4836.4]
  wire [47:0] _GEN_949; // @[Switch.scala 33:19:@4836.4]
  wire [47:0] _GEN_950; // @[Switch.scala 33:19:@4836.4]
  wire [47:0] _GEN_951; // @[Switch.scala 33:19:@4836.4]
  wire [47:0] _GEN_952; // @[Switch.scala 33:19:@4836.4]
  wire [47:0] _GEN_953; // @[Switch.scala 33:19:@4836.4]
  wire [47:0] _GEN_954; // @[Switch.scala 33:19:@4836.4]
  wire [47:0] _GEN_955; // @[Switch.scala 33:19:@4836.4]
  wire [47:0] _GEN_956; // @[Switch.scala 33:19:@4836.4]
  wire [47:0] _GEN_957; // @[Switch.scala 33:19:@4836.4]
  wire [47:0] _GEN_958; // @[Switch.scala 33:19:@4836.4]
  wire [7:0] _T_10520; // @[Switch.scala 34:32:@4843.4]
  wire [15:0] _T_10528; // @[Switch.scala 34:32:@4851.4]
  wire [7:0] _T_10535; // @[Switch.scala 34:32:@4858.4]
  wire [31:0] _T_10544; // @[Switch.scala 34:32:@4867.4]
  wire  _T_10548; // @[Switch.scala 30:53:@4870.4]
  wire  valid_30_0; // @[Switch.scala 30:36:@4871.4]
  wire  _T_10551; // @[Switch.scala 30:53:@4873.4]
  wire  valid_30_1; // @[Switch.scala 30:36:@4874.4]
  wire  _T_10554; // @[Switch.scala 30:53:@4876.4]
  wire  valid_30_2; // @[Switch.scala 30:36:@4877.4]
  wire  _T_10557; // @[Switch.scala 30:53:@4879.4]
  wire  valid_30_3; // @[Switch.scala 30:36:@4880.4]
  wire  _T_10560; // @[Switch.scala 30:53:@4882.4]
  wire  valid_30_4; // @[Switch.scala 30:36:@4883.4]
  wire  _T_10563; // @[Switch.scala 30:53:@4885.4]
  wire  valid_30_5; // @[Switch.scala 30:36:@4886.4]
  wire  _T_10566; // @[Switch.scala 30:53:@4888.4]
  wire  valid_30_6; // @[Switch.scala 30:36:@4889.4]
  wire  _T_10569; // @[Switch.scala 30:53:@4891.4]
  wire  valid_30_7; // @[Switch.scala 30:36:@4892.4]
  wire  _T_10572; // @[Switch.scala 30:53:@4894.4]
  wire  valid_30_8; // @[Switch.scala 30:36:@4895.4]
  wire  _T_10575; // @[Switch.scala 30:53:@4897.4]
  wire  valid_30_9; // @[Switch.scala 30:36:@4898.4]
  wire  _T_10578; // @[Switch.scala 30:53:@4900.4]
  wire  valid_30_10; // @[Switch.scala 30:36:@4901.4]
  wire  _T_10581; // @[Switch.scala 30:53:@4903.4]
  wire  valid_30_11; // @[Switch.scala 30:36:@4904.4]
  wire  _T_10584; // @[Switch.scala 30:53:@4906.4]
  wire  valid_30_12; // @[Switch.scala 30:36:@4907.4]
  wire  _T_10587; // @[Switch.scala 30:53:@4909.4]
  wire  valid_30_13; // @[Switch.scala 30:36:@4910.4]
  wire  _T_10590; // @[Switch.scala 30:53:@4912.4]
  wire  valid_30_14; // @[Switch.scala 30:36:@4913.4]
  wire  _T_10593; // @[Switch.scala 30:53:@4915.4]
  wire  valid_30_15; // @[Switch.scala 30:36:@4916.4]
  wire  _T_10596; // @[Switch.scala 30:53:@4918.4]
  wire  valid_30_16; // @[Switch.scala 30:36:@4919.4]
  wire  _T_10599; // @[Switch.scala 30:53:@4921.4]
  wire  valid_30_17; // @[Switch.scala 30:36:@4922.4]
  wire  _T_10602; // @[Switch.scala 30:53:@4924.4]
  wire  valid_30_18; // @[Switch.scala 30:36:@4925.4]
  wire  _T_10605; // @[Switch.scala 30:53:@4927.4]
  wire  valid_30_19; // @[Switch.scala 30:36:@4928.4]
  wire  _T_10608; // @[Switch.scala 30:53:@4930.4]
  wire  valid_30_20; // @[Switch.scala 30:36:@4931.4]
  wire  _T_10611; // @[Switch.scala 30:53:@4933.4]
  wire  valid_30_21; // @[Switch.scala 30:36:@4934.4]
  wire  _T_10614; // @[Switch.scala 30:53:@4936.4]
  wire  valid_30_22; // @[Switch.scala 30:36:@4937.4]
  wire  _T_10617; // @[Switch.scala 30:53:@4939.4]
  wire  valid_30_23; // @[Switch.scala 30:36:@4940.4]
  wire  _T_10620; // @[Switch.scala 30:53:@4942.4]
  wire  valid_30_24; // @[Switch.scala 30:36:@4943.4]
  wire  _T_10623; // @[Switch.scala 30:53:@4945.4]
  wire  valid_30_25; // @[Switch.scala 30:36:@4946.4]
  wire  _T_10626; // @[Switch.scala 30:53:@4948.4]
  wire  valid_30_26; // @[Switch.scala 30:36:@4949.4]
  wire  _T_10629; // @[Switch.scala 30:53:@4951.4]
  wire  valid_30_27; // @[Switch.scala 30:36:@4952.4]
  wire  _T_10632; // @[Switch.scala 30:53:@4954.4]
  wire  valid_30_28; // @[Switch.scala 30:36:@4955.4]
  wire  _T_10635; // @[Switch.scala 30:53:@4957.4]
  wire  valid_30_29; // @[Switch.scala 30:36:@4958.4]
  wire  _T_10638; // @[Switch.scala 30:53:@4960.4]
  wire  valid_30_30; // @[Switch.scala 30:36:@4961.4]
  wire  _T_10641; // @[Switch.scala 30:53:@4963.4]
  wire  valid_30_31; // @[Switch.scala 30:36:@4964.4]
  wire [4:0] _T_10675; // @[Mux.scala 31:69:@4966.4]
  wire [4:0] _T_10676; // @[Mux.scala 31:69:@4967.4]
  wire [4:0] _T_10677; // @[Mux.scala 31:69:@4968.4]
  wire [4:0] _T_10678; // @[Mux.scala 31:69:@4969.4]
  wire [4:0] _T_10679; // @[Mux.scala 31:69:@4970.4]
  wire [4:0] _T_10680; // @[Mux.scala 31:69:@4971.4]
  wire [4:0] _T_10681; // @[Mux.scala 31:69:@4972.4]
  wire [4:0] _T_10682; // @[Mux.scala 31:69:@4973.4]
  wire [4:0] _T_10683; // @[Mux.scala 31:69:@4974.4]
  wire [4:0] _T_10684; // @[Mux.scala 31:69:@4975.4]
  wire [4:0] _T_10685; // @[Mux.scala 31:69:@4976.4]
  wire [4:0] _T_10686; // @[Mux.scala 31:69:@4977.4]
  wire [4:0] _T_10687; // @[Mux.scala 31:69:@4978.4]
  wire [4:0] _T_10688; // @[Mux.scala 31:69:@4979.4]
  wire [4:0] _T_10689; // @[Mux.scala 31:69:@4980.4]
  wire [4:0] _T_10690; // @[Mux.scala 31:69:@4981.4]
  wire [4:0] _T_10691; // @[Mux.scala 31:69:@4982.4]
  wire [4:0] _T_10692; // @[Mux.scala 31:69:@4983.4]
  wire [4:0] _T_10693; // @[Mux.scala 31:69:@4984.4]
  wire [4:0] _T_10694; // @[Mux.scala 31:69:@4985.4]
  wire [4:0] _T_10695; // @[Mux.scala 31:69:@4986.4]
  wire [4:0] _T_10696; // @[Mux.scala 31:69:@4987.4]
  wire [4:0] _T_10697; // @[Mux.scala 31:69:@4988.4]
  wire [4:0] _T_10698; // @[Mux.scala 31:69:@4989.4]
  wire [4:0] _T_10699; // @[Mux.scala 31:69:@4990.4]
  wire [4:0] _T_10700; // @[Mux.scala 31:69:@4991.4]
  wire [4:0] _T_10701; // @[Mux.scala 31:69:@4992.4]
  wire [4:0] _T_10702; // @[Mux.scala 31:69:@4993.4]
  wire [4:0] _T_10703; // @[Mux.scala 31:69:@4994.4]
  wire [4:0] _T_10704; // @[Mux.scala 31:69:@4995.4]
  wire [4:0] select_30; // @[Mux.scala 31:69:@4996.4]
  wire [47:0] _GEN_961; // @[Switch.scala 33:19:@4998.4]
  wire [47:0] _GEN_962; // @[Switch.scala 33:19:@4998.4]
  wire [47:0] _GEN_963; // @[Switch.scala 33:19:@4998.4]
  wire [47:0] _GEN_964; // @[Switch.scala 33:19:@4998.4]
  wire [47:0] _GEN_965; // @[Switch.scala 33:19:@4998.4]
  wire [47:0] _GEN_966; // @[Switch.scala 33:19:@4998.4]
  wire [47:0] _GEN_967; // @[Switch.scala 33:19:@4998.4]
  wire [47:0] _GEN_968; // @[Switch.scala 33:19:@4998.4]
  wire [47:0] _GEN_969; // @[Switch.scala 33:19:@4998.4]
  wire [47:0] _GEN_970; // @[Switch.scala 33:19:@4998.4]
  wire [47:0] _GEN_971; // @[Switch.scala 33:19:@4998.4]
  wire [47:0] _GEN_972; // @[Switch.scala 33:19:@4998.4]
  wire [47:0] _GEN_973; // @[Switch.scala 33:19:@4998.4]
  wire [47:0] _GEN_974; // @[Switch.scala 33:19:@4998.4]
  wire [47:0] _GEN_975; // @[Switch.scala 33:19:@4998.4]
  wire [47:0] _GEN_976; // @[Switch.scala 33:19:@4998.4]
  wire [47:0] _GEN_977; // @[Switch.scala 33:19:@4998.4]
  wire [47:0] _GEN_978; // @[Switch.scala 33:19:@4998.4]
  wire [47:0] _GEN_979; // @[Switch.scala 33:19:@4998.4]
  wire [47:0] _GEN_980; // @[Switch.scala 33:19:@4998.4]
  wire [47:0] _GEN_981; // @[Switch.scala 33:19:@4998.4]
  wire [47:0] _GEN_982; // @[Switch.scala 33:19:@4998.4]
  wire [47:0] _GEN_983; // @[Switch.scala 33:19:@4998.4]
  wire [47:0] _GEN_984; // @[Switch.scala 33:19:@4998.4]
  wire [47:0] _GEN_985; // @[Switch.scala 33:19:@4998.4]
  wire [47:0] _GEN_986; // @[Switch.scala 33:19:@4998.4]
  wire [47:0] _GEN_987; // @[Switch.scala 33:19:@4998.4]
  wire [47:0] _GEN_988; // @[Switch.scala 33:19:@4998.4]
  wire [47:0] _GEN_989; // @[Switch.scala 33:19:@4998.4]
  wire [47:0] _GEN_990; // @[Switch.scala 33:19:@4998.4]
  wire [7:0] _T_10713; // @[Switch.scala 34:32:@5005.4]
  wire [15:0] _T_10721; // @[Switch.scala 34:32:@5013.4]
  wire [7:0] _T_10728; // @[Switch.scala 34:32:@5020.4]
  wire [31:0] _T_10737; // @[Switch.scala 34:32:@5029.4]
  wire  _T_10741; // @[Switch.scala 30:53:@5032.4]
  wire  valid_31_0; // @[Switch.scala 30:36:@5033.4]
  wire  _T_10744; // @[Switch.scala 30:53:@5035.4]
  wire  valid_31_1; // @[Switch.scala 30:36:@5036.4]
  wire  _T_10747; // @[Switch.scala 30:53:@5038.4]
  wire  valid_31_2; // @[Switch.scala 30:36:@5039.4]
  wire  _T_10750; // @[Switch.scala 30:53:@5041.4]
  wire  valid_31_3; // @[Switch.scala 30:36:@5042.4]
  wire  _T_10753; // @[Switch.scala 30:53:@5044.4]
  wire  valid_31_4; // @[Switch.scala 30:36:@5045.4]
  wire  _T_10756; // @[Switch.scala 30:53:@5047.4]
  wire  valid_31_5; // @[Switch.scala 30:36:@5048.4]
  wire  _T_10759; // @[Switch.scala 30:53:@5050.4]
  wire  valid_31_6; // @[Switch.scala 30:36:@5051.4]
  wire  _T_10762; // @[Switch.scala 30:53:@5053.4]
  wire  valid_31_7; // @[Switch.scala 30:36:@5054.4]
  wire  _T_10765; // @[Switch.scala 30:53:@5056.4]
  wire  valid_31_8; // @[Switch.scala 30:36:@5057.4]
  wire  _T_10768; // @[Switch.scala 30:53:@5059.4]
  wire  valid_31_9; // @[Switch.scala 30:36:@5060.4]
  wire  _T_10771; // @[Switch.scala 30:53:@5062.4]
  wire  valid_31_10; // @[Switch.scala 30:36:@5063.4]
  wire  _T_10774; // @[Switch.scala 30:53:@5065.4]
  wire  valid_31_11; // @[Switch.scala 30:36:@5066.4]
  wire  _T_10777; // @[Switch.scala 30:53:@5068.4]
  wire  valid_31_12; // @[Switch.scala 30:36:@5069.4]
  wire  _T_10780; // @[Switch.scala 30:53:@5071.4]
  wire  valid_31_13; // @[Switch.scala 30:36:@5072.4]
  wire  _T_10783; // @[Switch.scala 30:53:@5074.4]
  wire  valid_31_14; // @[Switch.scala 30:36:@5075.4]
  wire  _T_10786; // @[Switch.scala 30:53:@5077.4]
  wire  valid_31_15; // @[Switch.scala 30:36:@5078.4]
  wire  _T_10789; // @[Switch.scala 30:53:@5080.4]
  wire  valid_31_16; // @[Switch.scala 30:36:@5081.4]
  wire  _T_10792; // @[Switch.scala 30:53:@5083.4]
  wire  valid_31_17; // @[Switch.scala 30:36:@5084.4]
  wire  _T_10795; // @[Switch.scala 30:53:@5086.4]
  wire  valid_31_18; // @[Switch.scala 30:36:@5087.4]
  wire  _T_10798; // @[Switch.scala 30:53:@5089.4]
  wire  valid_31_19; // @[Switch.scala 30:36:@5090.4]
  wire  _T_10801; // @[Switch.scala 30:53:@5092.4]
  wire  valid_31_20; // @[Switch.scala 30:36:@5093.4]
  wire  _T_10804; // @[Switch.scala 30:53:@5095.4]
  wire  valid_31_21; // @[Switch.scala 30:36:@5096.4]
  wire  _T_10807; // @[Switch.scala 30:53:@5098.4]
  wire  valid_31_22; // @[Switch.scala 30:36:@5099.4]
  wire  _T_10810; // @[Switch.scala 30:53:@5101.4]
  wire  valid_31_23; // @[Switch.scala 30:36:@5102.4]
  wire  _T_10813; // @[Switch.scala 30:53:@5104.4]
  wire  valid_31_24; // @[Switch.scala 30:36:@5105.4]
  wire  _T_10816; // @[Switch.scala 30:53:@5107.4]
  wire  valid_31_25; // @[Switch.scala 30:36:@5108.4]
  wire  _T_10819; // @[Switch.scala 30:53:@5110.4]
  wire  valid_31_26; // @[Switch.scala 30:36:@5111.4]
  wire  _T_10822; // @[Switch.scala 30:53:@5113.4]
  wire  valid_31_27; // @[Switch.scala 30:36:@5114.4]
  wire  _T_10825; // @[Switch.scala 30:53:@5116.4]
  wire  valid_31_28; // @[Switch.scala 30:36:@5117.4]
  wire  _T_10828; // @[Switch.scala 30:53:@5119.4]
  wire  valid_31_29; // @[Switch.scala 30:36:@5120.4]
  wire  _T_10831; // @[Switch.scala 30:53:@5122.4]
  wire  valid_31_30; // @[Switch.scala 30:36:@5123.4]
  wire  _T_10834; // @[Switch.scala 30:53:@5125.4]
  wire  valid_31_31; // @[Switch.scala 30:36:@5126.4]
  wire [4:0] _T_10868; // @[Mux.scala 31:69:@5128.4]
  wire [4:0] _T_10869; // @[Mux.scala 31:69:@5129.4]
  wire [4:0] _T_10870; // @[Mux.scala 31:69:@5130.4]
  wire [4:0] _T_10871; // @[Mux.scala 31:69:@5131.4]
  wire [4:0] _T_10872; // @[Mux.scala 31:69:@5132.4]
  wire [4:0] _T_10873; // @[Mux.scala 31:69:@5133.4]
  wire [4:0] _T_10874; // @[Mux.scala 31:69:@5134.4]
  wire [4:0] _T_10875; // @[Mux.scala 31:69:@5135.4]
  wire [4:0] _T_10876; // @[Mux.scala 31:69:@5136.4]
  wire [4:0] _T_10877; // @[Mux.scala 31:69:@5137.4]
  wire [4:0] _T_10878; // @[Mux.scala 31:69:@5138.4]
  wire [4:0] _T_10879; // @[Mux.scala 31:69:@5139.4]
  wire [4:0] _T_10880; // @[Mux.scala 31:69:@5140.4]
  wire [4:0] _T_10881; // @[Mux.scala 31:69:@5141.4]
  wire [4:0] _T_10882; // @[Mux.scala 31:69:@5142.4]
  wire [4:0] _T_10883; // @[Mux.scala 31:69:@5143.4]
  wire [4:0] _T_10884; // @[Mux.scala 31:69:@5144.4]
  wire [4:0] _T_10885; // @[Mux.scala 31:69:@5145.4]
  wire [4:0] _T_10886; // @[Mux.scala 31:69:@5146.4]
  wire [4:0] _T_10887; // @[Mux.scala 31:69:@5147.4]
  wire [4:0] _T_10888; // @[Mux.scala 31:69:@5148.4]
  wire [4:0] _T_10889; // @[Mux.scala 31:69:@5149.4]
  wire [4:0] _T_10890; // @[Mux.scala 31:69:@5150.4]
  wire [4:0] _T_10891; // @[Mux.scala 31:69:@5151.4]
  wire [4:0] _T_10892; // @[Mux.scala 31:69:@5152.4]
  wire [4:0] _T_10893; // @[Mux.scala 31:69:@5153.4]
  wire [4:0] _T_10894; // @[Mux.scala 31:69:@5154.4]
  wire [4:0] _T_10895; // @[Mux.scala 31:69:@5155.4]
  wire [4:0] _T_10896; // @[Mux.scala 31:69:@5156.4]
  wire [4:0] _T_10897; // @[Mux.scala 31:69:@5157.4]
  wire [4:0] select_31; // @[Mux.scala 31:69:@5158.4]
  wire [47:0] _GEN_993; // @[Switch.scala 33:19:@5160.4]
  wire [47:0] _GEN_994; // @[Switch.scala 33:19:@5160.4]
  wire [47:0] _GEN_995; // @[Switch.scala 33:19:@5160.4]
  wire [47:0] _GEN_996; // @[Switch.scala 33:19:@5160.4]
  wire [47:0] _GEN_997; // @[Switch.scala 33:19:@5160.4]
  wire [47:0] _GEN_998; // @[Switch.scala 33:19:@5160.4]
  wire [47:0] _GEN_999; // @[Switch.scala 33:19:@5160.4]
  wire [47:0] _GEN_1000; // @[Switch.scala 33:19:@5160.4]
  wire [47:0] _GEN_1001; // @[Switch.scala 33:19:@5160.4]
  wire [47:0] _GEN_1002; // @[Switch.scala 33:19:@5160.4]
  wire [47:0] _GEN_1003; // @[Switch.scala 33:19:@5160.4]
  wire [47:0] _GEN_1004; // @[Switch.scala 33:19:@5160.4]
  wire [47:0] _GEN_1005; // @[Switch.scala 33:19:@5160.4]
  wire [47:0] _GEN_1006; // @[Switch.scala 33:19:@5160.4]
  wire [47:0] _GEN_1007; // @[Switch.scala 33:19:@5160.4]
  wire [47:0] _GEN_1008; // @[Switch.scala 33:19:@5160.4]
  wire [47:0] _GEN_1009; // @[Switch.scala 33:19:@5160.4]
  wire [47:0] _GEN_1010; // @[Switch.scala 33:19:@5160.4]
  wire [47:0] _GEN_1011; // @[Switch.scala 33:19:@5160.4]
  wire [47:0] _GEN_1012; // @[Switch.scala 33:19:@5160.4]
  wire [47:0] _GEN_1013; // @[Switch.scala 33:19:@5160.4]
  wire [47:0] _GEN_1014; // @[Switch.scala 33:19:@5160.4]
  wire [47:0] _GEN_1015; // @[Switch.scala 33:19:@5160.4]
  wire [47:0] _GEN_1016; // @[Switch.scala 33:19:@5160.4]
  wire [47:0] _GEN_1017; // @[Switch.scala 33:19:@5160.4]
  wire [47:0] _GEN_1018; // @[Switch.scala 33:19:@5160.4]
  wire [47:0] _GEN_1019; // @[Switch.scala 33:19:@5160.4]
  wire [47:0] _GEN_1020; // @[Switch.scala 33:19:@5160.4]
  wire [47:0] _GEN_1021; // @[Switch.scala 33:19:@5160.4]
  wire [47:0] _GEN_1022; // @[Switch.scala 33:19:@5160.4]
  wire [7:0] _T_10906; // @[Switch.scala 34:32:@5167.4]
  wire [15:0] _T_10914; // @[Switch.scala 34:32:@5175.4]
  wire [7:0] _T_10921; // @[Switch.scala 34:32:@5182.4]
  wire [31:0] _T_10930; // @[Switch.scala 34:32:@5191.4]
  wire  _T_15428; // @[Switch.scala 41:52:@5195.4]
  wire  output_0_0; // @[Switch.scala 41:38:@5196.4]
  wire  _T_15431; // @[Switch.scala 41:52:@5198.4]
  wire  output_0_1; // @[Switch.scala 41:38:@5199.4]
  wire  _T_15434; // @[Switch.scala 41:52:@5201.4]
  wire  output_0_2; // @[Switch.scala 41:38:@5202.4]
  wire  _T_15437; // @[Switch.scala 41:52:@5204.4]
  wire  output_0_3; // @[Switch.scala 41:38:@5205.4]
  wire  _T_15440; // @[Switch.scala 41:52:@5207.4]
  wire  output_0_4; // @[Switch.scala 41:38:@5208.4]
  wire  _T_15443; // @[Switch.scala 41:52:@5210.4]
  wire  output_0_5; // @[Switch.scala 41:38:@5211.4]
  wire  _T_15446; // @[Switch.scala 41:52:@5213.4]
  wire  output_0_6; // @[Switch.scala 41:38:@5214.4]
  wire  _T_15449; // @[Switch.scala 41:52:@5216.4]
  wire  output_0_7; // @[Switch.scala 41:38:@5217.4]
  wire  _T_15452; // @[Switch.scala 41:52:@5219.4]
  wire  output_0_8; // @[Switch.scala 41:38:@5220.4]
  wire  _T_15455; // @[Switch.scala 41:52:@5222.4]
  wire  output_0_9; // @[Switch.scala 41:38:@5223.4]
  wire  _T_15458; // @[Switch.scala 41:52:@5225.4]
  wire  output_0_10; // @[Switch.scala 41:38:@5226.4]
  wire  _T_15461; // @[Switch.scala 41:52:@5228.4]
  wire  output_0_11; // @[Switch.scala 41:38:@5229.4]
  wire  _T_15464; // @[Switch.scala 41:52:@5231.4]
  wire  output_0_12; // @[Switch.scala 41:38:@5232.4]
  wire  _T_15467; // @[Switch.scala 41:52:@5234.4]
  wire  output_0_13; // @[Switch.scala 41:38:@5235.4]
  wire  _T_15470; // @[Switch.scala 41:52:@5237.4]
  wire  output_0_14; // @[Switch.scala 41:38:@5238.4]
  wire  _T_15473; // @[Switch.scala 41:52:@5240.4]
  wire  output_0_15; // @[Switch.scala 41:38:@5241.4]
  wire  _T_15476; // @[Switch.scala 41:52:@5243.4]
  wire  output_0_16; // @[Switch.scala 41:38:@5244.4]
  wire  _T_15479; // @[Switch.scala 41:52:@5246.4]
  wire  output_0_17; // @[Switch.scala 41:38:@5247.4]
  wire  _T_15482; // @[Switch.scala 41:52:@5249.4]
  wire  output_0_18; // @[Switch.scala 41:38:@5250.4]
  wire  _T_15485; // @[Switch.scala 41:52:@5252.4]
  wire  output_0_19; // @[Switch.scala 41:38:@5253.4]
  wire  _T_15488; // @[Switch.scala 41:52:@5255.4]
  wire  output_0_20; // @[Switch.scala 41:38:@5256.4]
  wire  _T_15491; // @[Switch.scala 41:52:@5258.4]
  wire  output_0_21; // @[Switch.scala 41:38:@5259.4]
  wire  _T_15494; // @[Switch.scala 41:52:@5261.4]
  wire  output_0_22; // @[Switch.scala 41:38:@5262.4]
  wire  _T_15497; // @[Switch.scala 41:52:@5264.4]
  wire  output_0_23; // @[Switch.scala 41:38:@5265.4]
  wire  _T_15500; // @[Switch.scala 41:52:@5267.4]
  wire  output_0_24; // @[Switch.scala 41:38:@5268.4]
  wire  _T_15503; // @[Switch.scala 41:52:@5270.4]
  wire  output_0_25; // @[Switch.scala 41:38:@5271.4]
  wire  _T_15506; // @[Switch.scala 41:52:@5273.4]
  wire  output_0_26; // @[Switch.scala 41:38:@5274.4]
  wire  _T_15509; // @[Switch.scala 41:52:@5276.4]
  wire  output_0_27; // @[Switch.scala 41:38:@5277.4]
  wire  _T_15512; // @[Switch.scala 41:52:@5279.4]
  wire  output_0_28; // @[Switch.scala 41:38:@5280.4]
  wire  _T_15515; // @[Switch.scala 41:52:@5282.4]
  wire  output_0_29; // @[Switch.scala 41:38:@5283.4]
  wire  _T_15518; // @[Switch.scala 41:52:@5285.4]
  wire  output_0_30; // @[Switch.scala 41:38:@5286.4]
  wire  _T_15521; // @[Switch.scala 41:52:@5288.4]
  wire  output_0_31; // @[Switch.scala 41:38:@5289.4]
  wire [7:0] _T_15529; // @[Switch.scala 43:31:@5297.4]
  wire [15:0] _T_15537; // @[Switch.scala 43:31:@5305.4]
  wire [7:0] _T_15544; // @[Switch.scala 43:31:@5312.4]
  wire [31:0] _T_15553; // @[Switch.scala 43:31:@5321.4]
  wire  _T_15557; // @[Switch.scala 41:52:@5324.4]
  wire  output_1_0; // @[Switch.scala 41:38:@5325.4]
  wire  _T_15560; // @[Switch.scala 41:52:@5327.4]
  wire  output_1_1; // @[Switch.scala 41:38:@5328.4]
  wire  _T_15563; // @[Switch.scala 41:52:@5330.4]
  wire  output_1_2; // @[Switch.scala 41:38:@5331.4]
  wire  _T_15566; // @[Switch.scala 41:52:@5333.4]
  wire  output_1_3; // @[Switch.scala 41:38:@5334.4]
  wire  _T_15569; // @[Switch.scala 41:52:@5336.4]
  wire  output_1_4; // @[Switch.scala 41:38:@5337.4]
  wire  _T_15572; // @[Switch.scala 41:52:@5339.4]
  wire  output_1_5; // @[Switch.scala 41:38:@5340.4]
  wire  _T_15575; // @[Switch.scala 41:52:@5342.4]
  wire  output_1_6; // @[Switch.scala 41:38:@5343.4]
  wire  _T_15578; // @[Switch.scala 41:52:@5345.4]
  wire  output_1_7; // @[Switch.scala 41:38:@5346.4]
  wire  _T_15581; // @[Switch.scala 41:52:@5348.4]
  wire  output_1_8; // @[Switch.scala 41:38:@5349.4]
  wire  _T_15584; // @[Switch.scala 41:52:@5351.4]
  wire  output_1_9; // @[Switch.scala 41:38:@5352.4]
  wire  _T_15587; // @[Switch.scala 41:52:@5354.4]
  wire  output_1_10; // @[Switch.scala 41:38:@5355.4]
  wire  _T_15590; // @[Switch.scala 41:52:@5357.4]
  wire  output_1_11; // @[Switch.scala 41:38:@5358.4]
  wire  _T_15593; // @[Switch.scala 41:52:@5360.4]
  wire  output_1_12; // @[Switch.scala 41:38:@5361.4]
  wire  _T_15596; // @[Switch.scala 41:52:@5363.4]
  wire  output_1_13; // @[Switch.scala 41:38:@5364.4]
  wire  _T_15599; // @[Switch.scala 41:52:@5366.4]
  wire  output_1_14; // @[Switch.scala 41:38:@5367.4]
  wire  _T_15602; // @[Switch.scala 41:52:@5369.4]
  wire  output_1_15; // @[Switch.scala 41:38:@5370.4]
  wire  _T_15605; // @[Switch.scala 41:52:@5372.4]
  wire  output_1_16; // @[Switch.scala 41:38:@5373.4]
  wire  _T_15608; // @[Switch.scala 41:52:@5375.4]
  wire  output_1_17; // @[Switch.scala 41:38:@5376.4]
  wire  _T_15611; // @[Switch.scala 41:52:@5378.4]
  wire  output_1_18; // @[Switch.scala 41:38:@5379.4]
  wire  _T_15614; // @[Switch.scala 41:52:@5381.4]
  wire  output_1_19; // @[Switch.scala 41:38:@5382.4]
  wire  _T_15617; // @[Switch.scala 41:52:@5384.4]
  wire  output_1_20; // @[Switch.scala 41:38:@5385.4]
  wire  _T_15620; // @[Switch.scala 41:52:@5387.4]
  wire  output_1_21; // @[Switch.scala 41:38:@5388.4]
  wire  _T_15623; // @[Switch.scala 41:52:@5390.4]
  wire  output_1_22; // @[Switch.scala 41:38:@5391.4]
  wire  _T_15626; // @[Switch.scala 41:52:@5393.4]
  wire  output_1_23; // @[Switch.scala 41:38:@5394.4]
  wire  _T_15629; // @[Switch.scala 41:52:@5396.4]
  wire  output_1_24; // @[Switch.scala 41:38:@5397.4]
  wire  _T_15632; // @[Switch.scala 41:52:@5399.4]
  wire  output_1_25; // @[Switch.scala 41:38:@5400.4]
  wire  _T_15635; // @[Switch.scala 41:52:@5402.4]
  wire  output_1_26; // @[Switch.scala 41:38:@5403.4]
  wire  _T_15638; // @[Switch.scala 41:52:@5405.4]
  wire  output_1_27; // @[Switch.scala 41:38:@5406.4]
  wire  _T_15641; // @[Switch.scala 41:52:@5408.4]
  wire  output_1_28; // @[Switch.scala 41:38:@5409.4]
  wire  _T_15644; // @[Switch.scala 41:52:@5411.4]
  wire  output_1_29; // @[Switch.scala 41:38:@5412.4]
  wire  _T_15647; // @[Switch.scala 41:52:@5414.4]
  wire  output_1_30; // @[Switch.scala 41:38:@5415.4]
  wire  _T_15650; // @[Switch.scala 41:52:@5417.4]
  wire  output_1_31; // @[Switch.scala 41:38:@5418.4]
  wire [7:0] _T_15658; // @[Switch.scala 43:31:@5426.4]
  wire [15:0] _T_15666; // @[Switch.scala 43:31:@5434.4]
  wire [7:0] _T_15673; // @[Switch.scala 43:31:@5441.4]
  wire [31:0] _T_15682; // @[Switch.scala 43:31:@5450.4]
  wire  _T_15686; // @[Switch.scala 41:52:@5453.4]
  wire  output_2_0; // @[Switch.scala 41:38:@5454.4]
  wire  _T_15689; // @[Switch.scala 41:52:@5456.4]
  wire  output_2_1; // @[Switch.scala 41:38:@5457.4]
  wire  _T_15692; // @[Switch.scala 41:52:@5459.4]
  wire  output_2_2; // @[Switch.scala 41:38:@5460.4]
  wire  _T_15695; // @[Switch.scala 41:52:@5462.4]
  wire  output_2_3; // @[Switch.scala 41:38:@5463.4]
  wire  _T_15698; // @[Switch.scala 41:52:@5465.4]
  wire  output_2_4; // @[Switch.scala 41:38:@5466.4]
  wire  _T_15701; // @[Switch.scala 41:52:@5468.4]
  wire  output_2_5; // @[Switch.scala 41:38:@5469.4]
  wire  _T_15704; // @[Switch.scala 41:52:@5471.4]
  wire  output_2_6; // @[Switch.scala 41:38:@5472.4]
  wire  _T_15707; // @[Switch.scala 41:52:@5474.4]
  wire  output_2_7; // @[Switch.scala 41:38:@5475.4]
  wire  _T_15710; // @[Switch.scala 41:52:@5477.4]
  wire  output_2_8; // @[Switch.scala 41:38:@5478.4]
  wire  _T_15713; // @[Switch.scala 41:52:@5480.4]
  wire  output_2_9; // @[Switch.scala 41:38:@5481.4]
  wire  _T_15716; // @[Switch.scala 41:52:@5483.4]
  wire  output_2_10; // @[Switch.scala 41:38:@5484.4]
  wire  _T_15719; // @[Switch.scala 41:52:@5486.4]
  wire  output_2_11; // @[Switch.scala 41:38:@5487.4]
  wire  _T_15722; // @[Switch.scala 41:52:@5489.4]
  wire  output_2_12; // @[Switch.scala 41:38:@5490.4]
  wire  _T_15725; // @[Switch.scala 41:52:@5492.4]
  wire  output_2_13; // @[Switch.scala 41:38:@5493.4]
  wire  _T_15728; // @[Switch.scala 41:52:@5495.4]
  wire  output_2_14; // @[Switch.scala 41:38:@5496.4]
  wire  _T_15731; // @[Switch.scala 41:52:@5498.4]
  wire  output_2_15; // @[Switch.scala 41:38:@5499.4]
  wire  _T_15734; // @[Switch.scala 41:52:@5501.4]
  wire  output_2_16; // @[Switch.scala 41:38:@5502.4]
  wire  _T_15737; // @[Switch.scala 41:52:@5504.4]
  wire  output_2_17; // @[Switch.scala 41:38:@5505.4]
  wire  _T_15740; // @[Switch.scala 41:52:@5507.4]
  wire  output_2_18; // @[Switch.scala 41:38:@5508.4]
  wire  _T_15743; // @[Switch.scala 41:52:@5510.4]
  wire  output_2_19; // @[Switch.scala 41:38:@5511.4]
  wire  _T_15746; // @[Switch.scala 41:52:@5513.4]
  wire  output_2_20; // @[Switch.scala 41:38:@5514.4]
  wire  _T_15749; // @[Switch.scala 41:52:@5516.4]
  wire  output_2_21; // @[Switch.scala 41:38:@5517.4]
  wire  _T_15752; // @[Switch.scala 41:52:@5519.4]
  wire  output_2_22; // @[Switch.scala 41:38:@5520.4]
  wire  _T_15755; // @[Switch.scala 41:52:@5522.4]
  wire  output_2_23; // @[Switch.scala 41:38:@5523.4]
  wire  _T_15758; // @[Switch.scala 41:52:@5525.4]
  wire  output_2_24; // @[Switch.scala 41:38:@5526.4]
  wire  _T_15761; // @[Switch.scala 41:52:@5528.4]
  wire  output_2_25; // @[Switch.scala 41:38:@5529.4]
  wire  _T_15764; // @[Switch.scala 41:52:@5531.4]
  wire  output_2_26; // @[Switch.scala 41:38:@5532.4]
  wire  _T_15767; // @[Switch.scala 41:52:@5534.4]
  wire  output_2_27; // @[Switch.scala 41:38:@5535.4]
  wire  _T_15770; // @[Switch.scala 41:52:@5537.4]
  wire  output_2_28; // @[Switch.scala 41:38:@5538.4]
  wire  _T_15773; // @[Switch.scala 41:52:@5540.4]
  wire  output_2_29; // @[Switch.scala 41:38:@5541.4]
  wire  _T_15776; // @[Switch.scala 41:52:@5543.4]
  wire  output_2_30; // @[Switch.scala 41:38:@5544.4]
  wire  _T_15779; // @[Switch.scala 41:52:@5546.4]
  wire  output_2_31; // @[Switch.scala 41:38:@5547.4]
  wire [7:0] _T_15787; // @[Switch.scala 43:31:@5555.4]
  wire [15:0] _T_15795; // @[Switch.scala 43:31:@5563.4]
  wire [7:0] _T_15802; // @[Switch.scala 43:31:@5570.4]
  wire [31:0] _T_15811; // @[Switch.scala 43:31:@5579.4]
  wire  _T_15815; // @[Switch.scala 41:52:@5582.4]
  wire  output_3_0; // @[Switch.scala 41:38:@5583.4]
  wire  _T_15818; // @[Switch.scala 41:52:@5585.4]
  wire  output_3_1; // @[Switch.scala 41:38:@5586.4]
  wire  _T_15821; // @[Switch.scala 41:52:@5588.4]
  wire  output_3_2; // @[Switch.scala 41:38:@5589.4]
  wire  _T_15824; // @[Switch.scala 41:52:@5591.4]
  wire  output_3_3; // @[Switch.scala 41:38:@5592.4]
  wire  _T_15827; // @[Switch.scala 41:52:@5594.4]
  wire  output_3_4; // @[Switch.scala 41:38:@5595.4]
  wire  _T_15830; // @[Switch.scala 41:52:@5597.4]
  wire  output_3_5; // @[Switch.scala 41:38:@5598.4]
  wire  _T_15833; // @[Switch.scala 41:52:@5600.4]
  wire  output_3_6; // @[Switch.scala 41:38:@5601.4]
  wire  _T_15836; // @[Switch.scala 41:52:@5603.4]
  wire  output_3_7; // @[Switch.scala 41:38:@5604.4]
  wire  _T_15839; // @[Switch.scala 41:52:@5606.4]
  wire  output_3_8; // @[Switch.scala 41:38:@5607.4]
  wire  _T_15842; // @[Switch.scala 41:52:@5609.4]
  wire  output_3_9; // @[Switch.scala 41:38:@5610.4]
  wire  _T_15845; // @[Switch.scala 41:52:@5612.4]
  wire  output_3_10; // @[Switch.scala 41:38:@5613.4]
  wire  _T_15848; // @[Switch.scala 41:52:@5615.4]
  wire  output_3_11; // @[Switch.scala 41:38:@5616.4]
  wire  _T_15851; // @[Switch.scala 41:52:@5618.4]
  wire  output_3_12; // @[Switch.scala 41:38:@5619.4]
  wire  _T_15854; // @[Switch.scala 41:52:@5621.4]
  wire  output_3_13; // @[Switch.scala 41:38:@5622.4]
  wire  _T_15857; // @[Switch.scala 41:52:@5624.4]
  wire  output_3_14; // @[Switch.scala 41:38:@5625.4]
  wire  _T_15860; // @[Switch.scala 41:52:@5627.4]
  wire  output_3_15; // @[Switch.scala 41:38:@5628.4]
  wire  _T_15863; // @[Switch.scala 41:52:@5630.4]
  wire  output_3_16; // @[Switch.scala 41:38:@5631.4]
  wire  _T_15866; // @[Switch.scala 41:52:@5633.4]
  wire  output_3_17; // @[Switch.scala 41:38:@5634.4]
  wire  _T_15869; // @[Switch.scala 41:52:@5636.4]
  wire  output_3_18; // @[Switch.scala 41:38:@5637.4]
  wire  _T_15872; // @[Switch.scala 41:52:@5639.4]
  wire  output_3_19; // @[Switch.scala 41:38:@5640.4]
  wire  _T_15875; // @[Switch.scala 41:52:@5642.4]
  wire  output_3_20; // @[Switch.scala 41:38:@5643.4]
  wire  _T_15878; // @[Switch.scala 41:52:@5645.4]
  wire  output_3_21; // @[Switch.scala 41:38:@5646.4]
  wire  _T_15881; // @[Switch.scala 41:52:@5648.4]
  wire  output_3_22; // @[Switch.scala 41:38:@5649.4]
  wire  _T_15884; // @[Switch.scala 41:52:@5651.4]
  wire  output_3_23; // @[Switch.scala 41:38:@5652.4]
  wire  _T_15887; // @[Switch.scala 41:52:@5654.4]
  wire  output_3_24; // @[Switch.scala 41:38:@5655.4]
  wire  _T_15890; // @[Switch.scala 41:52:@5657.4]
  wire  output_3_25; // @[Switch.scala 41:38:@5658.4]
  wire  _T_15893; // @[Switch.scala 41:52:@5660.4]
  wire  output_3_26; // @[Switch.scala 41:38:@5661.4]
  wire  _T_15896; // @[Switch.scala 41:52:@5663.4]
  wire  output_3_27; // @[Switch.scala 41:38:@5664.4]
  wire  _T_15899; // @[Switch.scala 41:52:@5666.4]
  wire  output_3_28; // @[Switch.scala 41:38:@5667.4]
  wire  _T_15902; // @[Switch.scala 41:52:@5669.4]
  wire  output_3_29; // @[Switch.scala 41:38:@5670.4]
  wire  _T_15905; // @[Switch.scala 41:52:@5672.4]
  wire  output_3_30; // @[Switch.scala 41:38:@5673.4]
  wire  _T_15908; // @[Switch.scala 41:52:@5675.4]
  wire  output_3_31; // @[Switch.scala 41:38:@5676.4]
  wire [7:0] _T_15916; // @[Switch.scala 43:31:@5684.4]
  wire [15:0] _T_15924; // @[Switch.scala 43:31:@5692.4]
  wire [7:0] _T_15931; // @[Switch.scala 43:31:@5699.4]
  wire [31:0] _T_15940; // @[Switch.scala 43:31:@5708.4]
  wire  _T_15944; // @[Switch.scala 41:52:@5711.4]
  wire  output_4_0; // @[Switch.scala 41:38:@5712.4]
  wire  _T_15947; // @[Switch.scala 41:52:@5714.4]
  wire  output_4_1; // @[Switch.scala 41:38:@5715.4]
  wire  _T_15950; // @[Switch.scala 41:52:@5717.4]
  wire  output_4_2; // @[Switch.scala 41:38:@5718.4]
  wire  _T_15953; // @[Switch.scala 41:52:@5720.4]
  wire  output_4_3; // @[Switch.scala 41:38:@5721.4]
  wire  _T_15956; // @[Switch.scala 41:52:@5723.4]
  wire  output_4_4; // @[Switch.scala 41:38:@5724.4]
  wire  _T_15959; // @[Switch.scala 41:52:@5726.4]
  wire  output_4_5; // @[Switch.scala 41:38:@5727.4]
  wire  _T_15962; // @[Switch.scala 41:52:@5729.4]
  wire  output_4_6; // @[Switch.scala 41:38:@5730.4]
  wire  _T_15965; // @[Switch.scala 41:52:@5732.4]
  wire  output_4_7; // @[Switch.scala 41:38:@5733.4]
  wire  _T_15968; // @[Switch.scala 41:52:@5735.4]
  wire  output_4_8; // @[Switch.scala 41:38:@5736.4]
  wire  _T_15971; // @[Switch.scala 41:52:@5738.4]
  wire  output_4_9; // @[Switch.scala 41:38:@5739.4]
  wire  _T_15974; // @[Switch.scala 41:52:@5741.4]
  wire  output_4_10; // @[Switch.scala 41:38:@5742.4]
  wire  _T_15977; // @[Switch.scala 41:52:@5744.4]
  wire  output_4_11; // @[Switch.scala 41:38:@5745.4]
  wire  _T_15980; // @[Switch.scala 41:52:@5747.4]
  wire  output_4_12; // @[Switch.scala 41:38:@5748.4]
  wire  _T_15983; // @[Switch.scala 41:52:@5750.4]
  wire  output_4_13; // @[Switch.scala 41:38:@5751.4]
  wire  _T_15986; // @[Switch.scala 41:52:@5753.4]
  wire  output_4_14; // @[Switch.scala 41:38:@5754.4]
  wire  _T_15989; // @[Switch.scala 41:52:@5756.4]
  wire  output_4_15; // @[Switch.scala 41:38:@5757.4]
  wire  _T_15992; // @[Switch.scala 41:52:@5759.4]
  wire  output_4_16; // @[Switch.scala 41:38:@5760.4]
  wire  _T_15995; // @[Switch.scala 41:52:@5762.4]
  wire  output_4_17; // @[Switch.scala 41:38:@5763.4]
  wire  _T_15998; // @[Switch.scala 41:52:@5765.4]
  wire  output_4_18; // @[Switch.scala 41:38:@5766.4]
  wire  _T_16001; // @[Switch.scala 41:52:@5768.4]
  wire  output_4_19; // @[Switch.scala 41:38:@5769.4]
  wire  _T_16004; // @[Switch.scala 41:52:@5771.4]
  wire  output_4_20; // @[Switch.scala 41:38:@5772.4]
  wire  _T_16007; // @[Switch.scala 41:52:@5774.4]
  wire  output_4_21; // @[Switch.scala 41:38:@5775.4]
  wire  _T_16010; // @[Switch.scala 41:52:@5777.4]
  wire  output_4_22; // @[Switch.scala 41:38:@5778.4]
  wire  _T_16013; // @[Switch.scala 41:52:@5780.4]
  wire  output_4_23; // @[Switch.scala 41:38:@5781.4]
  wire  _T_16016; // @[Switch.scala 41:52:@5783.4]
  wire  output_4_24; // @[Switch.scala 41:38:@5784.4]
  wire  _T_16019; // @[Switch.scala 41:52:@5786.4]
  wire  output_4_25; // @[Switch.scala 41:38:@5787.4]
  wire  _T_16022; // @[Switch.scala 41:52:@5789.4]
  wire  output_4_26; // @[Switch.scala 41:38:@5790.4]
  wire  _T_16025; // @[Switch.scala 41:52:@5792.4]
  wire  output_4_27; // @[Switch.scala 41:38:@5793.4]
  wire  _T_16028; // @[Switch.scala 41:52:@5795.4]
  wire  output_4_28; // @[Switch.scala 41:38:@5796.4]
  wire  _T_16031; // @[Switch.scala 41:52:@5798.4]
  wire  output_4_29; // @[Switch.scala 41:38:@5799.4]
  wire  _T_16034; // @[Switch.scala 41:52:@5801.4]
  wire  output_4_30; // @[Switch.scala 41:38:@5802.4]
  wire  _T_16037; // @[Switch.scala 41:52:@5804.4]
  wire  output_4_31; // @[Switch.scala 41:38:@5805.4]
  wire [7:0] _T_16045; // @[Switch.scala 43:31:@5813.4]
  wire [15:0] _T_16053; // @[Switch.scala 43:31:@5821.4]
  wire [7:0] _T_16060; // @[Switch.scala 43:31:@5828.4]
  wire [31:0] _T_16069; // @[Switch.scala 43:31:@5837.4]
  wire  _T_16073; // @[Switch.scala 41:52:@5840.4]
  wire  output_5_0; // @[Switch.scala 41:38:@5841.4]
  wire  _T_16076; // @[Switch.scala 41:52:@5843.4]
  wire  output_5_1; // @[Switch.scala 41:38:@5844.4]
  wire  _T_16079; // @[Switch.scala 41:52:@5846.4]
  wire  output_5_2; // @[Switch.scala 41:38:@5847.4]
  wire  _T_16082; // @[Switch.scala 41:52:@5849.4]
  wire  output_5_3; // @[Switch.scala 41:38:@5850.4]
  wire  _T_16085; // @[Switch.scala 41:52:@5852.4]
  wire  output_5_4; // @[Switch.scala 41:38:@5853.4]
  wire  _T_16088; // @[Switch.scala 41:52:@5855.4]
  wire  output_5_5; // @[Switch.scala 41:38:@5856.4]
  wire  _T_16091; // @[Switch.scala 41:52:@5858.4]
  wire  output_5_6; // @[Switch.scala 41:38:@5859.4]
  wire  _T_16094; // @[Switch.scala 41:52:@5861.4]
  wire  output_5_7; // @[Switch.scala 41:38:@5862.4]
  wire  _T_16097; // @[Switch.scala 41:52:@5864.4]
  wire  output_5_8; // @[Switch.scala 41:38:@5865.4]
  wire  _T_16100; // @[Switch.scala 41:52:@5867.4]
  wire  output_5_9; // @[Switch.scala 41:38:@5868.4]
  wire  _T_16103; // @[Switch.scala 41:52:@5870.4]
  wire  output_5_10; // @[Switch.scala 41:38:@5871.4]
  wire  _T_16106; // @[Switch.scala 41:52:@5873.4]
  wire  output_5_11; // @[Switch.scala 41:38:@5874.4]
  wire  _T_16109; // @[Switch.scala 41:52:@5876.4]
  wire  output_5_12; // @[Switch.scala 41:38:@5877.4]
  wire  _T_16112; // @[Switch.scala 41:52:@5879.4]
  wire  output_5_13; // @[Switch.scala 41:38:@5880.4]
  wire  _T_16115; // @[Switch.scala 41:52:@5882.4]
  wire  output_5_14; // @[Switch.scala 41:38:@5883.4]
  wire  _T_16118; // @[Switch.scala 41:52:@5885.4]
  wire  output_5_15; // @[Switch.scala 41:38:@5886.4]
  wire  _T_16121; // @[Switch.scala 41:52:@5888.4]
  wire  output_5_16; // @[Switch.scala 41:38:@5889.4]
  wire  _T_16124; // @[Switch.scala 41:52:@5891.4]
  wire  output_5_17; // @[Switch.scala 41:38:@5892.4]
  wire  _T_16127; // @[Switch.scala 41:52:@5894.4]
  wire  output_5_18; // @[Switch.scala 41:38:@5895.4]
  wire  _T_16130; // @[Switch.scala 41:52:@5897.4]
  wire  output_5_19; // @[Switch.scala 41:38:@5898.4]
  wire  _T_16133; // @[Switch.scala 41:52:@5900.4]
  wire  output_5_20; // @[Switch.scala 41:38:@5901.4]
  wire  _T_16136; // @[Switch.scala 41:52:@5903.4]
  wire  output_5_21; // @[Switch.scala 41:38:@5904.4]
  wire  _T_16139; // @[Switch.scala 41:52:@5906.4]
  wire  output_5_22; // @[Switch.scala 41:38:@5907.4]
  wire  _T_16142; // @[Switch.scala 41:52:@5909.4]
  wire  output_5_23; // @[Switch.scala 41:38:@5910.4]
  wire  _T_16145; // @[Switch.scala 41:52:@5912.4]
  wire  output_5_24; // @[Switch.scala 41:38:@5913.4]
  wire  _T_16148; // @[Switch.scala 41:52:@5915.4]
  wire  output_5_25; // @[Switch.scala 41:38:@5916.4]
  wire  _T_16151; // @[Switch.scala 41:52:@5918.4]
  wire  output_5_26; // @[Switch.scala 41:38:@5919.4]
  wire  _T_16154; // @[Switch.scala 41:52:@5921.4]
  wire  output_5_27; // @[Switch.scala 41:38:@5922.4]
  wire  _T_16157; // @[Switch.scala 41:52:@5924.4]
  wire  output_5_28; // @[Switch.scala 41:38:@5925.4]
  wire  _T_16160; // @[Switch.scala 41:52:@5927.4]
  wire  output_5_29; // @[Switch.scala 41:38:@5928.4]
  wire  _T_16163; // @[Switch.scala 41:52:@5930.4]
  wire  output_5_30; // @[Switch.scala 41:38:@5931.4]
  wire  _T_16166; // @[Switch.scala 41:52:@5933.4]
  wire  output_5_31; // @[Switch.scala 41:38:@5934.4]
  wire [7:0] _T_16174; // @[Switch.scala 43:31:@5942.4]
  wire [15:0] _T_16182; // @[Switch.scala 43:31:@5950.4]
  wire [7:0] _T_16189; // @[Switch.scala 43:31:@5957.4]
  wire [31:0] _T_16198; // @[Switch.scala 43:31:@5966.4]
  wire  _T_16202; // @[Switch.scala 41:52:@5969.4]
  wire  output_6_0; // @[Switch.scala 41:38:@5970.4]
  wire  _T_16205; // @[Switch.scala 41:52:@5972.4]
  wire  output_6_1; // @[Switch.scala 41:38:@5973.4]
  wire  _T_16208; // @[Switch.scala 41:52:@5975.4]
  wire  output_6_2; // @[Switch.scala 41:38:@5976.4]
  wire  _T_16211; // @[Switch.scala 41:52:@5978.4]
  wire  output_6_3; // @[Switch.scala 41:38:@5979.4]
  wire  _T_16214; // @[Switch.scala 41:52:@5981.4]
  wire  output_6_4; // @[Switch.scala 41:38:@5982.4]
  wire  _T_16217; // @[Switch.scala 41:52:@5984.4]
  wire  output_6_5; // @[Switch.scala 41:38:@5985.4]
  wire  _T_16220; // @[Switch.scala 41:52:@5987.4]
  wire  output_6_6; // @[Switch.scala 41:38:@5988.4]
  wire  _T_16223; // @[Switch.scala 41:52:@5990.4]
  wire  output_6_7; // @[Switch.scala 41:38:@5991.4]
  wire  _T_16226; // @[Switch.scala 41:52:@5993.4]
  wire  output_6_8; // @[Switch.scala 41:38:@5994.4]
  wire  _T_16229; // @[Switch.scala 41:52:@5996.4]
  wire  output_6_9; // @[Switch.scala 41:38:@5997.4]
  wire  _T_16232; // @[Switch.scala 41:52:@5999.4]
  wire  output_6_10; // @[Switch.scala 41:38:@6000.4]
  wire  _T_16235; // @[Switch.scala 41:52:@6002.4]
  wire  output_6_11; // @[Switch.scala 41:38:@6003.4]
  wire  _T_16238; // @[Switch.scala 41:52:@6005.4]
  wire  output_6_12; // @[Switch.scala 41:38:@6006.4]
  wire  _T_16241; // @[Switch.scala 41:52:@6008.4]
  wire  output_6_13; // @[Switch.scala 41:38:@6009.4]
  wire  _T_16244; // @[Switch.scala 41:52:@6011.4]
  wire  output_6_14; // @[Switch.scala 41:38:@6012.4]
  wire  _T_16247; // @[Switch.scala 41:52:@6014.4]
  wire  output_6_15; // @[Switch.scala 41:38:@6015.4]
  wire  _T_16250; // @[Switch.scala 41:52:@6017.4]
  wire  output_6_16; // @[Switch.scala 41:38:@6018.4]
  wire  _T_16253; // @[Switch.scala 41:52:@6020.4]
  wire  output_6_17; // @[Switch.scala 41:38:@6021.4]
  wire  _T_16256; // @[Switch.scala 41:52:@6023.4]
  wire  output_6_18; // @[Switch.scala 41:38:@6024.4]
  wire  _T_16259; // @[Switch.scala 41:52:@6026.4]
  wire  output_6_19; // @[Switch.scala 41:38:@6027.4]
  wire  _T_16262; // @[Switch.scala 41:52:@6029.4]
  wire  output_6_20; // @[Switch.scala 41:38:@6030.4]
  wire  _T_16265; // @[Switch.scala 41:52:@6032.4]
  wire  output_6_21; // @[Switch.scala 41:38:@6033.4]
  wire  _T_16268; // @[Switch.scala 41:52:@6035.4]
  wire  output_6_22; // @[Switch.scala 41:38:@6036.4]
  wire  _T_16271; // @[Switch.scala 41:52:@6038.4]
  wire  output_6_23; // @[Switch.scala 41:38:@6039.4]
  wire  _T_16274; // @[Switch.scala 41:52:@6041.4]
  wire  output_6_24; // @[Switch.scala 41:38:@6042.4]
  wire  _T_16277; // @[Switch.scala 41:52:@6044.4]
  wire  output_6_25; // @[Switch.scala 41:38:@6045.4]
  wire  _T_16280; // @[Switch.scala 41:52:@6047.4]
  wire  output_6_26; // @[Switch.scala 41:38:@6048.4]
  wire  _T_16283; // @[Switch.scala 41:52:@6050.4]
  wire  output_6_27; // @[Switch.scala 41:38:@6051.4]
  wire  _T_16286; // @[Switch.scala 41:52:@6053.4]
  wire  output_6_28; // @[Switch.scala 41:38:@6054.4]
  wire  _T_16289; // @[Switch.scala 41:52:@6056.4]
  wire  output_6_29; // @[Switch.scala 41:38:@6057.4]
  wire  _T_16292; // @[Switch.scala 41:52:@6059.4]
  wire  output_6_30; // @[Switch.scala 41:38:@6060.4]
  wire  _T_16295; // @[Switch.scala 41:52:@6062.4]
  wire  output_6_31; // @[Switch.scala 41:38:@6063.4]
  wire [7:0] _T_16303; // @[Switch.scala 43:31:@6071.4]
  wire [15:0] _T_16311; // @[Switch.scala 43:31:@6079.4]
  wire [7:0] _T_16318; // @[Switch.scala 43:31:@6086.4]
  wire [31:0] _T_16327; // @[Switch.scala 43:31:@6095.4]
  wire  _T_16331; // @[Switch.scala 41:52:@6098.4]
  wire  output_7_0; // @[Switch.scala 41:38:@6099.4]
  wire  _T_16334; // @[Switch.scala 41:52:@6101.4]
  wire  output_7_1; // @[Switch.scala 41:38:@6102.4]
  wire  _T_16337; // @[Switch.scala 41:52:@6104.4]
  wire  output_7_2; // @[Switch.scala 41:38:@6105.4]
  wire  _T_16340; // @[Switch.scala 41:52:@6107.4]
  wire  output_7_3; // @[Switch.scala 41:38:@6108.4]
  wire  _T_16343; // @[Switch.scala 41:52:@6110.4]
  wire  output_7_4; // @[Switch.scala 41:38:@6111.4]
  wire  _T_16346; // @[Switch.scala 41:52:@6113.4]
  wire  output_7_5; // @[Switch.scala 41:38:@6114.4]
  wire  _T_16349; // @[Switch.scala 41:52:@6116.4]
  wire  output_7_6; // @[Switch.scala 41:38:@6117.4]
  wire  _T_16352; // @[Switch.scala 41:52:@6119.4]
  wire  output_7_7; // @[Switch.scala 41:38:@6120.4]
  wire  _T_16355; // @[Switch.scala 41:52:@6122.4]
  wire  output_7_8; // @[Switch.scala 41:38:@6123.4]
  wire  _T_16358; // @[Switch.scala 41:52:@6125.4]
  wire  output_7_9; // @[Switch.scala 41:38:@6126.4]
  wire  _T_16361; // @[Switch.scala 41:52:@6128.4]
  wire  output_7_10; // @[Switch.scala 41:38:@6129.4]
  wire  _T_16364; // @[Switch.scala 41:52:@6131.4]
  wire  output_7_11; // @[Switch.scala 41:38:@6132.4]
  wire  _T_16367; // @[Switch.scala 41:52:@6134.4]
  wire  output_7_12; // @[Switch.scala 41:38:@6135.4]
  wire  _T_16370; // @[Switch.scala 41:52:@6137.4]
  wire  output_7_13; // @[Switch.scala 41:38:@6138.4]
  wire  _T_16373; // @[Switch.scala 41:52:@6140.4]
  wire  output_7_14; // @[Switch.scala 41:38:@6141.4]
  wire  _T_16376; // @[Switch.scala 41:52:@6143.4]
  wire  output_7_15; // @[Switch.scala 41:38:@6144.4]
  wire  _T_16379; // @[Switch.scala 41:52:@6146.4]
  wire  output_7_16; // @[Switch.scala 41:38:@6147.4]
  wire  _T_16382; // @[Switch.scala 41:52:@6149.4]
  wire  output_7_17; // @[Switch.scala 41:38:@6150.4]
  wire  _T_16385; // @[Switch.scala 41:52:@6152.4]
  wire  output_7_18; // @[Switch.scala 41:38:@6153.4]
  wire  _T_16388; // @[Switch.scala 41:52:@6155.4]
  wire  output_7_19; // @[Switch.scala 41:38:@6156.4]
  wire  _T_16391; // @[Switch.scala 41:52:@6158.4]
  wire  output_7_20; // @[Switch.scala 41:38:@6159.4]
  wire  _T_16394; // @[Switch.scala 41:52:@6161.4]
  wire  output_7_21; // @[Switch.scala 41:38:@6162.4]
  wire  _T_16397; // @[Switch.scala 41:52:@6164.4]
  wire  output_7_22; // @[Switch.scala 41:38:@6165.4]
  wire  _T_16400; // @[Switch.scala 41:52:@6167.4]
  wire  output_7_23; // @[Switch.scala 41:38:@6168.4]
  wire  _T_16403; // @[Switch.scala 41:52:@6170.4]
  wire  output_7_24; // @[Switch.scala 41:38:@6171.4]
  wire  _T_16406; // @[Switch.scala 41:52:@6173.4]
  wire  output_7_25; // @[Switch.scala 41:38:@6174.4]
  wire  _T_16409; // @[Switch.scala 41:52:@6176.4]
  wire  output_7_26; // @[Switch.scala 41:38:@6177.4]
  wire  _T_16412; // @[Switch.scala 41:52:@6179.4]
  wire  output_7_27; // @[Switch.scala 41:38:@6180.4]
  wire  _T_16415; // @[Switch.scala 41:52:@6182.4]
  wire  output_7_28; // @[Switch.scala 41:38:@6183.4]
  wire  _T_16418; // @[Switch.scala 41:52:@6185.4]
  wire  output_7_29; // @[Switch.scala 41:38:@6186.4]
  wire  _T_16421; // @[Switch.scala 41:52:@6188.4]
  wire  output_7_30; // @[Switch.scala 41:38:@6189.4]
  wire  _T_16424; // @[Switch.scala 41:52:@6191.4]
  wire  output_7_31; // @[Switch.scala 41:38:@6192.4]
  wire [7:0] _T_16432; // @[Switch.scala 43:31:@6200.4]
  wire [15:0] _T_16440; // @[Switch.scala 43:31:@6208.4]
  wire [7:0] _T_16447; // @[Switch.scala 43:31:@6215.4]
  wire [31:0] _T_16456; // @[Switch.scala 43:31:@6224.4]
  wire  _T_16460; // @[Switch.scala 41:52:@6227.4]
  wire  output_8_0; // @[Switch.scala 41:38:@6228.4]
  wire  _T_16463; // @[Switch.scala 41:52:@6230.4]
  wire  output_8_1; // @[Switch.scala 41:38:@6231.4]
  wire  _T_16466; // @[Switch.scala 41:52:@6233.4]
  wire  output_8_2; // @[Switch.scala 41:38:@6234.4]
  wire  _T_16469; // @[Switch.scala 41:52:@6236.4]
  wire  output_8_3; // @[Switch.scala 41:38:@6237.4]
  wire  _T_16472; // @[Switch.scala 41:52:@6239.4]
  wire  output_8_4; // @[Switch.scala 41:38:@6240.4]
  wire  _T_16475; // @[Switch.scala 41:52:@6242.4]
  wire  output_8_5; // @[Switch.scala 41:38:@6243.4]
  wire  _T_16478; // @[Switch.scala 41:52:@6245.4]
  wire  output_8_6; // @[Switch.scala 41:38:@6246.4]
  wire  _T_16481; // @[Switch.scala 41:52:@6248.4]
  wire  output_8_7; // @[Switch.scala 41:38:@6249.4]
  wire  _T_16484; // @[Switch.scala 41:52:@6251.4]
  wire  output_8_8; // @[Switch.scala 41:38:@6252.4]
  wire  _T_16487; // @[Switch.scala 41:52:@6254.4]
  wire  output_8_9; // @[Switch.scala 41:38:@6255.4]
  wire  _T_16490; // @[Switch.scala 41:52:@6257.4]
  wire  output_8_10; // @[Switch.scala 41:38:@6258.4]
  wire  _T_16493; // @[Switch.scala 41:52:@6260.4]
  wire  output_8_11; // @[Switch.scala 41:38:@6261.4]
  wire  _T_16496; // @[Switch.scala 41:52:@6263.4]
  wire  output_8_12; // @[Switch.scala 41:38:@6264.4]
  wire  _T_16499; // @[Switch.scala 41:52:@6266.4]
  wire  output_8_13; // @[Switch.scala 41:38:@6267.4]
  wire  _T_16502; // @[Switch.scala 41:52:@6269.4]
  wire  output_8_14; // @[Switch.scala 41:38:@6270.4]
  wire  _T_16505; // @[Switch.scala 41:52:@6272.4]
  wire  output_8_15; // @[Switch.scala 41:38:@6273.4]
  wire  _T_16508; // @[Switch.scala 41:52:@6275.4]
  wire  output_8_16; // @[Switch.scala 41:38:@6276.4]
  wire  _T_16511; // @[Switch.scala 41:52:@6278.4]
  wire  output_8_17; // @[Switch.scala 41:38:@6279.4]
  wire  _T_16514; // @[Switch.scala 41:52:@6281.4]
  wire  output_8_18; // @[Switch.scala 41:38:@6282.4]
  wire  _T_16517; // @[Switch.scala 41:52:@6284.4]
  wire  output_8_19; // @[Switch.scala 41:38:@6285.4]
  wire  _T_16520; // @[Switch.scala 41:52:@6287.4]
  wire  output_8_20; // @[Switch.scala 41:38:@6288.4]
  wire  _T_16523; // @[Switch.scala 41:52:@6290.4]
  wire  output_8_21; // @[Switch.scala 41:38:@6291.4]
  wire  _T_16526; // @[Switch.scala 41:52:@6293.4]
  wire  output_8_22; // @[Switch.scala 41:38:@6294.4]
  wire  _T_16529; // @[Switch.scala 41:52:@6296.4]
  wire  output_8_23; // @[Switch.scala 41:38:@6297.4]
  wire  _T_16532; // @[Switch.scala 41:52:@6299.4]
  wire  output_8_24; // @[Switch.scala 41:38:@6300.4]
  wire  _T_16535; // @[Switch.scala 41:52:@6302.4]
  wire  output_8_25; // @[Switch.scala 41:38:@6303.4]
  wire  _T_16538; // @[Switch.scala 41:52:@6305.4]
  wire  output_8_26; // @[Switch.scala 41:38:@6306.4]
  wire  _T_16541; // @[Switch.scala 41:52:@6308.4]
  wire  output_8_27; // @[Switch.scala 41:38:@6309.4]
  wire  _T_16544; // @[Switch.scala 41:52:@6311.4]
  wire  output_8_28; // @[Switch.scala 41:38:@6312.4]
  wire  _T_16547; // @[Switch.scala 41:52:@6314.4]
  wire  output_8_29; // @[Switch.scala 41:38:@6315.4]
  wire  _T_16550; // @[Switch.scala 41:52:@6317.4]
  wire  output_8_30; // @[Switch.scala 41:38:@6318.4]
  wire  _T_16553; // @[Switch.scala 41:52:@6320.4]
  wire  output_8_31; // @[Switch.scala 41:38:@6321.4]
  wire [7:0] _T_16561; // @[Switch.scala 43:31:@6329.4]
  wire [15:0] _T_16569; // @[Switch.scala 43:31:@6337.4]
  wire [7:0] _T_16576; // @[Switch.scala 43:31:@6344.4]
  wire [31:0] _T_16585; // @[Switch.scala 43:31:@6353.4]
  wire  _T_16589; // @[Switch.scala 41:52:@6356.4]
  wire  output_9_0; // @[Switch.scala 41:38:@6357.4]
  wire  _T_16592; // @[Switch.scala 41:52:@6359.4]
  wire  output_9_1; // @[Switch.scala 41:38:@6360.4]
  wire  _T_16595; // @[Switch.scala 41:52:@6362.4]
  wire  output_9_2; // @[Switch.scala 41:38:@6363.4]
  wire  _T_16598; // @[Switch.scala 41:52:@6365.4]
  wire  output_9_3; // @[Switch.scala 41:38:@6366.4]
  wire  _T_16601; // @[Switch.scala 41:52:@6368.4]
  wire  output_9_4; // @[Switch.scala 41:38:@6369.4]
  wire  _T_16604; // @[Switch.scala 41:52:@6371.4]
  wire  output_9_5; // @[Switch.scala 41:38:@6372.4]
  wire  _T_16607; // @[Switch.scala 41:52:@6374.4]
  wire  output_9_6; // @[Switch.scala 41:38:@6375.4]
  wire  _T_16610; // @[Switch.scala 41:52:@6377.4]
  wire  output_9_7; // @[Switch.scala 41:38:@6378.4]
  wire  _T_16613; // @[Switch.scala 41:52:@6380.4]
  wire  output_9_8; // @[Switch.scala 41:38:@6381.4]
  wire  _T_16616; // @[Switch.scala 41:52:@6383.4]
  wire  output_9_9; // @[Switch.scala 41:38:@6384.4]
  wire  _T_16619; // @[Switch.scala 41:52:@6386.4]
  wire  output_9_10; // @[Switch.scala 41:38:@6387.4]
  wire  _T_16622; // @[Switch.scala 41:52:@6389.4]
  wire  output_9_11; // @[Switch.scala 41:38:@6390.4]
  wire  _T_16625; // @[Switch.scala 41:52:@6392.4]
  wire  output_9_12; // @[Switch.scala 41:38:@6393.4]
  wire  _T_16628; // @[Switch.scala 41:52:@6395.4]
  wire  output_9_13; // @[Switch.scala 41:38:@6396.4]
  wire  _T_16631; // @[Switch.scala 41:52:@6398.4]
  wire  output_9_14; // @[Switch.scala 41:38:@6399.4]
  wire  _T_16634; // @[Switch.scala 41:52:@6401.4]
  wire  output_9_15; // @[Switch.scala 41:38:@6402.4]
  wire  _T_16637; // @[Switch.scala 41:52:@6404.4]
  wire  output_9_16; // @[Switch.scala 41:38:@6405.4]
  wire  _T_16640; // @[Switch.scala 41:52:@6407.4]
  wire  output_9_17; // @[Switch.scala 41:38:@6408.4]
  wire  _T_16643; // @[Switch.scala 41:52:@6410.4]
  wire  output_9_18; // @[Switch.scala 41:38:@6411.4]
  wire  _T_16646; // @[Switch.scala 41:52:@6413.4]
  wire  output_9_19; // @[Switch.scala 41:38:@6414.4]
  wire  _T_16649; // @[Switch.scala 41:52:@6416.4]
  wire  output_9_20; // @[Switch.scala 41:38:@6417.4]
  wire  _T_16652; // @[Switch.scala 41:52:@6419.4]
  wire  output_9_21; // @[Switch.scala 41:38:@6420.4]
  wire  _T_16655; // @[Switch.scala 41:52:@6422.4]
  wire  output_9_22; // @[Switch.scala 41:38:@6423.4]
  wire  _T_16658; // @[Switch.scala 41:52:@6425.4]
  wire  output_9_23; // @[Switch.scala 41:38:@6426.4]
  wire  _T_16661; // @[Switch.scala 41:52:@6428.4]
  wire  output_9_24; // @[Switch.scala 41:38:@6429.4]
  wire  _T_16664; // @[Switch.scala 41:52:@6431.4]
  wire  output_9_25; // @[Switch.scala 41:38:@6432.4]
  wire  _T_16667; // @[Switch.scala 41:52:@6434.4]
  wire  output_9_26; // @[Switch.scala 41:38:@6435.4]
  wire  _T_16670; // @[Switch.scala 41:52:@6437.4]
  wire  output_9_27; // @[Switch.scala 41:38:@6438.4]
  wire  _T_16673; // @[Switch.scala 41:52:@6440.4]
  wire  output_9_28; // @[Switch.scala 41:38:@6441.4]
  wire  _T_16676; // @[Switch.scala 41:52:@6443.4]
  wire  output_9_29; // @[Switch.scala 41:38:@6444.4]
  wire  _T_16679; // @[Switch.scala 41:52:@6446.4]
  wire  output_9_30; // @[Switch.scala 41:38:@6447.4]
  wire  _T_16682; // @[Switch.scala 41:52:@6449.4]
  wire  output_9_31; // @[Switch.scala 41:38:@6450.4]
  wire [7:0] _T_16690; // @[Switch.scala 43:31:@6458.4]
  wire [15:0] _T_16698; // @[Switch.scala 43:31:@6466.4]
  wire [7:0] _T_16705; // @[Switch.scala 43:31:@6473.4]
  wire [31:0] _T_16714; // @[Switch.scala 43:31:@6482.4]
  wire  _T_16718; // @[Switch.scala 41:52:@6485.4]
  wire  output_10_0; // @[Switch.scala 41:38:@6486.4]
  wire  _T_16721; // @[Switch.scala 41:52:@6488.4]
  wire  output_10_1; // @[Switch.scala 41:38:@6489.4]
  wire  _T_16724; // @[Switch.scala 41:52:@6491.4]
  wire  output_10_2; // @[Switch.scala 41:38:@6492.4]
  wire  _T_16727; // @[Switch.scala 41:52:@6494.4]
  wire  output_10_3; // @[Switch.scala 41:38:@6495.4]
  wire  _T_16730; // @[Switch.scala 41:52:@6497.4]
  wire  output_10_4; // @[Switch.scala 41:38:@6498.4]
  wire  _T_16733; // @[Switch.scala 41:52:@6500.4]
  wire  output_10_5; // @[Switch.scala 41:38:@6501.4]
  wire  _T_16736; // @[Switch.scala 41:52:@6503.4]
  wire  output_10_6; // @[Switch.scala 41:38:@6504.4]
  wire  _T_16739; // @[Switch.scala 41:52:@6506.4]
  wire  output_10_7; // @[Switch.scala 41:38:@6507.4]
  wire  _T_16742; // @[Switch.scala 41:52:@6509.4]
  wire  output_10_8; // @[Switch.scala 41:38:@6510.4]
  wire  _T_16745; // @[Switch.scala 41:52:@6512.4]
  wire  output_10_9; // @[Switch.scala 41:38:@6513.4]
  wire  _T_16748; // @[Switch.scala 41:52:@6515.4]
  wire  output_10_10; // @[Switch.scala 41:38:@6516.4]
  wire  _T_16751; // @[Switch.scala 41:52:@6518.4]
  wire  output_10_11; // @[Switch.scala 41:38:@6519.4]
  wire  _T_16754; // @[Switch.scala 41:52:@6521.4]
  wire  output_10_12; // @[Switch.scala 41:38:@6522.4]
  wire  _T_16757; // @[Switch.scala 41:52:@6524.4]
  wire  output_10_13; // @[Switch.scala 41:38:@6525.4]
  wire  _T_16760; // @[Switch.scala 41:52:@6527.4]
  wire  output_10_14; // @[Switch.scala 41:38:@6528.4]
  wire  _T_16763; // @[Switch.scala 41:52:@6530.4]
  wire  output_10_15; // @[Switch.scala 41:38:@6531.4]
  wire  _T_16766; // @[Switch.scala 41:52:@6533.4]
  wire  output_10_16; // @[Switch.scala 41:38:@6534.4]
  wire  _T_16769; // @[Switch.scala 41:52:@6536.4]
  wire  output_10_17; // @[Switch.scala 41:38:@6537.4]
  wire  _T_16772; // @[Switch.scala 41:52:@6539.4]
  wire  output_10_18; // @[Switch.scala 41:38:@6540.4]
  wire  _T_16775; // @[Switch.scala 41:52:@6542.4]
  wire  output_10_19; // @[Switch.scala 41:38:@6543.4]
  wire  _T_16778; // @[Switch.scala 41:52:@6545.4]
  wire  output_10_20; // @[Switch.scala 41:38:@6546.4]
  wire  _T_16781; // @[Switch.scala 41:52:@6548.4]
  wire  output_10_21; // @[Switch.scala 41:38:@6549.4]
  wire  _T_16784; // @[Switch.scala 41:52:@6551.4]
  wire  output_10_22; // @[Switch.scala 41:38:@6552.4]
  wire  _T_16787; // @[Switch.scala 41:52:@6554.4]
  wire  output_10_23; // @[Switch.scala 41:38:@6555.4]
  wire  _T_16790; // @[Switch.scala 41:52:@6557.4]
  wire  output_10_24; // @[Switch.scala 41:38:@6558.4]
  wire  _T_16793; // @[Switch.scala 41:52:@6560.4]
  wire  output_10_25; // @[Switch.scala 41:38:@6561.4]
  wire  _T_16796; // @[Switch.scala 41:52:@6563.4]
  wire  output_10_26; // @[Switch.scala 41:38:@6564.4]
  wire  _T_16799; // @[Switch.scala 41:52:@6566.4]
  wire  output_10_27; // @[Switch.scala 41:38:@6567.4]
  wire  _T_16802; // @[Switch.scala 41:52:@6569.4]
  wire  output_10_28; // @[Switch.scala 41:38:@6570.4]
  wire  _T_16805; // @[Switch.scala 41:52:@6572.4]
  wire  output_10_29; // @[Switch.scala 41:38:@6573.4]
  wire  _T_16808; // @[Switch.scala 41:52:@6575.4]
  wire  output_10_30; // @[Switch.scala 41:38:@6576.4]
  wire  _T_16811; // @[Switch.scala 41:52:@6578.4]
  wire  output_10_31; // @[Switch.scala 41:38:@6579.4]
  wire [7:0] _T_16819; // @[Switch.scala 43:31:@6587.4]
  wire [15:0] _T_16827; // @[Switch.scala 43:31:@6595.4]
  wire [7:0] _T_16834; // @[Switch.scala 43:31:@6602.4]
  wire [31:0] _T_16843; // @[Switch.scala 43:31:@6611.4]
  wire  _T_16847; // @[Switch.scala 41:52:@6614.4]
  wire  output_11_0; // @[Switch.scala 41:38:@6615.4]
  wire  _T_16850; // @[Switch.scala 41:52:@6617.4]
  wire  output_11_1; // @[Switch.scala 41:38:@6618.4]
  wire  _T_16853; // @[Switch.scala 41:52:@6620.4]
  wire  output_11_2; // @[Switch.scala 41:38:@6621.4]
  wire  _T_16856; // @[Switch.scala 41:52:@6623.4]
  wire  output_11_3; // @[Switch.scala 41:38:@6624.4]
  wire  _T_16859; // @[Switch.scala 41:52:@6626.4]
  wire  output_11_4; // @[Switch.scala 41:38:@6627.4]
  wire  _T_16862; // @[Switch.scala 41:52:@6629.4]
  wire  output_11_5; // @[Switch.scala 41:38:@6630.4]
  wire  _T_16865; // @[Switch.scala 41:52:@6632.4]
  wire  output_11_6; // @[Switch.scala 41:38:@6633.4]
  wire  _T_16868; // @[Switch.scala 41:52:@6635.4]
  wire  output_11_7; // @[Switch.scala 41:38:@6636.4]
  wire  _T_16871; // @[Switch.scala 41:52:@6638.4]
  wire  output_11_8; // @[Switch.scala 41:38:@6639.4]
  wire  _T_16874; // @[Switch.scala 41:52:@6641.4]
  wire  output_11_9; // @[Switch.scala 41:38:@6642.4]
  wire  _T_16877; // @[Switch.scala 41:52:@6644.4]
  wire  output_11_10; // @[Switch.scala 41:38:@6645.4]
  wire  _T_16880; // @[Switch.scala 41:52:@6647.4]
  wire  output_11_11; // @[Switch.scala 41:38:@6648.4]
  wire  _T_16883; // @[Switch.scala 41:52:@6650.4]
  wire  output_11_12; // @[Switch.scala 41:38:@6651.4]
  wire  _T_16886; // @[Switch.scala 41:52:@6653.4]
  wire  output_11_13; // @[Switch.scala 41:38:@6654.4]
  wire  _T_16889; // @[Switch.scala 41:52:@6656.4]
  wire  output_11_14; // @[Switch.scala 41:38:@6657.4]
  wire  _T_16892; // @[Switch.scala 41:52:@6659.4]
  wire  output_11_15; // @[Switch.scala 41:38:@6660.4]
  wire  _T_16895; // @[Switch.scala 41:52:@6662.4]
  wire  output_11_16; // @[Switch.scala 41:38:@6663.4]
  wire  _T_16898; // @[Switch.scala 41:52:@6665.4]
  wire  output_11_17; // @[Switch.scala 41:38:@6666.4]
  wire  _T_16901; // @[Switch.scala 41:52:@6668.4]
  wire  output_11_18; // @[Switch.scala 41:38:@6669.4]
  wire  _T_16904; // @[Switch.scala 41:52:@6671.4]
  wire  output_11_19; // @[Switch.scala 41:38:@6672.4]
  wire  _T_16907; // @[Switch.scala 41:52:@6674.4]
  wire  output_11_20; // @[Switch.scala 41:38:@6675.4]
  wire  _T_16910; // @[Switch.scala 41:52:@6677.4]
  wire  output_11_21; // @[Switch.scala 41:38:@6678.4]
  wire  _T_16913; // @[Switch.scala 41:52:@6680.4]
  wire  output_11_22; // @[Switch.scala 41:38:@6681.4]
  wire  _T_16916; // @[Switch.scala 41:52:@6683.4]
  wire  output_11_23; // @[Switch.scala 41:38:@6684.4]
  wire  _T_16919; // @[Switch.scala 41:52:@6686.4]
  wire  output_11_24; // @[Switch.scala 41:38:@6687.4]
  wire  _T_16922; // @[Switch.scala 41:52:@6689.4]
  wire  output_11_25; // @[Switch.scala 41:38:@6690.4]
  wire  _T_16925; // @[Switch.scala 41:52:@6692.4]
  wire  output_11_26; // @[Switch.scala 41:38:@6693.4]
  wire  _T_16928; // @[Switch.scala 41:52:@6695.4]
  wire  output_11_27; // @[Switch.scala 41:38:@6696.4]
  wire  _T_16931; // @[Switch.scala 41:52:@6698.4]
  wire  output_11_28; // @[Switch.scala 41:38:@6699.4]
  wire  _T_16934; // @[Switch.scala 41:52:@6701.4]
  wire  output_11_29; // @[Switch.scala 41:38:@6702.4]
  wire  _T_16937; // @[Switch.scala 41:52:@6704.4]
  wire  output_11_30; // @[Switch.scala 41:38:@6705.4]
  wire  _T_16940; // @[Switch.scala 41:52:@6707.4]
  wire  output_11_31; // @[Switch.scala 41:38:@6708.4]
  wire [7:0] _T_16948; // @[Switch.scala 43:31:@6716.4]
  wire [15:0] _T_16956; // @[Switch.scala 43:31:@6724.4]
  wire [7:0] _T_16963; // @[Switch.scala 43:31:@6731.4]
  wire [31:0] _T_16972; // @[Switch.scala 43:31:@6740.4]
  wire  _T_16976; // @[Switch.scala 41:52:@6743.4]
  wire  output_12_0; // @[Switch.scala 41:38:@6744.4]
  wire  _T_16979; // @[Switch.scala 41:52:@6746.4]
  wire  output_12_1; // @[Switch.scala 41:38:@6747.4]
  wire  _T_16982; // @[Switch.scala 41:52:@6749.4]
  wire  output_12_2; // @[Switch.scala 41:38:@6750.4]
  wire  _T_16985; // @[Switch.scala 41:52:@6752.4]
  wire  output_12_3; // @[Switch.scala 41:38:@6753.4]
  wire  _T_16988; // @[Switch.scala 41:52:@6755.4]
  wire  output_12_4; // @[Switch.scala 41:38:@6756.4]
  wire  _T_16991; // @[Switch.scala 41:52:@6758.4]
  wire  output_12_5; // @[Switch.scala 41:38:@6759.4]
  wire  _T_16994; // @[Switch.scala 41:52:@6761.4]
  wire  output_12_6; // @[Switch.scala 41:38:@6762.4]
  wire  _T_16997; // @[Switch.scala 41:52:@6764.4]
  wire  output_12_7; // @[Switch.scala 41:38:@6765.4]
  wire  _T_17000; // @[Switch.scala 41:52:@6767.4]
  wire  output_12_8; // @[Switch.scala 41:38:@6768.4]
  wire  _T_17003; // @[Switch.scala 41:52:@6770.4]
  wire  output_12_9; // @[Switch.scala 41:38:@6771.4]
  wire  _T_17006; // @[Switch.scala 41:52:@6773.4]
  wire  output_12_10; // @[Switch.scala 41:38:@6774.4]
  wire  _T_17009; // @[Switch.scala 41:52:@6776.4]
  wire  output_12_11; // @[Switch.scala 41:38:@6777.4]
  wire  _T_17012; // @[Switch.scala 41:52:@6779.4]
  wire  output_12_12; // @[Switch.scala 41:38:@6780.4]
  wire  _T_17015; // @[Switch.scala 41:52:@6782.4]
  wire  output_12_13; // @[Switch.scala 41:38:@6783.4]
  wire  _T_17018; // @[Switch.scala 41:52:@6785.4]
  wire  output_12_14; // @[Switch.scala 41:38:@6786.4]
  wire  _T_17021; // @[Switch.scala 41:52:@6788.4]
  wire  output_12_15; // @[Switch.scala 41:38:@6789.4]
  wire  _T_17024; // @[Switch.scala 41:52:@6791.4]
  wire  output_12_16; // @[Switch.scala 41:38:@6792.4]
  wire  _T_17027; // @[Switch.scala 41:52:@6794.4]
  wire  output_12_17; // @[Switch.scala 41:38:@6795.4]
  wire  _T_17030; // @[Switch.scala 41:52:@6797.4]
  wire  output_12_18; // @[Switch.scala 41:38:@6798.4]
  wire  _T_17033; // @[Switch.scala 41:52:@6800.4]
  wire  output_12_19; // @[Switch.scala 41:38:@6801.4]
  wire  _T_17036; // @[Switch.scala 41:52:@6803.4]
  wire  output_12_20; // @[Switch.scala 41:38:@6804.4]
  wire  _T_17039; // @[Switch.scala 41:52:@6806.4]
  wire  output_12_21; // @[Switch.scala 41:38:@6807.4]
  wire  _T_17042; // @[Switch.scala 41:52:@6809.4]
  wire  output_12_22; // @[Switch.scala 41:38:@6810.4]
  wire  _T_17045; // @[Switch.scala 41:52:@6812.4]
  wire  output_12_23; // @[Switch.scala 41:38:@6813.4]
  wire  _T_17048; // @[Switch.scala 41:52:@6815.4]
  wire  output_12_24; // @[Switch.scala 41:38:@6816.4]
  wire  _T_17051; // @[Switch.scala 41:52:@6818.4]
  wire  output_12_25; // @[Switch.scala 41:38:@6819.4]
  wire  _T_17054; // @[Switch.scala 41:52:@6821.4]
  wire  output_12_26; // @[Switch.scala 41:38:@6822.4]
  wire  _T_17057; // @[Switch.scala 41:52:@6824.4]
  wire  output_12_27; // @[Switch.scala 41:38:@6825.4]
  wire  _T_17060; // @[Switch.scala 41:52:@6827.4]
  wire  output_12_28; // @[Switch.scala 41:38:@6828.4]
  wire  _T_17063; // @[Switch.scala 41:52:@6830.4]
  wire  output_12_29; // @[Switch.scala 41:38:@6831.4]
  wire  _T_17066; // @[Switch.scala 41:52:@6833.4]
  wire  output_12_30; // @[Switch.scala 41:38:@6834.4]
  wire  _T_17069; // @[Switch.scala 41:52:@6836.4]
  wire  output_12_31; // @[Switch.scala 41:38:@6837.4]
  wire [7:0] _T_17077; // @[Switch.scala 43:31:@6845.4]
  wire [15:0] _T_17085; // @[Switch.scala 43:31:@6853.4]
  wire [7:0] _T_17092; // @[Switch.scala 43:31:@6860.4]
  wire [31:0] _T_17101; // @[Switch.scala 43:31:@6869.4]
  wire  _T_17105; // @[Switch.scala 41:52:@6872.4]
  wire  output_13_0; // @[Switch.scala 41:38:@6873.4]
  wire  _T_17108; // @[Switch.scala 41:52:@6875.4]
  wire  output_13_1; // @[Switch.scala 41:38:@6876.4]
  wire  _T_17111; // @[Switch.scala 41:52:@6878.4]
  wire  output_13_2; // @[Switch.scala 41:38:@6879.4]
  wire  _T_17114; // @[Switch.scala 41:52:@6881.4]
  wire  output_13_3; // @[Switch.scala 41:38:@6882.4]
  wire  _T_17117; // @[Switch.scala 41:52:@6884.4]
  wire  output_13_4; // @[Switch.scala 41:38:@6885.4]
  wire  _T_17120; // @[Switch.scala 41:52:@6887.4]
  wire  output_13_5; // @[Switch.scala 41:38:@6888.4]
  wire  _T_17123; // @[Switch.scala 41:52:@6890.4]
  wire  output_13_6; // @[Switch.scala 41:38:@6891.4]
  wire  _T_17126; // @[Switch.scala 41:52:@6893.4]
  wire  output_13_7; // @[Switch.scala 41:38:@6894.4]
  wire  _T_17129; // @[Switch.scala 41:52:@6896.4]
  wire  output_13_8; // @[Switch.scala 41:38:@6897.4]
  wire  _T_17132; // @[Switch.scala 41:52:@6899.4]
  wire  output_13_9; // @[Switch.scala 41:38:@6900.4]
  wire  _T_17135; // @[Switch.scala 41:52:@6902.4]
  wire  output_13_10; // @[Switch.scala 41:38:@6903.4]
  wire  _T_17138; // @[Switch.scala 41:52:@6905.4]
  wire  output_13_11; // @[Switch.scala 41:38:@6906.4]
  wire  _T_17141; // @[Switch.scala 41:52:@6908.4]
  wire  output_13_12; // @[Switch.scala 41:38:@6909.4]
  wire  _T_17144; // @[Switch.scala 41:52:@6911.4]
  wire  output_13_13; // @[Switch.scala 41:38:@6912.4]
  wire  _T_17147; // @[Switch.scala 41:52:@6914.4]
  wire  output_13_14; // @[Switch.scala 41:38:@6915.4]
  wire  _T_17150; // @[Switch.scala 41:52:@6917.4]
  wire  output_13_15; // @[Switch.scala 41:38:@6918.4]
  wire  _T_17153; // @[Switch.scala 41:52:@6920.4]
  wire  output_13_16; // @[Switch.scala 41:38:@6921.4]
  wire  _T_17156; // @[Switch.scala 41:52:@6923.4]
  wire  output_13_17; // @[Switch.scala 41:38:@6924.4]
  wire  _T_17159; // @[Switch.scala 41:52:@6926.4]
  wire  output_13_18; // @[Switch.scala 41:38:@6927.4]
  wire  _T_17162; // @[Switch.scala 41:52:@6929.4]
  wire  output_13_19; // @[Switch.scala 41:38:@6930.4]
  wire  _T_17165; // @[Switch.scala 41:52:@6932.4]
  wire  output_13_20; // @[Switch.scala 41:38:@6933.4]
  wire  _T_17168; // @[Switch.scala 41:52:@6935.4]
  wire  output_13_21; // @[Switch.scala 41:38:@6936.4]
  wire  _T_17171; // @[Switch.scala 41:52:@6938.4]
  wire  output_13_22; // @[Switch.scala 41:38:@6939.4]
  wire  _T_17174; // @[Switch.scala 41:52:@6941.4]
  wire  output_13_23; // @[Switch.scala 41:38:@6942.4]
  wire  _T_17177; // @[Switch.scala 41:52:@6944.4]
  wire  output_13_24; // @[Switch.scala 41:38:@6945.4]
  wire  _T_17180; // @[Switch.scala 41:52:@6947.4]
  wire  output_13_25; // @[Switch.scala 41:38:@6948.4]
  wire  _T_17183; // @[Switch.scala 41:52:@6950.4]
  wire  output_13_26; // @[Switch.scala 41:38:@6951.4]
  wire  _T_17186; // @[Switch.scala 41:52:@6953.4]
  wire  output_13_27; // @[Switch.scala 41:38:@6954.4]
  wire  _T_17189; // @[Switch.scala 41:52:@6956.4]
  wire  output_13_28; // @[Switch.scala 41:38:@6957.4]
  wire  _T_17192; // @[Switch.scala 41:52:@6959.4]
  wire  output_13_29; // @[Switch.scala 41:38:@6960.4]
  wire  _T_17195; // @[Switch.scala 41:52:@6962.4]
  wire  output_13_30; // @[Switch.scala 41:38:@6963.4]
  wire  _T_17198; // @[Switch.scala 41:52:@6965.4]
  wire  output_13_31; // @[Switch.scala 41:38:@6966.4]
  wire [7:0] _T_17206; // @[Switch.scala 43:31:@6974.4]
  wire [15:0] _T_17214; // @[Switch.scala 43:31:@6982.4]
  wire [7:0] _T_17221; // @[Switch.scala 43:31:@6989.4]
  wire [31:0] _T_17230; // @[Switch.scala 43:31:@6998.4]
  wire  _T_17234; // @[Switch.scala 41:52:@7001.4]
  wire  output_14_0; // @[Switch.scala 41:38:@7002.4]
  wire  _T_17237; // @[Switch.scala 41:52:@7004.4]
  wire  output_14_1; // @[Switch.scala 41:38:@7005.4]
  wire  _T_17240; // @[Switch.scala 41:52:@7007.4]
  wire  output_14_2; // @[Switch.scala 41:38:@7008.4]
  wire  _T_17243; // @[Switch.scala 41:52:@7010.4]
  wire  output_14_3; // @[Switch.scala 41:38:@7011.4]
  wire  _T_17246; // @[Switch.scala 41:52:@7013.4]
  wire  output_14_4; // @[Switch.scala 41:38:@7014.4]
  wire  _T_17249; // @[Switch.scala 41:52:@7016.4]
  wire  output_14_5; // @[Switch.scala 41:38:@7017.4]
  wire  _T_17252; // @[Switch.scala 41:52:@7019.4]
  wire  output_14_6; // @[Switch.scala 41:38:@7020.4]
  wire  _T_17255; // @[Switch.scala 41:52:@7022.4]
  wire  output_14_7; // @[Switch.scala 41:38:@7023.4]
  wire  _T_17258; // @[Switch.scala 41:52:@7025.4]
  wire  output_14_8; // @[Switch.scala 41:38:@7026.4]
  wire  _T_17261; // @[Switch.scala 41:52:@7028.4]
  wire  output_14_9; // @[Switch.scala 41:38:@7029.4]
  wire  _T_17264; // @[Switch.scala 41:52:@7031.4]
  wire  output_14_10; // @[Switch.scala 41:38:@7032.4]
  wire  _T_17267; // @[Switch.scala 41:52:@7034.4]
  wire  output_14_11; // @[Switch.scala 41:38:@7035.4]
  wire  _T_17270; // @[Switch.scala 41:52:@7037.4]
  wire  output_14_12; // @[Switch.scala 41:38:@7038.4]
  wire  _T_17273; // @[Switch.scala 41:52:@7040.4]
  wire  output_14_13; // @[Switch.scala 41:38:@7041.4]
  wire  _T_17276; // @[Switch.scala 41:52:@7043.4]
  wire  output_14_14; // @[Switch.scala 41:38:@7044.4]
  wire  _T_17279; // @[Switch.scala 41:52:@7046.4]
  wire  output_14_15; // @[Switch.scala 41:38:@7047.4]
  wire  _T_17282; // @[Switch.scala 41:52:@7049.4]
  wire  output_14_16; // @[Switch.scala 41:38:@7050.4]
  wire  _T_17285; // @[Switch.scala 41:52:@7052.4]
  wire  output_14_17; // @[Switch.scala 41:38:@7053.4]
  wire  _T_17288; // @[Switch.scala 41:52:@7055.4]
  wire  output_14_18; // @[Switch.scala 41:38:@7056.4]
  wire  _T_17291; // @[Switch.scala 41:52:@7058.4]
  wire  output_14_19; // @[Switch.scala 41:38:@7059.4]
  wire  _T_17294; // @[Switch.scala 41:52:@7061.4]
  wire  output_14_20; // @[Switch.scala 41:38:@7062.4]
  wire  _T_17297; // @[Switch.scala 41:52:@7064.4]
  wire  output_14_21; // @[Switch.scala 41:38:@7065.4]
  wire  _T_17300; // @[Switch.scala 41:52:@7067.4]
  wire  output_14_22; // @[Switch.scala 41:38:@7068.4]
  wire  _T_17303; // @[Switch.scala 41:52:@7070.4]
  wire  output_14_23; // @[Switch.scala 41:38:@7071.4]
  wire  _T_17306; // @[Switch.scala 41:52:@7073.4]
  wire  output_14_24; // @[Switch.scala 41:38:@7074.4]
  wire  _T_17309; // @[Switch.scala 41:52:@7076.4]
  wire  output_14_25; // @[Switch.scala 41:38:@7077.4]
  wire  _T_17312; // @[Switch.scala 41:52:@7079.4]
  wire  output_14_26; // @[Switch.scala 41:38:@7080.4]
  wire  _T_17315; // @[Switch.scala 41:52:@7082.4]
  wire  output_14_27; // @[Switch.scala 41:38:@7083.4]
  wire  _T_17318; // @[Switch.scala 41:52:@7085.4]
  wire  output_14_28; // @[Switch.scala 41:38:@7086.4]
  wire  _T_17321; // @[Switch.scala 41:52:@7088.4]
  wire  output_14_29; // @[Switch.scala 41:38:@7089.4]
  wire  _T_17324; // @[Switch.scala 41:52:@7091.4]
  wire  output_14_30; // @[Switch.scala 41:38:@7092.4]
  wire  _T_17327; // @[Switch.scala 41:52:@7094.4]
  wire  output_14_31; // @[Switch.scala 41:38:@7095.4]
  wire [7:0] _T_17335; // @[Switch.scala 43:31:@7103.4]
  wire [15:0] _T_17343; // @[Switch.scala 43:31:@7111.4]
  wire [7:0] _T_17350; // @[Switch.scala 43:31:@7118.4]
  wire [31:0] _T_17359; // @[Switch.scala 43:31:@7127.4]
  wire  _T_17363; // @[Switch.scala 41:52:@7130.4]
  wire  output_15_0; // @[Switch.scala 41:38:@7131.4]
  wire  _T_17366; // @[Switch.scala 41:52:@7133.4]
  wire  output_15_1; // @[Switch.scala 41:38:@7134.4]
  wire  _T_17369; // @[Switch.scala 41:52:@7136.4]
  wire  output_15_2; // @[Switch.scala 41:38:@7137.4]
  wire  _T_17372; // @[Switch.scala 41:52:@7139.4]
  wire  output_15_3; // @[Switch.scala 41:38:@7140.4]
  wire  _T_17375; // @[Switch.scala 41:52:@7142.4]
  wire  output_15_4; // @[Switch.scala 41:38:@7143.4]
  wire  _T_17378; // @[Switch.scala 41:52:@7145.4]
  wire  output_15_5; // @[Switch.scala 41:38:@7146.4]
  wire  _T_17381; // @[Switch.scala 41:52:@7148.4]
  wire  output_15_6; // @[Switch.scala 41:38:@7149.4]
  wire  _T_17384; // @[Switch.scala 41:52:@7151.4]
  wire  output_15_7; // @[Switch.scala 41:38:@7152.4]
  wire  _T_17387; // @[Switch.scala 41:52:@7154.4]
  wire  output_15_8; // @[Switch.scala 41:38:@7155.4]
  wire  _T_17390; // @[Switch.scala 41:52:@7157.4]
  wire  output_15_9; // @[Switch.scala 41:38:@7158.4]
  wire  _T_17393; // @[Switch.scala 41:52:@7160.4]
  wire  output_15_10; // @[Switch.scala 41:38:@7161.4]
  wire  _T_17396; // @[Switch.scala 41:52:@7163.4]
  wire  output_15_11; // @[Switch.scala 41:38:@7164.4]
  wire  _T_17399; // @[Switch.scala 41:52:@7166.4]
  wire  output_15_12; // @[Switch.scala 41:38:@7167.4]
  wire  _T_17402; // @[Switch.scala 41:52:@7169.4]
  wire  output_15_13; // @[Switch.scala 41:38:@7170.4]
  wire  _T_17405; // @[Switch.scala 41:52:@7172.4]
  wire  output_15_14; // @[Switch.scala 41:38:@7173.4]
  wire  _T_17408; // @[Switch.scala 41:52:@7175.4]
  wire  output_15_15; // @[Switch.scala 41:38:@7176.4]
  wire  _T_17411; // @[Switch.scala 41:52:@7178.4]
  wire  output_15_16; // @[Switch.scala 41:38:@7179.4]
  wire  _T_17414; // @[Switch.scala 41:52:@7181.4]
  wire  output_15_17; // @[Switch.scala 41:38:@7182.4]
  wire  _T_17417; // @[Switch.scala 41:52:@7184.4]
  wire  output_15_18; // @[Switch.scala 41:38:@7185.4]
  wire  _T_17420; // @[Switch.scala 41:52:@7187.4]
  wire  output_15_19; // @[Switch.scala 41:38:@7188.4]
  wire  _T_17423; // @[Switch.scala 41:52:@7190.4]
  wire  output_15_20; // @[Switch.scala 41:38:@7191.4]
  wire  _T_17426; // @[Switch.scala 41:52:@7193.4]
  wire  output_15_21; // @[Switch.scala 41:38:@7194.4]
  wire  _T_17429; // @[Switch.scala 41:52:@7196.4]
  wire  output_15_22; // @[Switch.scala 41:38:@7197.4]
  wire  _T_17432; // @[Switch.scala 41:52:@7199.4]
  wire  output_15_23; // @[Switch.scala 41:38:@7200.4]
  wire  _T_17435; // @[Switch.scala 41:52:@7202.4]
  wire  output_15_24; // @[Switch.scala 41:38:@7203.4]
  wire  _T_17438; // @[Switch.scala 41:52:@7205.4]
  wire  output_15_25; // @[Switch.scala 41:38:@7206.4]
  wire  _T_17441; // @[Switch.scala 41:52:@7208.4]
  wire  output_15_26; // @[Switch.scala 41:38:@7209.4]
  wire  _T_17444; // @[Switch.scala 41:52:@7211.4]
  wire  output_15_27; // @[Switch.scala 41:38:@7212.4]
  wire  _T_17447; // @[Switch.scala 41:52:@7214.4]
  wire  output_15_28; // @[Switch.scala 41:38:@7215.4]
  wire  _T_17450; // @[Switch.scala 41:52:@7217.4]
  wire  output_15_29; // @[Switch.scala 41:38:@7218.4]
  wire  _T_17453; // @[Switch.scala 41:52:@7220.4]
  wire  output_15_30; // @[Switch.scala 41:38:@7221.4]
  wire  _T_17456; // @[Switch.scala 41:52:@7223.4]
  wire  output_15_31; // @[Switch.scala 41:38:@7224.4]
  wire [7:0] _T_17464; // @[Switch.scala 43:31:@7232.4]
  wire [15:0] _T_17472; // @[Switch.scala 43:31:@7240.4]
  wire [7:0] _T_17479; // @[Switch.scala 43:31:@7247.4]
  wire [31:0] _T_17488; // @[Switch.scala 43:31:@7256.4]
  wire  _T_17492; // @[Switch.scala 41:52:@7259.4]
  wire  output_16_0; // @[Switch.scala 41:38:@7260.4]
  wire  _T_17495; // @[Switch.scala 41:52:@7262.4]
  wire  output_16_1; // @[Switch.scala 41:38:@7263.4]
  wire  _T_17498; // @[Switch.scala 41:52:@7265.4]
  wire  output_16_2; // @[Switch.scala 41:38:@7266.4]
  wire  _T_17501; // @[Switch.scala 41:52:@7268.4]
  wire  output_16_3; // @[Switch.scala 41:38:@7269.4]
  wire  _T_17504; // @[Switch.scala 41:52:@7271.4]
  wire  output_16_4; // @[Switch.scala 41:38:@7272.4]
  wire  _T_17507; // @[Switch.scala 41:52:@7274.4]
  wire  output_16_5; // @[Switch.scala 41:38:@7275.4]
  wire  _T_17510; // @[Switch.scala 41:52:@7277.4]
  wire  output_16_6; // @[Switch.scala 41:38:@7278.4]
  wire  _T_17513; // @[Switch.scala 41:52:@7280.4]
  wire  output_16_7; // @[Switch.scala 41:38:@7281.4]
  wire  _T_17516; // @[Switch.scala 41:52:@7283.4]
  wire  output_16_8; // @[Switch.scala 41:38:@7284.4]
  wire  _T_17519; // @[Switch.scala 41:52:@7286.4]
  wire  output_16_9; // @[Switch.scala 41:38:@7287.4]
  wire  _T_17522; // @[Switch.scala 41:52:@7289.4]
  wire  output_16_10; // @[Switch.scala 41:38:@7290.4]
  wire  _T_17525; // @[Switch.scala 41:52:@7292.4]
  wire  output_16_11; // @[Switch.scala 41:38:@7293.4]
  wire  _T_17528; // @[Switch.scala 41:52:@7295.4]
  wire  output_16_12; // @[Switch.scala 41:38:@7296.4]
  wire  _T_17531; // @[Switch.scala 41:52:@7298.4]
  wire  output_16_13; // @[Switch.scala 41:38:@7299.4]
  wire  _T_17534; // @[Switch.scala 41:52:@7301.4]
  wire  output_16_14; // @[Switch.scala 41:38:@7302.4]
  wire  _T_17537; // @[Switch.scala 41:52:@7304.4]
  wire  output_16_15; // @[Switch.scala 41:38:@7305.4]
  wire  _T_17540; // @[Switch.scala 41:52:@7307.4]
  wire  output_16_16; // @[Switch.scala 41:38:@7308.4]
  wire  _T_17543; // @[Switch.scala 41:52:@7310.4]
  wire  output_16_17; // @[Switch.scala 41:38:@7311.4]
  wire  _T_17546; // @[Switch.scala 41:52:@7313.4]
  wire  output_16_18; // @[Switch.scala 41:38:@7314.4]
  wire  _T_17549; // @[Switch.scala 41:52:@7316.4]
  wire  output_16_19; // @[Switch.scala 41:38:@7317.4]
  wire  _T_17552; // @[Switch.scala 41:52:@7319.4]
  wire  output_16_20; // @[Switch.scala 41:38:@7320.4]
  wire  _T_17555; // @[Switch.scala 41:52:@7322.4]
  wire  output_16_21; // @[Switch.scala 41:38:@7323.4]
  wire  _T_17558; // @[Switch.scala 41:52:@7325.4]
  wire  output_16_22; // @[Switch.scala 41:38:@7326.4]
  wire  _T_17561; // @[Switch.scala 41:52:@7328.4]
  wire  output_16_23; // @[Switch.scala 41:38:@7329.4]
  wire  _T_17564; // @[Switch.scala 41:52:@7331.4]
  wire  output_16_24; // @[Switch.scala 41:38:@7332.4]
  wire  _T_17567; // @[Switch.scala 41:52:@7334.4]
  wire  output_16_25; // @[Switch.scala 41:38:@7335.4]
  wire  _T_17570; // @[Switch.scala 41:52:@7337.4]
  wire  output_16_26; // @[Switch.scala 41:38:@7338.4]
  wire  _T_17573; // @[Switch.scala 41:52:@7340.4]
  wire  output_16_27; // @[Switch.scala 41:38:@7341.4]
  wire  _T_17576; // @[Switch.scala 41:52:@7343.4]
  wire  output_16_28; // @[Switch.scala 41:38:@7344.4]
  wire  _T_17579; // @[Switch.scala 41:52:@7346.4]
  wire  output_16_29; // @[Switch.scala 41:38:@7347.4]
  wire  _T_17582; // @[Switch.scala 41:52:@7349.4]
  wire  output_16_30; // @[Switch.scala 41:38:@7350.4]
  wire  _T_17585; // @[Switch.scala 41:52:@7352.4]
  wire  output_16_31; // @[Switch.scala 41:38:@7353.4]
  wire [7:0] _T_17593; // @[Switch.scala 43:31:@7361.4]
  wire [15:0] _T_17601; // @[Switch.scala 43:31:@7369.4]
  wire [7:0] _T_17608; // @[Switch.scala 43:31:@7376.4]
  wire [31:0] _T_17617; // @[Switch.scala 43:31:@7385.4]
  wire  _T_17621; // @[Switch.scala 41:52:@7388.4]
  wire  output_17_0; // @[Switch.scala 41:38:@7389.4]
  wire  _T_17624; // @[Switch.scala 41:52:@7391.4]
  wire  output_17_1; // @[Switch.scala 41:38:@7392.4]
  wire  _T_17627; // @[Switch.scala 41:52:@7394.4]
  wire  output_17_2; // @[Switch.scala 41:38:@7395.4]
  wire  _T_17630; // @[Switch.scala 41:52:@7397.4]
  wire  output_17_3; // @[Switch.scala 41:38:@7398.4]
  wire  _T_17633; // @[Switch.scala 41:52:@7400.4]
  wire  output_17_4; // @[Switch.scala 41:38:@7401.4]
  wire  _T_17636; // @[Switch.scala 41:52:@7403.4]
  wire  output_17_5; // @[Switch.scala 41:38:@7404.4]
  wire  _T_17639; // @[Switch.scala 41:52:@7406.4]
  wire  output_17_6; // @[Switch.scala 41:38:@7407.4]
  wire  _T_17642; // @[Switch.scala 41:52:@7409.4]
  wire  output_17_7; // @[Switch.scala 41:38:@7410.4]
  wire  _T_17645; // @[Switch.scala 41:52:@7412.4]
  wire  output_17_8; // @[Switch.scala 41:38:@7413.4]
  wire  _T_17648; // @[Switch.scala 41:52:@7415.4]
  wire  output_17_9; // @[Switch.scala 41:38:@7416.4]
  wire  _T_17651; // @[Switch.scala 41:52:@7418.4]
  wire  output_17_10; // @[Switch.scala 41:38:@7419.4]
  wire  _T_17654; // @[Switch.scala 41:52:@7421.4]
  wire  output_17_11; // @[Switch.scala 41:38:@7422.4]
  wire  _T_17657; // @[Switch.scala 41:52:@7424.4]
  wire  output_17_12; // @[Switch.scala 41:38:@7425.4]
  wire  _T_17660; // @[Switch.scala 41:52:@7427.4]
  wire  output_17_13; // @[Switch.scala 41:38:@7428.4]
  wire  _T_17663; // @[Switch.scala 41:52:@7430.4]
  wire  output_17_14; // @[Switch.scala 41:38:@7431.4]
  wire  _T_17666; // @[Switch.scala 41:52:@7433.4]
  wire  output_17_15; // @[Switch.scala 41:38:@7434.4]
  wire  _T_17669; // @[Switch.scala 41:52:@7436.4]
  wire  output_17_16; // @[Switch.scala 41:38:@7437.4]
  wire  _T_17672; // @[Switch.scala 41:52:@7439.4]
  wire  output_17_17; // @[Switch.scala 41:38:@7440.4]
  wire  _T_17675; // @[Switch.scala 41:52:@7442.4]
  wire  output_17_18; // @[Switch.scala 41:38:@7443.4]
  wire  _T_17678; // @[Switch.scala 41:52:@7445.4]
  wire  output_17_19; // @[Switch.scala 41:38:@7446.4]
  wire  _T_17681; // @[Switch.scala 41:52:@7448.4]
  wire  output_17_20; // @[Switch.scala 41:38:@7449.4]
  wire  _T_17684; // @[Switch.scala 41:52:@7451.4]
  wire  output_17_21; // @[Switch.scala 41:38:@7452.4]
  wire  _T_17687; // @[Switch.scala 41:52:@7454.4]
  wire  output_17_22; // @[Switch.scala 41:38:@7455.4]
  wire  _T_17690; // @[Switch.scala 41:52:@7457.4]
  wire  output_17_23; // @[Switch.scala 41:38:@7458.4]
  wire  _T_17693; // @[Switch.scala 41:52:@7460.4]
  wire  output_17_24; // @[Switch.scala 41:38:@7461.4]
  wire  _T_17696; // @[Switch.scala 41:52:@7463.4]
  wire  output_17_25; // @[Switch.scala 41:38:@7464.4]
  wire  _T_17699; // @[Switch.scala 41:52:@7466.4]
  wire  output_17_26; // @[Switch.scala 41:38:@7467.4]
  wire  _T_17702; // @[Switch.scala 41:52:@7469.4]
  wire  output_17_27; // @[Switch.scala 41:38:@7470.4]
  wire  _T_17705; // @[Switch.scala 41:52:@7472.4]
  wire  output_17_28; // @[Switch.scala 41:38:@7473.4]
  wire  _T_17708; // @[Switch.scala 41:52:@7475.4]
  wire  output_17_29; // @[Switch.scala 41:38:@7476.4]
  wire  _T_17711; // @[Switch.scala 41:52:@7478.4]
  wire  output_17_30; // @[Switch.scala 41:38:@7479.4]
  wire  _T_17714; // @[Switch.scala 41:52:@7481.4]
  wire  output_17_31; // @[Switch.scala 41:38:@7482.4]
  wire [7:0] _T_17722; // @[Switch.scala 43:31:@7490.4]
  wire [15:0] _T_17730; // @[Switch.scala 43:31:@7498.4]
  wire [7:0] _T_17737; // @[Switch.scala 43:31:@7505.4]
  wire [31:0] _T_17746; // @[Switch.scala 43:31:@7514.4]
  wire  _T_17750; // @[Switch.scala 41:52:@7517.4]
  wire  output_18_0; // @[Switch.scala 41:38:@7518.4]
  wire  _T_17753; // @[Switch.scala 41:52:@7520.4]
  wire  output_18_1; // @[Switch.scala 41:38:@7521.4]
  wire  _T_17756; // @[Switch.scala 41:52:@7523.4]
  wire  output_18_2; // @[Switch.scala 41:38:@7524.4]
  wire  _T_17759; // @[Switch.scala 41:52:@7526.4]
  wire  output_18_3; // @[Switch.scala 41:38:@7527.4]
  wire  _T_17762; // @[Switch.scala 41:52:@7529.4]
  wire  output_18_4; // @[Switch.scala 41:38:@7530.4]
  wire  _T_17765; // @[Switch.scala 41:52:@7532.4]
  wire  output_18_5; // @[Switch.scala 41:38:@7533.4]
  wire  _T_17768; // @[Switch.scala 41:52:@7535.4]
  wire  output_18_6; // @[Switch.scala 41:38:@7536.4]
  wire  _T_17771; // @[Switch.scala 41:52:@7538.4]
  wire  output_18_7; // @[Switch.scala 41:38:@7539.4]
  wire  _T_17774; // @[Switch.scala 41:52:@7541.4]
  wire  output_18_8; // @[Switch.scala 41:38:@7542.4]
  wire  _T_17777; // @[Switch.scala 41:52:@7544.4]
  wire  output_18_9; // @[Switch.scala 41:38:@7545.4]
  wire  _T_17780; // @[Switch.scala 41:52:@7547.4]
  wire  output_18_10; // @[Switch.scala 41:38:@7548.4]
  wire  _T_17783; // @[Switch.scala 41:52:@7550.4]
  wire  output_18_11; // @[Switch.scala 41:38:@7551.4]
  wire  _T_17786; // @[Switch.scala 41:52:@7553.4]
  wire  output_18_12; // @[Switch.scala 41:38:@7554.4]
  wire  _T_17789; // @[Switch.scala 41:52:@7556.4]
  wire  output_18_13; // @[Switch.scala 41:38:@7557.4]
  wire  _T_17792; // @[Switch.scala 41:52:@7559.4]
  wire  output_18_14; // @[Switch.scala 41:38:@7560.4]
  wire  _T_17795; // @[Switch.scala 41:52:@7562.4]
  wire  output_18_15; // @[Switch.scala 41:38:@7563.4]
  wire  _T_17798; // @[Switch.scala 41:52:@7565.4]
  wire  output_18_16; // @[Switch.scala 41:38:@7566.4]
  wire  _T_17801; // @[Switch.scala 41:52:@7568.4]
  wire  output_18_17; // @[Switch.scala 41:38:@7569.4]
  wire  _T_17804; // @[Switch.scala 41:52:@7571.4]
  wire  output_18_18; // @[Switch.scala 41:38:@7572.4]
  wire  _T_17807; // @[Switch.scala 41:52:@7574.4]
  wire  output_18_19; // @[Switch.scala 41:38:@7575.4]
  wire  _T_17810; // @[Switch.scala 41:52:@7577.4]
  wire  output_18_20; // @[Switch.scala 41:38:@7578.4]
  wire  _T_17813; // @[Switch.scala 41:52:@7580.4]
  wire  output_18_21; // @[Switch.scala 41:38:@7581.4]
  wire  _T_17816; // @[Switch.scala 41:52:@7583.4]
  wire  output_18_22; // @[Switch.scala 41:38:@7584.4]
  wire  _T_17819; // @[Switch.scala 41:52:@7586.4]
  wire  output_18_23; // @[Switch.scala 41:38:@7587.4]
  wire  _T_17822; // @[Switch.scala 41:52:@7589.4]
  wire  output_18_24; // @[Switch.scala 41:38:@7590.4]
  wire  _T_17825; // @[Switch.scala 41:52:@7592.4]
  wire  output_18_25; // @[Switch.scala 41:38:@7593.4]
  wire  _T_17828; // @[Switch.scala 41:52:@7595.4]
  wire  output_18_26; // @[Switch.scala 41:38:@7596.4]
  wire  _T_17831; // @[Switch.scala 41:52:@7598.4]
  wire  output_18_27; // @[Switch.scala 41:38:@7599.4]
  wire  _T_17834; // @[Switch.scala 41:52:@7601.4]
  wire  output_18_28; // @[Switch.scala 41:38:@7602.4]
  wire  _T_17837; // @[Switch.scala 41:52:@7604.4]
  wire  output_18_29; // @[Switch.scala 41:38:@7605.4]
  wire  _T_17840; // @[Switch.scala 41:52:@7607.4]
  wire  output_18_30; // @[Switch.scala 41:38:@7608.4]
  wire  _T_17843; // @[Switch.scala 41:52:@7610.4]
  wire  output_18_31; // @[Switch.scala 41:38:@7611.4]
  wire [7:0] _T_17851; // @[Switch.scala 43:31:@7619.4]
  wire [15:0] _T_17859; // @[Switch.scala 43:31:@7627.4]
  wire [7:0] _T_17866; // @[Switch.scala 43:31:@7634.4]
  wire [31:0] _T_17875; // @[Switch.scala 43:31:@7643.4]
  wire  _T_17879; // @[Switch.scala 41:52:@7646.4]
  wire  output_19_0; // @[Switch.scala 41:38:@7647.4]
  wire  _T_17882; // @[Switch.scala 41:52:@7649.4]
  wire  output_19_1; // @[Switch.scala 41:38:@7650.4]
  wire  _T_17885; // @[Switch.scala 41:52:@7652.4]
  wire  output_19_2; // @[Switch.scala 41:38:@7653.4]
  wire  _T_17888; // @[Switch.scala 41:52:@7655.4]
  wire  output_19_3; // @[Switch.scala 41:38:@7656.4]
  wire  _T_17891; // @[Switch.scala 41:52:@7658.4]
  wire  output_19_4; // @[Switch.scala 41:38:@7659.4]
  wire  _T_17894; // @[Switch.scala 41:52:@7661.4]
  wire  output_19_5; // @[Switch.scala 41:38:@7662.4]
  wire  _T_17897; // @[Switch.scala 41:52:@7664.4]
  wire  output_19_6; // @[Switch.scala 41:38:@7665.4]
  wire  _T_17900; // @[Switch.scala 41:52:@7667.4]
  wire  output_19_7; // @[Switch.scala 41:38:@7668.4]
  wire  _T_17903; // @[Switch.scala 41:52:@7670.4]
  wire  output_19_8; // @[Switch.scala 41:38:@7671.4]
  wire  _T_17906; // @[Switch.scala 41:52:@7673.4]
  wire  output_19_9; // @[Switch.scala 41:38:@7674.4]
  wire  _T_17909; // @[Switch.scala 41:52:@7676.4]
  wire  output_19_10; // @[Switch.scala 41:38:@7677.4]
  wire  _T_17912; // @[Switch.scala 41:52:@7679.4]
  wire  output_19_11; // @[Switch.scala 41:38:@7680.4]
  wire  _T_17915; // @[Switch.scala 41:52:@7682.4]
  wire  output_19_12; // @[Switch.scala 41:38:@7683.4]
  wire  _T_17918; // @[Switch.scala 41:52:@7685.4]
  wire  output_19_13; // @[Switch.scala 41:38:@7686.4]
  wire  _T_17921; // @[Switch.scala 41:52:@7688.4]
  wire  output_19_14; // @[Switch.scala 41:38:@7689.4]
  wire  _T_17924; // @[Switch.scala 41:52:@7691.4]
  wire  output_19_15; // @[Switch.scala 41:38:@7692.4]
  wire  _T_17927; // @[Switch.scala 41:52:@7694.4]
  wire  output_19_16; // @[Switch.scala 41:38:@7695.4]
  wire  _T_17930; // @[Switch.scala 41:52:@7697.4]
  wire  output_19_17; // @[Switch.scala 41:38:@7698.4]
  wire  _T_17933; // @[Switch.scala 41:52:@7700.4]
  wire  output_19_18; // @[Switch.scala 41:38:@7701.4]
  wire  _T_17936; // @[Switch.scala 41:52:@7703.4]
  wire  output_19_19; // @[Switch.scala 41:38:@7704.4]
  wire  _T_17939; // @[Switch.scala 41:52:@7706.4]
  wire  output_19_20; // @[Switch.scala 41:38:@7707.4]
  wire  _T_17942; // @[Switch.scala 41:52:@7709.4]
  wire  output_19_21; // @[Switch.scala 41:38:@7710.4]
  wire  _T_17945; // @[Switch.scala 41:52:@7712.4]
  wire  output_19_22; // @[Switch.scala 41:38:@7713.4]
  wire  _T_17948; // @[Switch.scala 41:52:@7715.4]
  wire  output_19_23; // @[Switch.scala 41:38:@7716.4]
  wire  _T_17951; // @[Switch.scala 41:52:@7718.4]
  wire  output_19_24; // @[Switch.scala 41:38:@7719.4]
  wire  _T_17954; // @[Switch.scala 41:52:@7721.4]
  wire  output_19_25; // @[Switch.scala 41:38:@7722.4]
  wire  _T_17957; // @[Switch.scala 41:52:@7724.4]
  wire  output_19_26; // @[Switch.scala 41:38:@7725.4]
  wire  _T_17960; // @[Switch.scala 41:52:@7727.4]
  wire  output_19_27; // @[Switch.scala 41:38:@7728.4]
  wire  _T_17963; // @[Switch.scala 41:52:@7730.4]
  wire  output_19_28; // @[Switch.scala 41:38:@7731.4]
  wire  _T_17966; // @[Switch.scala 41:52:@7733.4]
  wire  output_19_29; // @[Switch.scala 41:38:@7734.4]
  wire  _T_17969; // @[Switch.scala 41:52:@7736.4]
  wire  output_19_30; // @[Switch.scala 41:38:@7737.4]
  wire  _T_17972; // @[Switch.scala 41:52:@7739.4]
  wire  output_19_31; // @[Switch.scala 41:38:@7740.4]
  wire [7:0] _T_17980; // @[Switch.scala 43:31:@7748.4]
  wire [15:0] _T_17988; // @[Switch.scala 43:31:@7756.4]
  wire [7:0] _T_17995; // @[Switch.scala 43:31:@7763.4]
  wire [31:0] _T_18004; // @[Switch.scala 43:31:@7772.4]
  wire  _T_18008; // @[Switch.scala 41:52:@7775.4]
  wire  output_20_0; // @[Switch.scala 41:38:@7776.4]
  wire  _T_18011; // @[Switch.scala 41:52:@7778.4]
  wire  output_20_1; // @[Switch.scala 41:38:@7779.4]
  wire  _T_18014; // @[Switch.scala 41:52:@7781.4]
  wire  output_20_2; // @[Switch.scala 41:38:@7782.4]
  wire  _T_18017; // @[Switch.scala 41:52:@7784.4]
  wire  output_20_3; // @[Switch.scala 41:38:@7785.4]
  wire  _T_18020; // @[Switch.scala 41:52:@7787.4]
  wire  output_20_4; // @[Switch.scala 41:38:@7788.4]
  wire  _T_18023; // @[Switch.scala 41:52:@7790.4]
  wire  output_20_5; // @[Switch.scala 41:38:@7791.4]
  wire  _T_18026; // @[Switch.scala 41:52:@7793.4]
  wire  output_20_6; // @[Switch.scala 41:38:@7794.4]
  wire  _T_18029; // @[Switch.scala 41:52:@7796.4]
  wire  output_20_7; // @[Switch.scala 41:38:@7797.4]
  wire  _T_18032; // @[Switch.scala 41:52:@7799.4]
  wire  output_20_8; // @[Switch.scala 41:38:@7800.4]
  wire  _T_18035; // @[Switch.scala 41:52:@7802.4]
  wire  output_20_9; // @[Switch.scala 41:38:@7803.4]
  wire  _T_18038; // @[Switch.scala 41:52:@7805.4]
  wire  output_20_10; // @[Switch.scala 41:38:@7806.4]
  wire  _T_18041; // @[Switch.scala 41:52:@7808.4]
  wire  output_20_11; // @[Switch.scala 41:38:@7809.4]
  wire  _T_18044; // @[Switch.scala 41:52:@7811.4]
  wire  output_20_12; // @[Switch.scala 41:38:@7812.4]
  wire  _T_18047; // @[Switch.scala 41:52:@7814.4]
  wire  output_20_13; // @[Switch.scala 41:38:@7815.4]
  wire  _T_18050; // @[Switch.scala 41:52:@7817.4]
  wire  output_20_14; // @[Switch.scala 41:38:@7818.4]
  wire  _T_18053; // @[Switch.scala 41:52:@7820.4]
  wire  output_20_15; // @[Switch.scala 41:38:@7821.4]
  wire  _T_18056; // @[Switch.scala 41:52:@7823.4]
  wire  output_20_16; // @[Switch.scala 41:38:@7824.4]
  wire  _T_18059; // @[Switch.scala 41:52:@7826.4]
  wire  output_20_17; // @[Switch.scala 41:38:@7827.4]
  wire  _T_18062; // @[Switch.scala 41:52:@7829.4]
  wire  output_20_18; // @[Switch.scala 41:38:@7830.4]
  wire  _T_18065; // @[Switch.scala 41:52:@7832.4]
  wire  output_20_19; // @[Switch.scala 41:38:@7833.4]
  wire  _T_18068; // @[Switch.scala 41:52:@7835.4]
  wire  output_20_20; // @[Switch.scala 41:38:@7836.4]
  wire  _T_18071; // @[Switch.scala 41:52:@7838.4]
  wire  output_20_21; // @[Switch.scala 41:38:@7839.4]
  wire  _T_18074; // @[Switch.scala 41:52:@7841.4]
  wire  output_20_22; // @[Switch.scala 41:38:@7842.4]
  wire  _T_18077; // @[Switch.scala 41:52:@7844.4]
  wire  output_20_23; // @[Switch.scala 41:38:@7845.4]
  wire  _T_18080; // @[Switch.scala 41:52:@7847.4]
  wire  output_20_24; // @[Switch.scala 41:38:@7848.4]
  wire  _T_18083; // @[Switch.scala 41:52:@7850.4]
  wire  output_20_25; // @[Switch.scala 41:38:@7851.4]
  wire  _T_18086; // @[Switch.scala 41:52:@7853.4]
  wire  output_20_26; // @[Switch.scala 41:38:@7854.4]
  wire  _T_18089; // @[Switch.scala 41:52:@7856.4]
  wire  output_20_27; // @[Switch.scala 41:38:@7857.4]
  wire  _T_18092; // @[Switch.scala 41:52:@7859.4]
  wire  output_20_28; // @[Switch.scala 41:38:@7860.4]
  wire  _T_18095; // @[Switch.scala 41:52:@7862.4]
  wire  output_20_29; // @[Switch.scala 41:38:@7863.4]
  wire  _T_18098; // @[Switch.scala 41:52:@7865.4]
  wire  output_20_30; // @[Switch.scala 41:38:@7866.4]
  wire  _T_18101; // @[Switch.scala 41:52:@7868.4]
  wire  output_20_31; // @[Switch.scala 41:38:@7869.4]
  wire [7:0] _T_18109; // @[Switch.scala 43:31:@7877.4]
  wire [15:0] _T_18117; // @[Switch.scala 43:31:@7885.4]
  wire [7:0] _T_18124; // @[Switch.scala 43:31:@7892.4]
  wire [31:0] _T_18133; // @[Switch.scala 43:31:@7901.4]
  wire  _T_18137; // @[Switch.scala 41:52:@7904.4]
  wire  output_21_0; // @[Switch.scala 41:38:@7905.4]
  wire  _T_18140; // @[Switch.scala 41:52:@7907.4]
  wire  output_21_1; // @[Switch.scala 41:38:@7908.4]
  wire  _T_18143; // @[Switch.scala 41:52:@7910.4]
  wire  output_21_2; // @[Switch.scala 41:38:@7911.4]
  wire  _T_18146; // @[Switch.scala 41:52:@7913.4]
  wire  output_21_3; // @[Switch.scala 41:38:@7914.4]
  wire  _T_18149; // @[Switch.scala 41:52:@7916.4]
  wire  output_21_4; // @[Switch.scala 41:38:@7917.4]
  wire  _T_18152; // @[Switch.scala 41:52:@7919.4]
  wire  output_21_5; // @[Switch.scala 41:38:@7920.4]
  wire  _T_18155; // @[Switch.scala 41:52:@7922.4]
  wire  output_21_6; // @[Switch.scala 41:38:@7923.4]
  wire  _T_18158; // @[Switch.scala 41:52:@7925.4]
  wire  output_21_7; // @[Switch.scala 41:38:@7926.4]
  wire  _T_18161; // @[Switch.scala 41:52:@7928.4]
  wire  output_21_8; // @[Switch.scala 41:38:@7929.4]
  wire  _T_18164; // @[Switch.scala 41:52:@7931.4]
  wire  output_21_9; // @[Switch.scala 41:38:@7932.4]
  wire  _T_18167; // @[Switch.scala 41:52:@7934.4]
  wire  output_21_10; // @[Switch.scala 41:38:@7935.4]
  wire  _T_18170; // @[Switch.scala 41:52:@7937.4]
  wire  output_21_11; // @[Switch.scala 41:38:@7938.4]
  wire  _T_18173; // @[Switch.scala 41:52:@7940.4]
  wire  output_21_12; // @[Switch.scala 41:38:@7941.4]
  wire  _T_18176; // @[Switch.scala 41:52:@7943.4]
  wire  output_21_13; // @[Switch.scala 41:38:@7944.4]
  wire  _T_18179; // @[Switch.scala 41:52:@7946.4]
  wire  output_21_14; // @[Switch.scala 41:38:@7947.4]
  wire  _T_18182; // @[Switch.scala 41:52:@7949.4]
  wire  output_21_15; // @[Switch.scala 41:38:@7950.4]
  wire  _T_18185; // @[Switch.scala 41:52:@7952.4]
  wire  output_21_16; // @[Switch.scala 41:38:@7953.4]
  wire  _T_18188; // @[Switch.scala 41:52:@7955.4]
  wire  output_21_17; // @[Switch.scala 41:38:@7956.4]
  wire  _T_18191; // @[Switch.scala 41:52:@7958.4]
  wire  output_21_18; // @[Switch.scala 41:38:@7959.4]
  wire  _T_18194; // @[Switch.scala 41:52:@7961.4]
  wire  output_21_19; // @[Switch.scala 41:38:@7962.4]
  wire  _T_18197; // @[Switch.scala 41:52:@7964.4]
  wire  output_21_20; // @[Switch.scala 41:38:@7965.4]
  wire  _T_18200; // @[Switch.scala 41:52:@7967.4]
  wire  output_21_21; // @[Switch.scala 41:38:@7968.4]
  wire  _T_18203; // @[Switch.scala 41:52:@7970.4]
  wire  output_21_22; // @[Switch.scala 41:38:@7971.4]
  wire  _T_18206; // @[Switch.scala 41:52:@7973.4]
  wire  output_21_23; // @[Switch.scala 41:38:@7974.4]
  wire  _T_18209; // @[Switch.scala 41:52:@7976.4]
  wire  output_21_24; // @[Switch.scala 41:38:@7977.4]
  wire  _T_18212; // @[Switch.scala 41:52:@7979.4]
  wire  output_21_25; // @[Switch.scala 41:38:@7980.4]
  wire  _T_18215; // @[Switch.scala 41:52:@7982.4]
  wire  output_21_26; // @[Switch.scala 41:38:@7983.4]
  wire  _T_18218; // @[Switch.scala 41:52:@7985.4]
  wire  output_21_27; // @[Switch.scala 41:38:@7986.4]
  wire  _T_18221; // @[Switch.scala 41:52:@7988.4]
  wire  output_21_28; // @[Switch.scala 41:38:@7989.4]
  wire  _T_18224; // @[Switch.scala 41:52:@7991.4]
  wire  output_21_29; // @[Switch.scala 41:38:@7992.4]
  wire  _T_18227; // @[Switch.scala 41:52:@7994.4]
  wire  output_21_30; // @[Switch.scala 41:38:@7995.4]
  wire  _T_18230; // @[Switch.scala 41:52:@7997.4]
  wire  output_21_31; // @[Switch.scala 41:38:@7998.4]
  wire [7:0] _T_18238; // @[Switch.scala 43:31:@8006.4]
  wire [15:0] _T_18246; // @[Switch.scala 43:31:@8014.4]
  wire [7:0] _T_18253; // @[Switch.scala 43:31:@8021.4]
  wire [31:0] _T_18262; // @[Switch.scala 43:31:@8030.4]
  wire  _T_18266; // @[Switch.scala 41:52:@8033.4]
  wire  output_22_0; // @[Switch.scala 41:38:@8034.4]
  wire  _T_18269; // @[Switch.scala 41:52:@8036.4]
  wire  output_22_1; // @[Switch.scala 41:38:@8037.4]
  wire  _T_18272; // @[Switch.scala 41:52:@8039.4]
  wire  output_22_2; // @[Switch.scala 41:38:@8040.4]
  wire  _T_18275; // @[Switch.scala 41:52:@8042.4]
  wire  output_22_3; // @[Switch.scala 41:38:@8043.4]
  wire  _T_18278; // @[Switch.scala 41:52:@8045.4]
  wire  output_22_4; // @[Switch.scala 41:38:@8046.4]
  wire  _T_18281; // @[Switch.scala 41:52:@8048.4]
  wire  output_22_5; // @[Switch.scala 41:38:@8049.4]
  wire  _T_18284; // @[Switch.scala 41:52:@8051.4]
  wire  output_22_6; // @[Switch.scala 41:38:@8052.4]
  wire  _T_18287; // @[Switch.scala 41:52:@8054.4]
  wire  output_22_7; // @[Switch.scala 41:38:@8055.4]
  wire  _T_18290; // @[Switch.scala 41:52:@8057.4]
  wire  output_22_8; // @[Switch.scala 41:38:@8058.4]
  wire  _T_18293; // @[Switch.scala 41:52:@8060.4]
  wire  output_22_9; // @[Switch.scala 41:38:@8061.4]
  wire  _T_18296; // @[Switch.scala 41:52:@8063.4]
  wire  output_22_10; // @[Switch.scala 41:38:@8064.4]
  wire  _T_18299; // @[Switch.scala 41:52:@8066.4]
  wire  output_22_11; // @[Switch.scala 41:38:@8067.4]
  wire  _T_18302; // @[Switch.scala 41:52:@8069.4]
  wire  output_22_12; // @[Switch.scala 41:38:@8070.4]
  wire  _T_18305; // @[Switch.scala 41:52:@8072.4]
  wire  output_22_13; // @[Switch.scala 41:38:@8073.4]
  wire  _T_18308; // @[Switch.scala 41:52:@8075.4]
  wire  output_22_14; // @[Switch.scala 41:38:@8076.4]
  wire  _T_18311; // @[Switch.scala 41:52:@8078.4]
  wire  output_22_15; // @[Switch.scala 41:38:@8079.4]
  wire  _T_18314; // @[Switch.scala 41:52:@8081.4]
  wire  output_22_16; // @[Switch.scala 41:38:@8082.4]
  wire  _T_18317; // @[Switch.scala 41:52:@8084.4]
  wire  output_22_17; // @[Switch.scala 41:38:@8085.4]
  wire  _T_18320; // @[Switch.scala 41:52:@8087.4]
  wire  output_22_18; // @[Switch.scala 41:38:@8088.4]
  wire  _T_18323; // @[Switch.scala 41:52:@8090.4]
  wire  output_22_19; // @[Switch.scala 41:38:@8091.4]
  wire  _T_18326; // @[Switch.scala 41:52:@8093.4]
  wire  output_22_20; // @[Switch.scala 41:38:@8094.4]
  wire  _T_18329; // @[Switch.scala 41:52:@8096.4]
  wire  output_22_21; // @[Switch.scala 41:38:@8097.4]
  wire  _T_18332; // @[Switch.scala 41:52:@8099.4]
  wire  output_22_22; // @[Switch.scala 41:38:@8100.4]
  wire  _T_18335; // @[Switch.scala 41:52:@8102.4]
  wire  output_22_23; // @[Switch.scala 41:38:@8103.4]
  wire  _T_18338; // @[Switch.scala 41:52:@8105.4]
  wire  output_22_24; // @[Switch.scala 41:38:@8106.4]
  wire  _T_18341; // @[Switch.scala 41:52:@8108.4]
  wire  output_22_25; // @[Switch.scala 41:38:@8109.4]
  wire  _T_18344; // @[Switch.scala 41:52:@8111.4]
  wire  output_22_26; // @[Switch.scala 41:38:@8112.4]
  wire  _T_18347; // @[Switch.scala 41:52:@8114.4]
  wire  output_22_27; // @[Switch.scala 41:38:@8115.4]
  wire  _T_18350; // @[Switch.scala 41:52:@8117.4]
  wire  output_22_28; // @[Switch.scala 41:38:@8118.4]
  wire  _T_18353; // @[Switch.scala 41:52:@8120.4]
  wire  output_22_29; // @[Switch.scala 41:38:@8121.4]
  wire  _T_18356; // @[Switch.scala 41:52:@8123.4]
  wire  output_22_30; // @[Switch.scala 41:38:@8124.4]
  wire  _T_18359; // @[Switch.scala 41:52:@8126.4]
  wire  output_22_31; // @[Switch.scala 41:38:@8127.4]
  wire [7:0] _T_18367; // @[Switch.scala 43:31:@8135.4]
  wire [15:0] _T_18375; // @[Switch.scala 43:31:@8143.4]
  wire [7:0] _T_18382; // @[Switch.scala 43:31:@8150.4]
  wire [31:0] _T_18391; // @[Switch.scala 43:31:@8159.4]
  wire  _T_18395; // @[Switch.scala 41:52:@8162.4]
  wire  output_23_0; // @[Switch.scala 41:38:@8163.4]
  wire  _T_18398; // @[Switch.scala 41:52:@8165.4]
  wire  output_23_1; // @[Switch.scala 41:38:@8166.4]
  wire  _T_18401; // @[Switch.scala 41:52:@8168.4]
  wire  output_23_2; // @[Switch.scala 41:38:@8169.4]
  wire  _T_18404; // @[Switch.scala 41:52:@8171.4]
  wire  output_23_3; // @[Switch.scala 41:38:@8172.4]
  wire  _T_18407; // @[Switch.scala 41:52:@8174.4]
  wire  output_23_4; // @[Switch.scala 41:38:@8175.4]
  wire  _T_18410; // @[Switch.scala 41:52:@8177.4]
  wire  output_23_5; // @[Switch.scala 41:38:@8178.4]
  wire  _T_18413; // @[Switch.scala 41:52:@8180.4]
  wire  output_23_6; // @[Switch.scala 41:38:@8181.4]
  wire  _T_18416; // @[Switch.scala 41:52:@8183.4]
  wire  output_23_7; // @[Switch.scala 41:38:@8184.4]
  wire  _T_18419; // @[Switch.scala 41:52:@8186.4]
  wire  output_23_8; // @[Switch.scala 41:38:@8187.4]
  wire  _T_18422; // @[Switch.scala 41:52:@8189.4]
  wire  output_23_9; // @[Switch.scala 41:38:@8190.4]
  wire  _T_18425; // @[Switch.scala 41:52:@8192.4]
  wire  output_23_10; // @[Switch.scala 41:38:@8193.4]
  wire  _T_18428; // @[Switch.scala 41:52:@8195.4]
  wire  output_23_11; // @[Switch.scala 41:38:@8196.4]
  wire  _T_18431; // @[Switch.scala 41:52:@8198.4]
  wire  output_23_12; // @[Switch.scala 41:38:@8199.4]
  wire  _T_18434; // @[Switch.scala 41:52:@8201.4]
  wire  output_23_13; // @[Switch.scala 41:38:@8202.4]
  wire  _T_18437; // @[Switch.scala 41:52:@8204.4]
  wire  output_23_14; // @[Switch.scala 41:38:@8205.4]
  wire  _T_18440; // @[Switch.scala 41:52:@8207.4]
  wire  output_23_15; // @[Switch.scala 41:38:@8208.4]
  wire  _T_18443; // @[Switch.scala 41:52:@8210.4]
  wire  output_23_16; // @[Switch.scala 41:38:@8211.4]
  wire  _T_18446; // @[Switch.scala 41:52:@8213.4]
  wire  output_23_17; // @[Switch.scala 41:38:@8214.4]
  wire  _T_18449; // @[Switch.scala 41:52:@8216.4]
  wire  output_23_18; // @[Switch.scala 41:38:@8217.4]
  wire  _T_18452; // @[Switch.scala 41:52:@8219.4]
  wire  output_23_19; // @[Switch.scala 41:38:@8220.4]
  wire  _T_18455; // @[Switch.scala 41:52:@8222.4]
  wire  output_23_20; // @[Switch.scala 41:38:@8223.4]
  wire  _T_18458; // @[Switch.scala 41:52:@8225.4]
  wire  output_23_21; // @[Switch.scala 41:38:@8226.4]
  wire  _T_18461; // @[Switch.scala 41:52:@8228.4]
  wire  output_23_22; // @[Switch.scala 41:38:@8229.4]
  wire  _T_18464; // @[Switch.scala 41:52:@8231.4]
  wire  output_23_23; // @[Switch.scala 41:38:@8232.4]
  wire  _T_18467; // @[Switch.scala 41:52:@8234.4]
  wire  output_23_24; // @[Switch.scala 41:38:@8235.4]
  wire  _T_18470; // @[Switch.scala 41:52:@8237.4]
  wire  output_23_25; // @[Switch.scala 41:38:@8238.4]
  wire  _T_18473; // @[Switch.scala 41:52:@8240.4]
  wire  output_23_26; // @[Switch.scala 41:38:@8241.4]
  wire  _T_18476; // @[Switch.scala 41:52:@8243.4]
  wire  output_23_27; // @[Switch.scala 41:38:@8244.4]
  wire  _T_18479; // @[Switch.scala 41:52:@8246.4]
  wire  output_23_28; // @[Switch.scala 41:38:@8247.4]
  wire  _T_18482; // @[Switch.scala 41:52:@8249.4]
  wire  output_23_29; // @[Switch.scala 41:38:@8250.4]
  wire  _T_18485; // @[Switch.scala 41:52:@8252.4]
  wire  output_23_30; // @[Switch.scala 41:38:@8253.4]
  wire  _T_18488; // @[Switch.scala 41:52:@8255.4]
  wire  output_23_31; // @[Switch.scala 41:38:@8256.4]
  wire [7:0] _T_18496; // @[Switch.scala 43:31:@8264.4]
  wire [15:0] _T_18504; // @[Switch.scala 43:31:@8272.4]
  wire [7:0] _T_18511; // @[Switch.scala 43:31:@8279.4]
  wire [31:0] _T_18520; // @[Switch.scala 43:31:@8288.4]
  wire  _T_18524; // @[Switch.scala 41:52:@8291.4]
  wire  output_24_0; // @[Switch.scala 41:38:@8292.4]
  wire  _T_18527; // @[Switch.scala 41:52:@8294.4]
  wire  output_24_1; // @[Switch.scala 41:38:@8295.4]
  wire  _T_18530; // @[Switch.scala 41:52:@8297.4]
  wire  output_24_2; // @[Switch.scala 41:38:@8298.4]
  wire  _T_18533; // @[Switch.scala 41:52:@8300.4]
  wire  output_24_3; // @[Switch.scala 41:38:@8301.4]
  wire  _T_18536; // @[Switch.scala 41:52:@8303.4]
  wire  output_24_4; // @[Switch.scala 41:38:@8304.4]
  wire  _T_18539; // @[Switch.scala 41:52:@8306.4]
  wire  output_24_5; // @[Switch.scala 41:38:@8307.4]
  wire  _T_18542; // @[Switch.scala 41:52:@8309.4]
  wire  output_24_6; // @[Switch.scala 41:38:@8310.4]
  wire  _T_18545; // @[Switch.scala 41:52:@8312.4]
  wire  output_24_7; // @[Switch.scala 41:38:@8313.4]
  wire  _T_18548; // @[Switch.scala 41:52:@8315.4]
  wire  output_24_8; // @[Switch.scala 41:38:@8316.4]
  wire  _T_18551; // @[Switch.scala 41:52:@8318.4]
  wire  output_24_9; // @[Switch.scala 41:38:@8319.4]
  wire  _T_18554; // @[Switch.scala 41:52:@8321.4]
  wire  output_24_10; // @[Switch.scala 41:38:@8322.4]
  wire  _T_18557; // @[Switch.scala 41:52:@8324.4]
  wire  output_24_11; // @[Switch.scala 41:38:@8325.4]
  wire  _T_18560; // @[Switch.scala 41:52:@8327.4]
  wire  output_24_12; // @[Switch.scala 41:38:@8328.4]
  wire  _T_18563; // @[Switch.scala 41:52:@8330.4]
  wire  output_24_13; // @[Switch.scala 41:38:@8331.4]
  wire  _T_18566; // @[Switch.scala 41:52:@8333.4]
  wire  output_24_14; // @[Switch.scala 41:38:@8334.4]
  wire  _T_18569; // @[Switch.scala 41:52:@8336.4]
  wire  output_24_15; // @[Switch.scala 41:38:@8337.4]
  wire  _T_18572; // @[Switch.scala 41:52:@8339.4]
  wire  output_24_16; // @[Switch.scala 41:38:@8340.4]
  wire  _T_18575; // @[Switch.scala 41:52:@8342.4]
  wire  output_24_17; // @[Switch.scala 41:38:@8343.4]
  wire  _T_18578; // @[Switch.scala 41:52:@8345.4]
  wire  output_24_18; // @[Switch.scala 41:38:@8346.4]
  wire  _T_18581; // @[Switch.scala 41:52:@8348.4]
  wire  output_24_19; // @[Switch.scala 41:38:@8349.4]
  wire  _T_18584; // @[Switch.scala 41:52:@8351.4]
  wire  output_24_20; // @[Switch.scala 41:38:@8352.4]
  wire  _T_18587; // @[Switch.scala 41:52:@8354.4]
  wire  output_24_21; // @[Switch.scala 41:38:@8355.4]
  wire  _T_18590; // @[Switch.scala 41:52:@8357.4]
  wire  output_24_22; // @[Switch.scala 41:38:@8358.4]
  wire  _T_18593; // @[Switch.scala 41:52:@8360.4]
  wire  output_24_23; // @[Switch.scala 41:38:@8361.4]
  wire  _T_18596; // @[Switch.scala 41:52:@8363.4]
  wire  output_24_24; // @[Switch.scala 41:38:@8364.4]
  wire  _T_18599; // @[Switch.scala 41:52:@8366.4]
  wire  output_24_25; // @[Switch.scala 41:38:@8367.4]
  wire  _T_18602; // @[Switch.scala 41:52:@8369.4]
  wire  output_24_26; // @[Switch.scala 41:38:@8370.4]
  wire  _T_18605; // @[Switch.scala 41:52:@8372.4]
  wire  output_24_27; // @[Switch.scala 41:38:@8373.4]
  wire  _T_18608; // @[Switch.scala 41:52:@8375.4]
  wire  output_24_28; // @[Switch.scala 41:38:@8376.4]
  wire  _T_18611; // @[Switch.scala 41:52:@8378.4]
  wire  output_24_29; // @[Switch.scala 41:38:@8379.4]
  wire  _T_18614; // @[Switch.scala 41:52:@8381.4]
  wire  output_24_30; // @[Switch.scala 41:38:@8382.4]
  wire  _T_18617; // @[Switch.scala 41:52:@8384.4]
  wire  output_24_31; // @[Switch.scala 41:38:@8385.4]
  wire [7:0] _T_18625; // @[Switch.scala 43:31:@8393.4]
  wire [15:0] _T_18633; // @[Switch.scala 43:31:@8401.4]
  wire [7:0] _T_18640; // @[Switch.scala 43:31:@8408.4]
  wire [31:0] _T_18649; // @[Switch.scala 43:31:@8417.4]
  wire  _T_18653; // @[Switch.scala 41:52:@8420.4]
  wire  output_25_0; // @[Switch.scala 41:38:@8421.4]
  wire  _T_18656; // @[Switch.scala 41:52:@8423.4]
  wire  output_25_1; // @[Switch.scala 41:38:@8424.4]
  wire  _T_18659; // @[Switch.scala 41:52:@8426.4]
  wire  output_25_2; // @[Switch.scala 41:38:@8427.4]
  wire  _T_18662; // @[Switch.scala 41:52:@8429.4]
  wire  output_25_3; // @[Switch.scala 41:38:@8430.4]
  wire  _T_18665; // @[Switch.scala 41:52:@8432.4]
  wire  output_25_4; // @[Switch.scala 41:38:@8433.4]
  wire  _T_18668; // @[Switch.scala 41:52:@8435.4]
  wire  output_25_5; // @[Switch.scala 41:38:@8436.4]
  wire  _T_18671; // @[Switch.scala 41:52:@8438.4]
  wire  output_25_6; // @[Switch.scala 41:38:@8439.4]
  wire  _T_18674; // @[Switch.scala 41:52:@8441.4]
  wire  output_25_7; // @[Switch.scala 41:38:@8442.4]
  wire  _T_18677; // @[Switch.scala 41:52:@8444.4]
  wire  output_25_8; // @[Switch.scala 41:38:@8445.4]
  wire  _T_18680; // @[Switch.scala 41:52:@8447.4]
  wire  output_25_9; // @[Switch.scala 41:38:@8448.4]
  wire  _T_18683; // @[Switch.scala 41:52:@8450.4]
  wire  output_25_10; // @[Switch.scala 41:38:@8451.4]
  wire  _T_18686; // @[Switch.scala 41:52:@8453.4]
  wire  output_25_11; // @[Switch.scala 41:38:@8454.4]
  wire  _T_18689; // @[Switch.scala 41:52:@8456.4]
  wire  output_25_12; // @[Switch.scala 41:38:@8457.4]
  wire  _T_18692; // @[Switch.scala 41:52:@8459.4]
  wire  output_25_13; // @[Switch.scala 41:38:@8460.4]
  wire  _T_18695; // @[Switch.scala 41:52:@8462.4]
  wire  output_25_14; // @[Switch.scala 41:38:@8463.4]
  wire  _T_18698; // @[Switch.scala 41:52:@8465.4]
  wire  output_25_15; // @[Switch.scala 41:38:@8466.4]
  wire  _T_18701; // @[Switch.scala 41:52:@8468.4]
  wire  output_25_16; // @[Switch.scala 41:38:@8469.4]
  wire  _T_18704; // @[Switch.scala 41:52:@8471.4]
  wire  output_25_17; // @[Switch.scala 41:38:@8472.4]
  wire  _T_18707; // @[Switch.scala 41:52:@8474.4]
  wire  output_25_18; // @[Switch.scala 41:38:@8475.4]
  wire  _T_18710; // @[Switch.scala 41:52:@8477.4]
  wire  output_25_19; // @[Switch.scala 41:38:@8478.4]
  wire  _T_18713; // @[Switch.scala 41:52:@8480.4]
  wire  output_25_20; // @[Switch.scala 41:38:@8481.4]
  wire  _T_18716; // @[Switch.scala 41:52:@8483.4]
  wire  output_25_21; // @[Switch.scala 41:38:@8484.4]
  wire  _T_18719; // @[Switch.scala 41:52:@8486.4]
  wire  output_25_22; // @[Switch.scala 41:38:@8487.4]
  wire  _T_18722; // @[Switch.scala 41:52:@8489.4]
  wire  output_25_23; // @[Switch.scala 41:38:@8490.4]
  wire  _T_18725; // @[Switch.scala 41:52:@8492.4]
  wire  output_25_24; // @[Switch.scala 41:38:@8493.4]
  wire  _T_18728; // @[Switch.scala 41:52:@8495.4]
  wire  output_25_25; // @[Switch.scala 41:38:@8496.4]
  wire  _T_18731; // @[Switch.scala 41:52:@8498.4]
  wire  output_25_26; // @[Switch.scala 41:38:@8499.4]
  wire  _T_18734; // @[Switch.scala 41:52:@8501.4]
  wire  output_25_27; // @[Switch.scala 41:38:@8502.4]
  wire  _T_18737; // @[Switch.scala 41:52:@8504.4]
  wire  output_25_28; // @[Switch.scala 41:38:@8505.4]
  wire  _T_18740; // @[Switch.scala 41:52:@8507.4]
  wire  output_25_29; // @[Switch.scala 41:38:@8508.4]
  wire  _T_18743; // @[Switch.scala 41:52:@8510.4]
  wire  output_25_30; // @[Switch.scala 41:38:@8511.4]
  wire  _T_18746; // @[Switch.scala 41:52:@8513.4]
  wire  output_25_31; // @[Switch.scala 41:38:@8514.4]
  wire [7:0] _T_18754; // @[Switch.scala 43:31:@8522.4]
  wire [15:0] _T_18762; // @[Switch.scala 43:31:@8530.4]
  wire [7:0] _T_18769; // @[Switch.scala 43:31:@8537.4]
  wire [31:0] _T_18778; // @[Switch.scala 43:31:@8546.4]
  wire  _T_18782; // @[Switch.scala 41:52:@8549.4]
  wire  output_26_0; // @[Switch.scala 41:38:@8550.4]
  wire  _T_18785; // @[Switch.scala 41:52:@8552.4]
  wire  output_26_1; // @[Switch.scala 41:38:@8553.4]
  wire  _T_18788; // @[Switch.scala 41:52:@8555.4]
  wire  output_26_2; // @[Switch.scala 41:38:@8556.4]
  wire  _T_18791; // @[Switch.scala 41:52:@8558.4]
  wire  output_26_3; // @[Switch.scala 41:38:@8559.4]
  wire  _T_18794; // @[Switch.scala 41:52:@8561.4]
  wire  output_26_4; // @[Switch.scala 41:38:@8562.4]
  wire  _T_18797; // @[Switch.scala 41:52:@8564.4]
  wire  output_26_5; // @[Switch.scala 41:38:@8565.4]
  wire  _T_18800; // @[Switch.scala 41:52:@8567.4]
  wire  output_26_6; // @[Switch.scala 41:38:@8568.4]
  wire  _T_18803; // @[Switch.scala 41:52:@8570.4]
  wire  output_26_7; // @[Switch.scala 41:38:@8571.4]
  wire  _T_18806; // @[Switch.scala 41:52:@8573.4]
  wire  output_26_8; // @[Switch.scala 41:38:@8574.4]
  wire  _T_18809; // @[Switch.scala 41:52:@8576.4]
  wire  output_26_9; // @[Switch.scala 41:38:@8577.4]
  wire  _T_18812; // @[Switch.scala 41:52:@8579.4]
  wire  output_26_10; // @[Switch.scala 41:38:@8580.4]
  wire  _T_18815; // @[Switch.scala 41:52:@8582.4]
  wire  output_26_11; // @[Switch.scala 41:38:@8583.4]
  wire  _T_18818; // @[Switch.scala 41:52:@8585.4]
  wire  output_26_12; // @[Switch.scala 41:38:@8586.4]
  wire  _T_18821; // @[Switch.scala 41:52:@8588.4]
  wire  output_26_13; // @[Switch.scala 41:38:@8589.4]
  wire  _T_18824; // @[Switch.scala 41:52:@8591.4]
  wire  output_26_14; // @[Switch.scala 41:38:@8592.4]
  wire  _T_18827; // @[Switch.scala 41:52:@8594.4]
  wire  output_26_15; // @[Switch.scala 41:38:@8595.4]
  wire  _T_18830; // @[Switch.scala 41:52:@8597.4]
  wire  output_26_16; // @[Switch.scala 41:38:@8598.4]
  wire  _T_18833; // @[Switch.scala 41:52:@8600.4]
  wire  output_26_17; // @[Switch.scala 41:38:@8601.4]
  wire  _T_18836; // @[Switch.scala 41:52:@8603.4]
  wire  output_26_18; // @[Switch.scala 41:38:@8604.4]
  wire  _T_18839; // @[Switch.scala 41:52:@8606.4]
  wire  output_26_19; // @[Switch.scala 41:38:@8607.4]
  wire  _T_18842; // @[Switch.scala 41:52:@8609.4]
  wire  output_26_20; // @[Switch.scala 41:38:@8610.4]
  wire  _T_18845; // @[Switch.scala 41:52:@8612.4]
  wire  output_26_21; // @[Switch.scala 41:38:@8613.4]
  wire  _T_18848; // @[Switch.scala 41:52:@8615.4]
  wire  output_26_22; // @[Switch.scala 41:38:@8616.4]
  wire  _T_18851; // @[Switch.scala 41:52:@8618.4]
  wire  output_26_23; // @[Switch.scala 41:38:@8619.4]
  wire  _T_18854; // @[Switch.scala 41:52:@8621.4]
  wire  output_26_24; // @[Switch.scala 41:38:@8622.4]
  wire  _T_18857; // @[Switch.scala 41:52:@8624.4]
  wire  output_26_25; // @[Switch.scala 41:38:@8625.4]
  wire  _T_18860; // @[Switch.scala 41:52:@8627.4]
  wire  output_26_26; // @[Switch.scala 41:38:@8628.4]
  wire  _T_18863; // @[Switch.scala 41:52:@8630.4]
  wire  output_26_27; // @[Switch.scala 41:38:@8631.4]
  wire  _T_18866; // @[Switch.scala 41:52:@8633.4]
  wire  output_26_28; // @[Switch.scala 41:38:@8634.4]
  wire  _T_18869; // @[Switch.scala 41:52:@8636.4]
  wire  output_26_29; // @[Switch.scala 41:38:@8637.4]
  wire  _T_18872; // @[Switch.scala 41:52:@8639.4]
  wire  output_26_30; // @[Switch.scala 41:38:@8640.4]
  wire  _T_18875; // @[Switch.scala 41:52:@8642.4]
  wire  output_26_31; // @[Switch.scala 41:38:@8643.4]
  wire [7:0] _T_18883; // @[Switch.scala 43:31:@8651.4]
  wire [15:0] _T_18891; // @[Switch.scala 43:31:@8659.4]
  wire [7:0] _T_18898; // @[Switch.scala 43:31:@8666.4]
  wire [31:0] _T_18907; // @[Switch.scala 43:31:@8675.4]
  wire  _T_18911; // @[Switch.scala 41:52:@8678.4]
  wire  output_27_0; // @[Switch.scala 41:38:@8679.4]
  wire  _T_18914; // @[Switch.scala 41:52:@8681.4]
  wire  output_27_1; // @[Switch.scala 41:38:@8682.4]
  wire  _T_18917; // @[Switch.scala 41:52:@8684.4]
  wire  output_27_2; // @[Switch.scala 41:38:@8685.4]
  wire  _T_18920; // @[Switch.scala 41:52:@8687.4]
  wire  output_27_3; // @[Switch.scala 41:38:@8688.4]
  wire  _T_18923; // @[Switch.scala 41:52:@8690.4]
  wire  output_27_4; // @[Switch.scala 41:38:@8691.4]
  wire  _T_18926; // @[Switch.scala 41:52:@8693.4]
  wire  output_27_5; // @[Switch.scala 41:38:@8694.4]
  wire  _T_18929; // @[Switch.scala 41:52:@8696.4]
  wire  output_27_6; // @[Switch.scala 41:38:@8697.4]
  wire  _T_18932; // @[Switch.scala 41:52:@8699.4]
  wire  output_27_7; // @[Switch.scala 41:38:@8700.4]
  wire  _T_18935; // @[Switch.scala 41:52:@8702.4]
  wire  output_27_8; // @[Switch.scala 41:38:@8703.4]
  wire  _T_18938; // @[Switch.scala 41:52:@8705.4]
  wire  output_27_9; // @[Switch.scala 41:38:@8706.4]
  wire  _T_18941; // @[Switch.scala 41:52:@8708.4]
  wire  output_27_10; // @[Switch.scala 41:38:@8709.4]
  wire  _T_18944; // @[Switch.scala 41:52:@8711.4]
  wire  output_27_11; // @[Switch.scala 41:38:@8712.4]
  wire  _T_18947; // @[Switch.scala 41:52:@8714.4]
  wire  output_27_12; // @[Switch.scala 41:38:@8715.4]
  wire  _T_18950; // @[Switch.scala 41:52:@8717.4]
  wire  output_27_13; // @[Switch.scala 41:38:@8718.4]
  wire  _T_18953; // @[Switch.scala 41:52:@8720.4]
  wire  output_27_14; // @[Switch.scala 41:38:@8721.4]
  wire  _T_18956; // @[Switch.scala 41:52:@8723.4]
  wire  output_27_15; // @[Switch.scala 41:38:@8724.4]
  wire  _T_18959; // @[Switch.scala 41:52:@8726.4]
  wire  output_27_16; // @[Switch.scala 41:38:@8727.4]
  wire  _T_18962; // @[Switch.scala 41:52:@8729.4]
  wire  output_27_17; // @[Switch.scala 41:38:@8730.4]
  wire  _T_18965; // @[Switch.scala 41:52:@8732.4]
  wire  output_27_18; // @[Switch.scala 41:38:@8733.4]
  wire  _T_18968; // @[Switch.scala 41:52:@8735.4]
  wire  output_27_19; // @[Switch.scala 41:38:@8736.4]
  wire  _T_18971; // @[Switch.scala 41:52:@8738.4]
  wire  output_27_20; // @[Switch.scala 41:38:@8739.4]
  wire  _T_18974; // @[Switch.scala 41:52:@8741.4]
  wire  output_27_21; // @[Switch.scala 41:38:@8742.4]
  wire  _T_18977; // @[Switch.scala 41:52:@8744.4]
  wire  output_27_22; // @[Switch.scala 41:38:@8745.4]
  wire  _T_18980; // @[Switch.scala 41:52:@8747.4]
  wire  output_27_23; // @[Switch.scala 41:38:@8748.4]
  wire  _T_18983; // @[Switch.scala 41:52:@8750.4]
  wire  output_27_24; // @[Switch.scala 41:38:@8751.4]
  wire  _T_18986; // @[Switch.scala 41:52:@8753.4]
  wire  output_27_25; // @[Switch.scala 41:38:@8754.4]
  wire  _T_18989; // @[Switch.scala 41:52:@8756.4]
  wire  output_27_26; // @[Switch.scala 41:38:@8757.4]
  wire  _T_18992; // @[Switch.scala 41:52:@8759.4]
  wire  output_27_27; // @[Switch.scala 41:38:@8760.4]
  wire  _T_18995; // @[Switch.scala 41:52:@8762.4]
  wire  output_27_28; // @[Switch.scala 41:38:@8763.4]
  wire  _T_18998; // @[Switch.scala 41:52:@8765.4]
  wire  output_27_29; // @[Switch.scala 41:38:@8766.4]
  wire  _T_19001; // @[Switch.scala 41:52:@8768.4]
  wire  output_27_30; // @[Switch.scala 41:38:@8769.4]
  wire  _T_19004; // @[Switch.scala 41:52:@8771.4]
  wire  output_27_31; // @[Switch.scala 41:38:@8772.4]
  wire [7:0] _T_19012; // @[Switch.scala 43:31:@8780.4]
  wire [15:0] _T_19020; // @[Switch.scala 43:31:@8788.4]
  wire [7:0] _T_19027; // @[Switch.scala 43:31:@8795.4]
  wire [31:0] _T_19036; // @[Switch.scala 43:31:@8804.4]
  wire  _T_19040; // @[Switch.scala 41:52:@8807.4]
  wire  output_28_0; // @[Switch.scala 41:38:@8808.4]
  wire  _T_19043; // @[Switch.scala 41:52:@8810.4]
  wire  output_28_1; // @[Switch.scala 41:38:@8811.4]
  wire  _T_19046; // @[Switch.scala 41:52:@8813.4]
  wire  output_28_2; // @[Switch.scala 41:38:@8814.4]
  wire  _T_19049; // @[Switch.scala 41:52:@8816.4]
  wire  output_28_3; // @[Switch.scala 41:38:@8817.4]
  wire  _T_19052; // @[Switch.scala 41:52:@8819.4]
  wire  output_28_4; // @[Switch.scala 41:38:@8820.4]
  wire  _T_19055; // @[Switch.scala 41:52:@8822.4]
  wire  output_28_5; // @[Switch.scala 41:38:@8823.4]
  wire  _T_19058; // @[Switch.scala 41:52:@8825.4]
  wire  output_28_6; // @[Switch.scala 41:38:@8826.4]
  wire  _T_19061; // @[Switch.scala 41:52:@8828.4]
  wire  output_28_7; // @[Switch.scala 41:38:@8829.4]
  wire  _T_19064; // @[Switch.scala 41:52:@8831.4]
  wire  output_28_8; // @[Switch.scala 41:38:@8832.4]
  wire  _T_19067; // @[Switch.scala 41:52:@8834.4]
  wire  output_28_9; // @[Switch.scala 41:38:@8835.4]
  wire  _T_19070; // @[Switch.scala 41:52:@8837.4]
  wire  output_28_10; // @[Switch.scala 41:38:@8838.4]
  wire  _T_19073; // @[Switch.scala 41:52:@8840.4]
  wire  output_28_11; // @[Switch.scala 41:38:@8841.4]
  wire  _T_19076; // @[Switch.scala 41:52:@8843.4]
  wire  output_28_12; // @[Switch.scala 41:38:@8844.4]
  wire  _T_19079; // @[Switch.scala 41:52:@8846.4]
  wire  output_28_13; // @[Switch.scala 41:38:@8847.4]
  wire  _T_19082; // @[Switch.scala 41:52:@8849.4]
  wire  output_28_14; // @[Switch.scala 41:38:@8850.4]
  wire  _T_19085; // @[Switch.scala 41:52:@8852.4]
  wire  output_28_15; // @[Switch.scala 41:38:@8853.4]
  wire  _T_19088; // @[Switch.scala 41:52:@8855.4]
  wire  output_28_16; // @[Switch.scala 41:38:@8856.4]
  wire  _T_19091; // @[Switch.scala 41:52:@8858.4]
  wire  output_28_17; // @[Switch.scala 41:38:@8859.4]
  wire  _T_19094; // @[Switch.scala 41:52:@8861.4]
  wire  output_28_18; // @[Switch.scala 41:38:@8862.4]
  wire  _T_19097; // @[Switch.scala 41:52:@8864.4]
  wire  output_28_19; // @[Switch.scala 41:38:@8865.4]
  wire  _T_19100; // @[Switch.scala 41:52:@8867.4]
  wire  output_28_20; // @[Switch.scala 41:38:@8868.4]
  wire  _T_19103; // @[Switch.scala 41:52:@8870.4]
  wire  output_28_21; // @[Switch.scala 41:38:@8871.4]
  wire  _T_19106; // @[Switch.scala 41:52:@8873.4]
  wire  output_28_22; // @[Switch.scala 41:38:@8874.4]
  wire  _T_19109; // @[Switch.scala 41:52:@8876.4]
  wire  output_28_23; // @[Switch.scala 41:38:@8877.4]
  wire  _T_19112; // @[Switch.scala 41:52:@8879.4]
  wire  output_28_24; // @[Switch.scala 41:38:@8880.4]
  wire  _T_19115; // @[Switch.scala 41:52:@8882.4]
  wire  output_28_25; // @[Switch.scala 41:38:@8883.4]
  wire  _T_19118; // @[Switch.scala 41:52:@8885.4]
  wire  output_28_26; // @[Switch.scala 41:38:@8886.4]
  wire  _T_19121; // @[Switch.scala 41:52:@8888.4]
  wire  output_28_27; // @[Switch.scala 41:38:@8889.4]
  wire  _T_19124; // @[Switch.scala 41:52:@8891.4]
  wire  output_28_28; // @[Switch.scala 41:38:@8892.4]
  wire  _T_19127; // @[Switch.scala 41:52:@8894.4]
  wire  output_28_29; // @[Switch.scala 41:38:@8895.4]
  wire  _T_19130; // @[Switch.scala 41:52:@8897.4]
  wire  output_28_30; // @[Switch.scala 41:38:@8898.4]
  wire  _T_19133; // @[Switch.scala 41:52:@8900.4]
  wire  output_28_31; // @[Switch.scala 41:38:@8901.4]
  wire [7:0] _T_19141; // @[Switch.scala 43:31:@8909.4]
  wire [15:0] _T_19149; // @[Switch.scala 43:31:@8917.4]
  wire [7:0] _T_19156; // @[Switch.scala 43:31:@8924.4]
  wire [31:0] _T_19165; // @[Switch.scala 43:31:@8933.4]
  wire  _T_19169; // @[Switch.scala 41:52:@8936.4]
  wire  output_29_0; // @[Switch.scala 41:38:@8937.4]
  wire  _T_19172; // @[Switch.scala 41:52:@8939.4]
  wire  output_29_1; // @[Switch.scala 41:38:@8940.4]
  wire  _T_19175; // @[Switch.scala 41:52:@8942.4]
  wire  output_29_2; // @[Switch.scala 41:38:@8943.4]
  wire  _T_19178; // @[Switch.scala 41:52:@8945.4]
  wire  output_29_3; // @[Switch.scala 41:38:@8946.4]
  wire  _T_19181; // @[Switch.scala 41:52:@8948.4]
  wire  output_29_4; // @[Switch.scala 41:38:@8949.4]
  wire  _T_19184; // @[Switch.scala 41:52:@8951.4]
  wire  output_29_5; // @[Switch.scala 41:38:@8952.4]
  wire  _T_19187; // @[Switch.scala 41:52:@8954.4]
  wire  output_29_6; // @[Switch.scala 41:38:@8955.4]
  wire  _T_19190; // @[Switch.scala 41:52:@8957.4]
  wire  output_29_7; // @[Switch.scala 41:38:@8958.4]
  wire  _T_19193; // @[Switch.scala 41:52:@8960.4]
  wire  output_29_8; // @[Switch.scala 41:38:@8961.4]
  wire  _T_19196; // @[Switch.scala 41:52:@8963.4]
  wire  output_29_9; // @[Switch.scala 41:38:@8964.4]
  wire  _T_19199; // @[Switch.scala 41:52:@8966.4]
  wire  output_29_10; // @[Switch.scala 41:38:@8967.4]
  wire  _T_19202; // @[Switch.scala 41:52:@8969.4]
  wire  output_29_11; // @[Switch.scala 41:38:@8970.4]
  wire  _T_19205; // @[Switch.scala 41:52:@8972.4]
  wire  output_29_12; // @[Switch.scala 41:38:@8973.4]
  wire  _T_19208; // @[Switch.scala 41:52:@8975.4]
  wire  output_29_13; // @[Switch.scala 41:38:@8976.4]
  wire  _T_19211; // @[Switch.scala 41:52:@8978.4]
  wire  output_29_14; // @[Switch.scala 41:38:@8979.4]
  wire  _T_19214; // @[Switch.scala 41:52:@8981.4]
  wire  output_29_15; // @[Switch.scala 41:38:@8982.4]
  wire  _T_19217; // @[Switch.scala 41:52:@8984.4]
  wire  output_29_16; // @[Switch.scala 41:38:@8985.4]
  wire  _T_19220; // @[Switch.scala 41:52:@8987.4]
  wire  output_29_17; // @[Switch.scala 41:38:@8988.4]
  wire  _T_19223; // @[Switch.scala 41:52:@8990.4]
  wire  output_29_18; // @[Switch.scala 41:38:@8991.4]
  wire  _T_19226; // @[Switch.scala 41:52:@8993.4]
  wire  output_29_19; // @[Switch.scala 41:38:@8994.4]
  wire  _T_19229; // @[Switch.scala 41:52:@8996.4]
  wire  output_29_20; // @[Switch.scala 41:38:@8997.4]
  wire  _T_19232; // @[Switch.scala 41:52:@8999.4]
  wire  output_29_21; // @[Switch.scala 41:38:@9000.4]
  wire  _T_19235; // @[Switch.scala 41:52:@9002.4]
  wire  output_29_22; // @[Switch.scala 41:38:@9003.4]
  wire  _T_19238; // @[Switch.scala 41:52:@9005.4]
  wire  output_29_23; // @[Switch.scala 41:38:@9006.4]
  wire  _T_19241; // @[Switch.scala 41:52:@9008.4]
  wire  output_29_24; // @[Switch.scala 41:38:@9009.4]
  wire  _T_19244; // @[Switch.scala 41:52:@9011.4]
  wire  output_29_25; // @[Switch.scala 41:38:@9012.4]
  wire  _T_19247; // @[Switch.scala 41:52:@9014.4]
  wire  output_29_26; // @[Switch.scala 41:38:@9015.4]
  wire  _T_19250; // @[Switch.scala 41:52:@9017.4]
  wire  output_29_27; // @[Switch.scala 41:38:@9018.4]
  wire  _T_19253; // @[Switch.scala 41:52:@9020.4]
  wire  output_29_28; // @[Switch.scala 41:38:@9021.4]
  wire  _T_19256; // @[Switch.scala 41:52:@9023.4]
  wire  output_29_29; // @[Switch.scala 41:38:@9024.4]
  wire  _T_19259; // @[Switch.scala 41:52:@9026.4]
  wire  output_29_30; // @[Switch.scala 41:38:@9027.4]
  wire  _T_19262; // @[Switch.scala 41:52:@9029.4]
  wire  output_29_31; // @[Switch.scala 41:38:@9030.4]
  wire [7:0] _T_19270; // @[Switch.scala 43:31:@9038.4]
  wire [15:0] _T_19278; // @[Switch.scala 43:31:@9046.4]
  wire [7:0] _T_19285; // @[Switch.scala 43:31:@9053.4]
  wire [31:0] _T_19294; // @[Switch.scala 43:31:@9062.4]
  wire  _T_19298; // @[Switch.scala 41:52:@9065.4]
  wire  output_30_0; // @[Switch.scala 41:38:@9066.4]
  wire  _T_19301; // @[Switch.scala 41:52:@9068.4]
  wire  output_30_1; // @[Switch.scala 41:38:@9069.4]
  wire  _T_19304; // @[Switch.scala 41:52:@9071.4]
  wire  output_30_2; // @[Switch.scala 41:38:@9072.4]
  wire  _T_19307; // @[Switch.scala 41:52:@9074.4]
  wire  output_30_3; // @[Switch.scala 41:38:@9075.4]
  wire  _T_19310; // @[Switch.scala 41:52:@9077.4]
  wire  output_30_4; // @[Switch.scala 41:38:@9078.4]
  wire  _T_19313; // @[Switch.scala 41:52:@9080.4]
  wire  output_30_5; // @[Switch.scala 41:38:@9081.4]
  wire  _T_19316; // @[Switch.scala 41:52:@9083.4]
  wire  output_30_6; // @[Switch.scala 41:38:@9084.4]
  wire  _T_19319; // @[Switch.scala 41:52:@9086.4]
  wire  output_30_7; // @[Switch.scala 41:38:@9087.4]
  wire  _T_19322; // @[Switch.scala 41:52:@9089.4]
  wire  output_30_8; // @[Switch.scala 41:38:@9090.4]
  wire  _T_19325; // @[Switch.scala 41:52:@9092.4]
  wire  output_30_9; // @[Switch.scala 41:38:@9093.4]
  wire  _T_19328; // @[Switch.scala 41:52:@9095.4]
  wire  output_30_10; // @[Switch.scala 41:38:@9096.4]
  wire  _T_19331; // @[Switch.scala 41:52:@9098.4]
  wire  output_30_11; // @[Switch.scala 41:38:@9099.4]
  wire  _T_19334; // @[Switch.scala 41:52:@9101.4]
  wire  output_30_12; // @[Switch.scala 41:38:@9102.4]
  wire  _T_19337; // @[Switch.scala 41:52:@9104.4]
  wire  output_30_13; // @[Switch.scala 41:38:@9105.4]
  wire  _T_19340; // @[Switch.scala 41:52:@9107.4]
  wire  output_30_14; // @[Switch.scala 41:38:@9108.4]
  wire  _T_19343; // @[Switch.scala 41:52:@9110.4]
  wire  output_30_15; // @[Switch.scala 41:38:@9111.4]
  wire  _T_19346; // @[Switch.scala 41:52:@9113.4]
  wire  output_30_16; // @[Switch.scala 41:38:@9114.4]
  wire  _T_19349; // @[Switch.scala 41:52:@9116.4]
  wire  output_30_17; // @[Switch.scala 41:38:@9117.4]
  wire  _T_19352; // @[Switch.scala 41:52:@9119.4]
  wire  output_30_18; // @[Switch.scala 41:38:@9120.4]
  wire  _T_19355; // @[Switch.scala 41:52:@9122.4]
  wire  output_30_19; // @[Switch.scala 41:38:@9123.4]
  wire  _T_19358; // @[Switch.scala 41:52:@9125.4]
  wire  output_30_20; // @[Switch.scala 41:38:@9126.4]
  wire  _T_19361; // @[Switch.scala 41:52:@9128.4]
  wire  output_30_21; // @[Switch.scala 41:38:@9129.4]
  wire  _T_19364; // @[Switch.scala 41:52:@9131.4]
  wire  output_30_22; // @[Switch.scala 41:38:@9132.4]
  wire  _T_19367; // @[Switch.scala 41:52:@9134.4]
  wire  output_30_23; // @[Switch.scala 41:38:@9135.4]
  wire  _T_19370; // @[Switch.scala 41:52:@9137.4]
  wire  output_30_24; // @[Switch.scala 41:38:@9138.4]
  wire  _T_19373; // @[Switch.scala 41:52:@9140.4]
  wire  output_30_25; // @[Switch.scala 41:38:@9141.4]
  wire  _T_19376; // @[Switch.scala 41:52:@9143.4]
  wire  output_30_26; // @[Switch.scala 41:38:@9144.4]
  wire  _T_19379; // @[Switch.scala 41:52:@9146.4]
  wire  output_30_27; // @[Switch.scala 41:38:@9147.4]
  wire  _T_19382; // @[Switch.scala 41:52:@9149.4]
  wire  output_30_28; // @[Switch.scala 41:38:@9150.4]
  wire  _T_19385; // @[Switch.scala 41:52:@9152.4]
  wire  output_30_29; // @[Switch.scala 41:38:@9153.4]
  wire  _T_19388; // @[Switch.scala 41:52:@9155.4]
  wire  output_30_30; // @[Switch.scala 41:38:@9156.4]
  wire  _T_19391; // @[Switch.scala 41:52:@9158.4]
  wire  output_30_31; // @[Switch.scala 41:38:@9159.4]
  wire [7:0] _T_19399; // @[Switch.scala 43:31:@9167.4]
  wire [15:0] _T_19407; // @[Switch.scala 43:31:@9175.4]
  wire [7:0] _T_19414; // @[Switch.scala 43:31:@9182.4]
  wire [31:0] _T_19423; // @[Switch.scala 43:31:@9191.4]
  wire  _T_19427; // @[Switch.scala 41:52:@9194.4]
  wire  output_31_0; // @[Switch.scala 41:38:@9195.4]
  wire  _T_19430; // @[Switch.scala 41:52:@9197.4]
  wire  output_31_1; // @[Switch.scala 41:38:@9198.4]
  wire  _T_19433; // @[Switch.scala 41:52:@9200.4]
  wire  output_31_2; // @[Switch.scala 41:38:@9201.4]
  wire  _T_19436; // @[Switch.scala 41:52:@9203.4]
  wire  output_31_3; // @[Switch.scala 41:38:@9204.4]
  wire  _T_19439; // @[Switch.scala 41:52:@9206.4]
  wire  output_31_4; // @[Switch.scala 41:38:@9207.4]
  wire  _T_19442; // @[Switch.scala 41:52:@9209.4]
  wire  output_31_5; // @[Switch.scala 41:38:@9210.4]
  wire  _T_19445; // @[Switch.scala 41:52:@9212.4]
  wire  output_31_6; // @[Switch.scala 41:38:@9213.4]
  wire  _T_19448; // @[Switch.scala 41:52:@9215.4]
  wire  output_31_7; // @[Switch.scala 41:38:@9216.4]
  wire  _T_19451; // @[Switch.scala 41:52:@9218.4]
  wire  output_31_8; // @[Switch.scala 41:38:@9219.4]
  wire  _T_19454; // @[Switch.scala 41:52:@9221.4]
  wire  output_31_9; // @[Switch.scala 41:38:@9222.4]
  wire  _T_19457; // @[Switch.scala 41:52:@9224.4]
  wire  output_31_10; // @[Switch.scala 41:38:@9225.4]
  wire  _T_19460; // @[Switch.scala 41:52:@9227.4]
  wire  output_31_11; // @[Switch.scala 41:38:@9228.4]
  wire  _T_19463; // @[Switch.scala 41:52:@9230.4]
  wire  output_31_12; // @[Switch.scala 41:38:@9231.4]
  wire  _T_19466; // @[Switch.scala 41:52:@9233.4]
  wire  output_31_13; // @[Switch.scala 41:38:@9234.4]
  wire  _T_19469; // @[Switch.scala 41:52:@9236.4]
  wire  output_31_14; // @[Switch.scala 41:38:@9237.4]
  wire  _T_19472; // @[Switch.scala 41:52:@9239.4]
  wire  output_31_15; // @[Switch.scala 41:38:@9240.4]
  wire  _T_19475; // @[Switch.scala 41:52:@9242.4]
  wire  output_31_16; // @[Switch.scala 41:38:@9243.4]
  wire  _T_19478; // @[Switch.scala 41:52:@9245.4]
  wire  output_31_17; // @[Switch.scala 41:38:@9246.4]
  wire  _T_19481; // @[Switch.scala 41:52:@9248.4]
  wire  output_31_18; // @[Switch.scala 41:38:@9249.4]
  wire  _T_19484; // @[Switch.scala 41:52:@9251.4]
  wire  output_31_19; // @[Switch.scala 41:38:@9252.4]
  wire  _T_19487; // @[Switch.scala 41:52:@9254.4]
  wire  output_31_20; // @[Switch.scala 41:38:@9255.4]
  wire  _T_19490; // @[Switch.scala 41:52:@9257.4]
  wire  output_31_21; // @[Switch.scala 41:38:@9258.4]
  wire  _T_19493; // @[Switch.scala 41:52:@9260.4]
  wire  output_31_22; // @[Switch.scala 41:38:@9261.4]
  wire  _T_19496; // @[Switch.scala 41:52:@9263.4]
  wire  output_31_23; // @[Switch.scala 41:38:@9264.4]
  wire  _T_19499; // @[Switch.scala 41:52:@9266.4]
  wire  output_31_24; // @[Switch.scala 41:38:@9267.4]
  wire  _T_19502; // @[Switch.scala 41:52:@9269.4]
  wire  output_31_25; // @[Switch.scala 41:38:@9270.4]
  wire  _T_19505; // @[Switch.scala 41:52:@9272.4]
  wire  output_31_26; // @[Switch.scala 41:38:@9273.4]
  wire  _T_19508; // @[Switch.scala 41:52:@9275.4]
  wire  output_31_27; // @[Switch.scala 41:38:@9276.4]
  wire  _T_19511; // @[Switch.scala 41:52:@9278.4]
  wire  output_31_28; // @[Switch.scala 41:38:@9279.4]
  wire  _T_19514; // @[Switch.scala 41:52:@9281.4]
  wire  output_31_29; // @[Switch.scala 41:38:@9282.4]
  wire  _T_19517; // @[Switch.scala 41:52:@9284.4]
  wire  output_31_30; // @[Switch.scala 41:38:@9285.4]
  wire  _T_19520; // @[Switch.scala 41:52:@9287.4]
  wire  output_31_31; // @[Switch.scala 41:38:@9288.4]
  wire [7:0] _T_19528; // @[Switch.scala 43:31:@9296.4]
  wire [15:0] _T_19536; // @[Switch.scala 43:31:@9304.4]
  wire [7:0] _T_19543; // @[Switch.scala 43:31:@9311.4]
  wire [31:0] _T_19552; // @[Switch.scala 43:31:@9320.4]
  assign _T_4758 = io_inAddr_0 == 5'h0; // @[Switch.scala 30:53:@10.4]
  assign valid_0_0 = io_inValid_0 & _T_4758; // @[Switch.scala 30:36:@11.4]
  assign _T_4761 = io_inAddr_1 == 5'h0; // @[Switch.scala 30:53:@13.4]
  assign valid_0_1 = io_inValid_1 & _T_4761; // @[Switch.scala 30:36:@14.4]
  assign _T_4764 = io_inAddr_2 == 5'h0; // @[Switch.scala 30:53:@16.4]
  assign valid_0_2 = io_inValid_2 & _T_4764; // @[Switch.scala 30:36:@17.4]
  assign _T_4767 = io_inAddr_3 == 5'h0; // @[Switch.scala 30:53:@19.4]
  assign valid_0_3 = io_inValid_3 & _T_4767; // @[Switch.scala 30:36:@20.4]
  assign _T_4770 = io_inAddr_4 == 5'h0; // @[Switch.scala 30:53:@22.4]
  assign valid_0_4 = io_inValid_4 & _T_4770; // @[Switch.scala 30:36:@23.4]
  assign _T_4773 = io_inAddr_5 == 5'h0; // @[Switch.scala 30:53:@25.4]
  assign valid_0_5 = io_inValid_5 & _T_4773; // @[Switch.scala 30:36:@26.4]
  assign _T_4776 = io_inAddr_6 == 5'h0; // @[Switch.scala 30:53:@28.4]
  assign valid_0_6 = io_inValid_6 & _T_4776; // @[Switch.scala 30:36:@29.4]
  assign _T_4779 = io_inAddr_7 == 5'h0; // @[Switch.scala 30:53:@31.4]
  assign valid_0_7 = io_inValid_7 & _T_4779; // @[Switch.scala 30:36:@32.4]
  assign _T_4782 = io_inAddr_8 == 5'h0; // @[Switch.scala 30:53:@34.4]
  assign valid_0_8 = io_inValid_8 & _T_4782; // @[Switch.scala 30:36:@35.4]
  assign _T_4785 = io_inAddr_9 == 5'h0; // @[Switch.scala 30:53:@37.4]
  assign valid_0_9 = io_inValid_9 & _T_4785; // @[Switch.scala 30:36:@38.4]
  assign _T_4788 = io_inAddr_10 == 5'h0; // @[Switch.scala 30:53:@40.4]
  assign valid_0_10 = io_inValid_10 & _T_4788; // @[Switch.scala 30:36:@41.4]
  assign _T_4791 = io_inAddr_11 == 5'h0; // @[Switch.scala 30:53:@43.4]
  assign valid_0_11 = io_inValid_11 & _T_4791; // @[Switch.scala 30:36:@44.4]
  assign _T_4794 = io_inAddr_12 == 5'h0; // @[Switch.scala 30:53:@46.4]
  assign valid_0_12 = io_inValid_12 & _T_4794; // @[Switch.scala 30:36:@47.4]
  assign _T_4797 = io_inAddr_13 == 5'h0; // @[Switch.scala 30:53:@49.4]
  assign valid_0_13 = io_inValid_13 & _T_4797; // @[Switch.scala 30:36:@50.4]
  assign _T_4800 = io_inAddr_14 == 5'h0; // @[Switch.scala 30:53:@52.4]
  assign valid_0_14 = io_inValid_14 & _T_4800; // @[Switch.scala 30:36:@53.4]
  assign _T_4803 = io_inAddr_15 == 5'h0; // @[Switch.scala 30:53:@55.4]
  assign valid_0_15 = io_inValid_15 & _T_4803; // @[Switch.scala 30:36:@56.4]
  assign _T_4806 = io_inAddr_16 == 5'h0; // @[Switch.scala 30:53:@58.4]
  assign valid_0_16 = io_inValid_16 & _T_4806; // @[Switch.scala 30:36:@59.4]
  assign _T_4809 = io_inAddr_17 == 5'h0; // @[Switch.scala 30:53:@61.4]
  assign valid_0_17 = io_inValid_17 & _T_4809; // @[Switch.scala 30:36:@62.4]
  assign _T_4812 = io_inAddr_18 == 5'h0; // @[Switch.scala 30:53:@64.4]
  assign valid_0_18 = io_inValid_18 & _T_4812; // @[Switch.scala 30:36:@65.4]
  assign _T_4815 = io_inAddr_19 == 5'h0; // @[Switch.scala 30:53:@67.4]
  assign valid_0_19 = io_inValid_19 & _T_4815; // @[Switch.scala 30:36:@68.4]
  assign _T_4818 = io_inAddr_20 == 5'h0; // @[Switch.scala 30:53:@70.4]
  assign valid_0_20 = io_inValid_20 & _T_4818; // @[Switch.scala 30:36:@71.4]
  assign _T_4821 = io_inAddr_21 == 5'h0; // @[Switch.scala 30:53:@73.4]
  assign valid_0_21 = io_inValid_21 & _T_4821; // @[Switch.scala 30:36:@74.4]
  assign _T_4824 = io_inAddr_22 == 5'h0; // @[Switch.scala 30:53:@76.4]
  assign valid_0_22 = io_inValid_22 & _T_4824; // @[Switch.scala 30:36:@77.4]
  assign _T_4827 = io_inAddr_23 == 5'h0; // @[Switch.scala 30:53:@79.4]
  assign valid_0_23 = io_inValid_23 & _T_4827; // @[Switch.scala 30:36:@80.4]
  assign _T_4830 = io_inAddr_24 == 5'h0; // @[Switch.scala 30:53:@82.4]
  assign valid_0_24 = io_inValid_24 & _T_4830; // @[Switch.scala 30:36:@83.4]
  assign _T_4833 = io_inAddr_25 == 5'h0; // @[Switch.scala 30:53:@85.4]
  assign valid_0_25 = io_inValid_25 & _T_4833; // @[Switch.scala 30:36:@86.4]
  assign _T_4836 = io_inAddr_26 == 5'h0; // @[Switch.scala 30:53:@88.4]
  assign valid_0_26 = io_inValid_26 & _T_4836; // @[Switch.scala 30:36:@89.4]
  assign _T_4839 = io_inAddr_27 == 5'h0; // @[Switch.scala 30:53:@91.4]
  assign valid_0_27 = io_inValid_27 & _T_4839; // @[Switch.scala 30:36:@92.4]
  assign _T_4842 = io_inAddr_28 == 5'h0; // @[Switch.scala 30:53:@94.4]
  assign valid_0_28 = io_inValid_28 & _T_4842; // @[Switch.scala 30:36:@95.4]
  assign _T_4845 = io_inAddr_29 == 5'h0; // @[Switch.scala 30:53:@97.4]
  assign valid_0_29 = io_inValid_29 & _T_4845; // @[Switch.scala 30:36:@98.4]
  assign _T_4848 = io_inAddr_30 == 5'h0; // @[Switch.scala 30:53:@100.4]
  assign valid_0_30 = io_inValid_30 & _T_4848; // @[Switch.scala 30:36:@101.4]
  assign _T_4851 = io_inAddr_31 == 5'h0; // @[Switch.scala 30:53:@103.4]
  assign valid_0_31 = io_inValid_31 & _T_4851; // @[Switch.scala 30:36:@104.4]
  assign _T_4885 = valid_0_30 ? 5'h1e : 5'h1f; // @[Mux.scala 31:69:@106.4]
  assign _T_4886 = valid_0_29 ? 5'h1d : _T_4885; // @[Mux.scala 31:69:@107.4]
  assign _T_4887 = valid_0_28 ? 5'h1c : _T_4886; // @[Mux.scala 31:69:@108.4]
  assign _T_4888 = valid_0_27 ? 5'h1b : _T_4887; // @[Mux.scala 31:69:@109.4]
  assign _T_4889 = valid_0_26 ? 5'h1a : _T_4888; // @[Mux.scala 31:69:@110.4]
  assign _T_4890 = valid_0_25 ? 5'h19 : _T_4889; // @[Mux.scala 31:69:@111.4]
  assign _T_4891 = valid_0_24 ? 5'h18 : _T_4890; // @[Mux.scala 31:69:@112.4]
  assign _T_4892 = valid_0_23 ? 5'h17 : _T_4891; // @[Mux.scala 31:69:@113.4]
  assign _T_4893 = valid_0_22 ? 5'h16 : _T_4892; // @[Mux.scala 31:69:@114.4]
  assign _T_4894 = valid_0_21 ? 5'h15 : _T_4893; // @[Mux.scala 31:69:@115.4]
  assign _T_4895 = valid_0_20 ? 5'h14 : _T_4894; // @[Mux.scala 31:69:@116.4]
  assign _T_4896 = valid_0_19 ? 5'h13 : _T_4895; // @[Mux.scala 31:69:@117.4]
  assign _T_4897 = valid_0_18 ? 5'h12 : _T_4896; // @[Mux.scala 31:69:@118.4]
  assign _T_4898 = valid_0_17 ? 5'h11 : _T_4897; // @[Mux.scala 31:69:@119.4]
  assign _T_4899 = valid_0_16 ? 5'h10 : _T_4898; // @[Mux.scala 31:69:@120.4]
  assign _T_4900 = valid_0_15 ? 5'hf : _T_4899; // @[Mux.scala 31:69:@121.4]
  assign _T_4901 = valid_0_14 ? 5'he : _T_4900; // @[Mux.scala 31:69:@122.4]
  assign _T_4902 = valid_0_13 ? 5'hd : _T_4901; // @[Mux.scala 31:69:@123.4]
  assign _T_4903 = valid_0_12 ? 5'hc : _T_4902; // @[Mux.scala 31:69:@124.4]
  assign _T_4904 = valid_0_11 ? 5'hb : _T_4903; // @[Mux.scala 31:69:@125.4]
  assign _T_4905 = valid_0_10 ? 5'ha : _T_4904; // @[Mux.scala 31:69:@126.4]
  assign _T_4906 = valid_0_9 ? 5'h9 : _T_4905; // @[Mux.scala 31:69:@127.4]
  assign _T_4907 = valid_0_8 ? 5'h8 : _T_4906; // @[Mux.scala 31:69:@128.4]
  assign _T_4908 = valid_0_7 ? 5'h7 : _T_4907; // @[Mux.scala 31:69:@129.4]
  assign _T_4909 = valid_0_6 ? 5'h6 : _T_4908; // @[Mux.scala 31:69:@130.4]
  assign _T_4910 = valid_0_5 ? 5'h5 : _T_4909; // @[Mux.scala 31:69:@131.4]
  assign _T_4911 = valid_0_4 ? 5'h4 : _T_4910; // @[Mux.scala 31:69:@132.4]
  assign _T_4912 = valid_0_3 ? 5'h3 : _T_4911; // @[Mux.scala 31:69:@133.4]
  assign _T_4913 = valid_0_2 ? 5'h2 : _T_4912; // @[Mux.scala 31:69:@134.4]
  assign _T_4914 = valid_0_1 ? 5'h1 : _T_4913; // @[Mux.scala 31:69:@135.4]
  assign select_0 = valid_0_0 ? 5'h0 : _T_4914; // @[Mux.scala 31:69:@136.4]
  assign _GEN_1 = 5'h1 == select_0 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@138.4]
  assign _GEN_2 = 5'h2 == select_0 ? io_inData_2 : _GEN_1; // @[Switch.scala 33:19:@138.4]
  assign _GEN_3 = 5'h3 == select_0 ? io_inData_3 : _GEN_2; // @[Switch.scala 33:19:@138.4]
  assign _GEN_4 = 5'h4 == select_0 ? io_inData_4 : _GEN_3; // @[Switch.scala 33:19:@138.4]
  assign _GEN_5 = 5'h5 == select_0 ? io_inData_5 : _GEN_4; // @[Switch.scala 33:19:@138.4]
  assign _GEN_6 = 5'h6 == select_0 ? io_inData_6 : _GEN_5; // @[Switch.scala 33:19:@138.4]
  assign _GEN_7 = 5'h7 == select_0 ? io_inData_7 : _GEN_6; // @[Switch.scala 33:19:@138.4]
  assign _GEN_8 = 5'h8 == select_0 ? io_inData_8 : _GEN_7; // @[Switch.scala 33:19:@138.4]
  assign _GEN_9 = 5'h9 == select_0 ? io_inData_9 : _GEN_8; // @[Switch.scala 33:19:@138.4]
  assign _GEN_10 = 5'ha == select_0 ? io_inData_10 : _GEN_9; // @[Switch.scala 33:19:@138.4]
  assign _GEN_11 = 5'hb == select_0 ? io_inData_11 : _GEN_10; // @[Switch.scala 33:19:@138.4]
  assign _GEN_12 = 5'hc == select_0 ? io_inData_12 : _GEN_11; // @[Switch.scala 33:19:@138.4]
  assign _GEN_13 = 5'hd == select_0 ? io_inData_13 : _GEN_12; // @[Switch.scala 33:19:@138.4]
  assign _GEN_14 = 5'he == select_0 ? io_inData_14 : _GEN_13; // @[Switch.scala 33:19:@138.4]
  assign _GEN_15 = 5'hf == select_0 ? io_inData_15 : _GEN_14; // @[Switch.scala 33:19:@138.4]
  assign _GEN_16 = 5'h10 == select_0 ? io_inData_16 : _GEN_15; // @[Switch.scala 33:19:@138.4]
  assign _GEN_17 = 5'h11 == select_0 ? io_inData_17 : _GEN_16; // @[Switch.scala 33:19:@138.4]
  assign _GEN_18 = 5'h12 == select_0 ? io_inData_18 : _GEN_17; // @[Switch.scala 33:19:@138.4]
  assign _GEN_19 = 5'h13 == select_0 ? io_inData_19 : _GEN_18; // @[Switch.scala 33:19:@138.4]
  assign _GEN_20 = 5'h14 == select_0 ? io_inData_20 : _GEN_19; // @[Switch.scala 33:19:@138.4]
  assign _GEN_21 = 5'h15 == select_0 ? io_inData_21 : _GEN_20; // @[Switch.scala 33:19:@138.4]
  assign _GEN_22 = 5'h16 == select_0 ? io_inData_22 : _GEN_21; // @[Switch.scala 33:19:@138.4]
  assign _GEN_23 = 5'h17 == select_0 ? io_inData_23 : _GEN_22; // @[Switch.scala 33:19:@138.4]
  assign _GEN_24 = 5'h18 == select_0 ? io_inData_24 : _GEN_23; // @[Switch.scala 33:19:@138.4]
  assign _GEN_25 = 5'h19 == select_0 ? io_inData_25 : _GEN_24; // @[Switch.scala 33:19:@138.4]
  assign _GEN_26 = 5'h1a == select_0 ? io_inData_26 : _GEN_25; // @[Switch.scala 33:19:@138.4]
  assign _GEN_27 = 5'h1b == select_0 ? io_inData_27 : _GEN_26; // @[Switch.scala 33:19:@138.4]
  assign _GEN_28 = 5'h1c == select_0 ? io_inData_28 : _GEN_27; // @[Switch.scala 33:19:@138.4]
  assign _GEN_29 = 5'h1d == select_0 ? io_inData_29 : _GEN_28; // @[Switch.scala 33:19:@138.4]
  assign _GEN_30 = 5'h1e == select_0 ? io_inData_30 : _GEN_29; // @[Switch.scala 33:19:@138.4]
  assign _T_4923 = {valid_0_7,valid_0_6,valid_0_5,valid_0_4,valid_0_3,valid_0_2,valid_0_1,valid_0_0}; // @[Switch.scala 34:32:@145.4]
  assign _T_4931 = {valid_0_15,valid_0_14,valid_0_13,valid_0_12,valid_0_11,valid_0_10,valid_0_9,valid_0_8,_T_4923}; // @[Switch.scala 34:32:@153.4]
  assign _T_4938 = {valid_0_23,valid_0_22,valid_0_21,valid_0_20,valid_0_19,valid_0_18,valid_0_17,valid_0_16}; // @[Switch.scala 34:32:@160.4]
  assign _T_4947 = {valid_0_31,valid_0_30,valid_0_29,valid_0_28,valid_0_27,valid_0_26,valid_0_25,valid_0_24,_T_4938,_T_4931}; // @[Switch.scala 34:32:@169.4]
  assign _T_4951 = io_inAddr_0 == 5'h1; // @[Switch.scala 30:53:@172.4]
  assign valid_1_0 = io_inValid_0 & _T_4951; // @[Switch.scala 30:36:@173.4]
  assign _T_4954 = io_inAddr_1 == 5'h1; // @[Switch.scala 30:53:@175.4]
  assign valid_1_1 = io_inValid_1 & _T_4954; // @[Switch.scala 30:36:@176.4]
  assign _T_4957 = io_inAddr_2 == 5'h1; // @[Switch.scala 30:53:@178.4]
  assign valid_1_2 = io_inValid_2 & _T_4957; // @[Switch.scala 30:36:@179.4]
  assign _T_4960 = io_inAddr_3 == 5'h1; // @[Switch.scala 30:53:@181.4]
  assign valid_1_3 = io_inValid_3 & _T_4960; // @[Switch.scala 30:36:@182.4]
  assign _T_4963 = io_inAddr_4 == 5'h1; // @[Switch.scala 30:53:@184.4]
  assign valid_1_4 = io_inValid_4 & _T_4963; // @[Switch.scala 30:36:@185.4]
  assign _T_4966 = io_inAddr_5 == 5'h1; // @[Switch.scala 30:53:@187.4]
  assign valid_1_5 = io_inValid_5 & _T_4966; // @[Switch.scala 30:36:@188.4]
  assign _T_4969 = io_inAddr_6 == 5'h1; // @[Switch.scala 30:53:@190.4]
  assign valid_1_6 = io_inValid_6 & _T_4969; // @[Switch.scala 30:36:@191.4]
  assign _T_4972 = io_inAddr_7 == 5'h1; // @[Switch.scala 30:53:@193.4]
  assign valid_1_7 = io_inValid_7 & _T_4972; // @[Switch.scala 30:36:@194.4]
  assign _T_4975 = io_inAddr_8 == 5'h1; // @[Switch.scala 30:53:@196.4]
  assign valid_1_8 = io_inValid_8 & _T_4975; // @[Switch.scala 30:36:@197.4]
  assign _T_4978 = io_inAddr_9 == 5'h1; // @[Switch.scala 30:53:@199.4]
  assign valid_1_9 = io_inValid_9 & _T_4978; // @[Switch.scala 30:36:@200.4]
  assign _T_4981 = io_inAddr_10 == 5'h1; // @[Switch.scala 30:53:@202.4]
  assign valid_1_10 = io_inValid_10 & _T_4981; // @[Switch.scala 30:36:@203.4]
  assign _T_4984 = io_inAddr_11 == 5'h1; // @[Switch.scala 30:53:@205.4]
  assign valid_1_11 = io_inValid_11 & _T_4984; // @[Switch.scala 30:36:@206.4]
  assign _T_4987 = io_inAddr_12 == 5'h1; // @[Switch.scala 30:53:@208.4]
  assign valid_1_12 = io_inValid_12 & _T_4987; // @[Switch.scala 30:36:@209.4]
  assign _T_4990 = io_inAddr_13 == 5'h1; // @[Switch.scala 30:53:@211.4]
  assign valid_1_13 = io_inValid_13 & _T_4990; // @[Switch.scala 30:36:@212.4]
  assign _T_4993 = io_inAddr_14 == 5'h1; // @[Switch.scala 30:53:@214.4]
  assign valid_1_14 = io_inValid_14 & _T_4993; // @[Switch.scala 30:36:@215.4]
  assign _T_4996 = io_inAddr_15 == 5'h1; // @[Switch.scala 30:53:@217.4]
  assign valid_1_15 = io_inValid_15 & _T_4996; // @[Switch.scala 30:36:@218.4]
  assign _T_4999 = io_inAddr_16 == 5'h1; // @[Switch.scala 30:53:@220.4]
  assign valid_1_16 = io_inValid_16 & _T_4999; // @[Switch.scala 30:36:@221.4]
  assign _T_5002 = io_inAddr_17 == 5'h1; // @[Switch.scala 30:53:@223.4]
  assign valid_1_17 = io_inValid_17 & _T_5002; // @[Switch.scala 30:36:@224.4]
  assign _T_5005 = io_inAddr_18 == 5'h1; // @[Switch.scala 30:53:@226.4]
  assign valid_1_18 = io_inValid_18 & _T_5005; // @[Switch.scala 30:36:@227.4]
  assign _T_5008 = io_inAddr_19 == 5'h1; // @[Switch.scala 30:53:@229.4]
  assign valid_1_19 = io_inValid_19 & _T_5008; // @[Switch.scala 30:36:@230.4]
  assign _T_5011 = io_inAddr_20 == 5'h1; // @[Switch.scala 30:53:@232.4]
  assign valid_1_20 = io_inValid_20 & _T_5011; // @[Switch.scala 30:36:@233.4]
  assign _T_5014 = io_inAddr_21 == 5'h1; // @[Switch.scala 30:53:@235.4]
  assign valid_1_21 = io_inValid_21 & _T_5014; // @[Switch.scala 30:36:@236.4]
  assign _T_5017 = io_inAddr_22 == 5'h1; // @[Switch.scala 30:53:@238.4]
  assign valid_1_22 = io_inValid_22 & _T_5017; // @[Switch.scala 30:36:@239.4]
  assign _T_5020 = io_inAddr_23 == 5'h1; // @[Switch.scala 30:53:@241.4]
  assign valid_1_23 = io_inValid_23 & _T_5020; // @[Switch.scala 30:36:@242.4]
  assign _T_5023 = io_inAddr_24 == 5'h1; // @[Switch.scala 30:53:@244.4]
  assign valid_1_24 = io_inValid_24 & _T_5023; // @[Switch.scala 30:36:@245.4]
  assign _T_5026 = io_inAddr_25 == 5'h1; // @[Switch.scala 30:53:@247.4]
  assign valid_1_25 = io_inValid_25 & _T_5026; // @[Switch.scala 30:36:@248.4]
  assign _T_5029 = io_inAddr_26 == 5'h1; // @[Switch.scala 30:53:@250.4]
  assign valid_1_26 = io_inValid_26 & _T_5029; // @[Switch.scala 30:36:@251.4]
  assign _T_5032 = io_inAddr_27 == 5'h1; // @[Switch.scala 30:53:@253.4]
  assign valid_1_27 = io_inValid_27 & _T_5032; // @[Switch.scala 30:36:@254.4]
  assign _T_5035 = io_inAddr_28 == 5'h1; // @[Switch.scala 30:53:@256.4]
  assign valid_1_28 = io_inValid_28 & _T_5035; // @[Switch.scala 30:36:@257.4]
  assign _T_5038 = io_inAddr_29 == 5'h1; // @[Switch.scala 30:53:@259.4]
  assign valid_1_29 = io_inValid_29 & _T_5038; // @[Switch.scala 30:36:@260.4]
  assign _T_5041 = io_inAddr_30 == 5'h1; // @[Switch.scala 30:53:@262.4]
  assign valid_1_30 = io_inValid_30 & _T_5041; // @[Switch.scala 30:36:@263.4]
  assign _T_5044 = io_inAddr_31 == 5'h1; // @[Switch.scala 30:53:@265.4]
  assign valid_1_31 = io_inValid_31 & _T_5044; // @[Switch.scala 30:36:@266.4]
  assign _T_5078 = valid_1_30 ? 5'h1e : 5'h1f; // @[Mux.scala 31:69:@268.4]
  assign _T_5079 = valid_1_29 ? 5'h1d : _T_5078; // @[Mux.scala 31:69:@269.4]
  assign _T_5080 = valid_1_28 ? 5'h1c : _T_5079; // @[Mux.scala 31:69:@270.4]
  assign _T_5081 = valid_1_27 ? 5'h1b : _T_5080; // @[Mux.scala 31:69:@271.4]
  assign _T_5082 = valid_1_26 ? 5'h1a : _T_5081; // @[Mux.scala 31:69:@272.4]
  assign _T_5083 = valid_1_25 ? 5'h19 : _T_5082; // @[Mux.scala 31:69:@273.4]
  assign _T_5084 = valid_1_24 ? 5'h18 : _T_5083; // @[Mux.scala 31:69:@274.4]
  assign _T_5085 = valid_1_23 ? 5'h17 : _T_5084; // @[Mux.scala 31:69:@275.4]
  assign _T_5086 = valid_1_22 ? 5'h16 : _T_5085; // @[Mux.scala 31:69:@276.4]
  assign _T_5087 = valid_1_21 ? 5'h15 : _T_5086; // @[Mux.scala 31:69:@277.4]
  assign _T_5088 = valid_1_20 ? 5'h14 : _T_5087; // @[Mux.scala 31:69:@278.4]
  assign _T_5089 = valid_1_19 ? 5'h13 : _T_5088; // @[Mux.scala 31:69:@279.4]
  assign _T_5090 = valid_1_18 ? 5'h12 : _T_5089; // @[Mux.scala 31:69:@280.4]
  assign _T_5091 = valid_1_17 ? 5'h11 : _T_5090; // @[Mux.scala 31:69:@281.4]
  assign _T_5092 = valid_1_16 ? 5'h10 : _T_5091; // @[Mux.scala 31:69:@282.4]
  assign _T_5093 = valid_1_15 ? 5'hf : _T_5092; // @[Mux.scala 31:69:@283.4]
  assign _T_5094 = valid_1_14 ? 5'he : _T_5093; // @[Mux.scala 31:69:@284.4]
  assign _T_5095 = valid_1_13 ? 5'hd : _T_5094; // @[Mux.scala 31:69:@285.4]
  assign _T_5096 = valid_1_12 ? 5'hc : _T_5095; // @[Mux.scala 31:69:@286.4]
  assign _T_5097 = valid_1_11 ? 5'hb : _T_5096; // @[Mux.scala 31:69:@287.4]
  assign _T_5098 = valid_1_10 ? 5'ha : _T_5097; // @[Mux.scala 31:69:@288.4]
  assign _T_5099 = valid_1_9 ? 5'h9 : _T_5098; // @[Mux.scala 31:69:@289.4]
  assign _T_5100 = valid_1_8 ? 5'h8 : _T_5099; // @[Mux.scala 31:69:@290.4]
  assign _T_5101 = valid_1_7 ? 5'h7 : _T_5100; // @[Mux.scala 31:69:@291.4]
  assign _T_5102 = valid_1_6 ? 5'h6 : _T_5101; // @[Mux.scala 31:69:@292.4]
  assign _T_5103 = valid_1_5 ? 5'h5 : _T_5102; // @[Mux.scala 31:69:@293.4]
  assign _T_5104 = valid_1_4 ? 5'h4 : _T_5103; // @[Mux.scala 31:69:@294.4]
  assign _T_5105 = valid_1_3 ? 5'h3 : _T_5104; // @[Mux.scala 31:69:@295.4]
  assign _T_5106 = valid_1_2 ? 5'h2 : _T_5105; // @[Mux.scala 31:69:@296.4]
  assign _T_5107 = valid_1_1 ? 5'h1 : _T_5106; // @[Mux.scala 31:69:@297.4]
  assign select_1 = valid_1_0 ? 5'h0 : _T_5107; // @[Mux.scala 31:69:@298.4]
  assign _GEN_33 = 5'h1 == select_1 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@300.4]
  assign _GEN_34 = 5'h2 == select_1 ? io_inData_2 : _GEN_33; // @[Switch.scala 33:19:@300.4]
  assign _GEN_35 = 5'h3 == select_1 ? io_inData_3 : _GEN_34; // @[Switch.scala 33:19:@300.4]
  assign _GEN_36 = 5'h4 == select_1 ? io_inData_4 : _GEN_35; // @[Switch.scala 33:19:@300.4]
  assign _GEN_37 = 5'h5 == select_1 ? io_inData_5 : _GEN_36; // @[Switch.scala 33:19:@300.4]
  assign _GEN_38 = 5'h6 == select_1 ? io_inData_6 : _GEN_37; // @[Switch.scala 33:19:@300.4]
  assign _GEN_39 = 5'h7 == select_1 ? io_inData_7 : _GEN_38; // @[Switch.scala 33:19:@300.4]
  assign _GEN_40 = 5'h8 == select_1 ? io_inData_8 : _GEN_39; // @[Switch.scala 33:19:@300.4]
  assign _GEN_41 = 5'h9 == select_1 ? io_inData_9 : _GEN_40; // @[Switch.scala 33:19:@300.4]
  assign _GEN_42 = 5'ha == select_1 ? io_inData_10 : _GEN_41; // @[Switch.scala 33:19:@300.4]
  assign _GEN_43 = 5'hb == select_1 ? io_inData_11 : _GEN_42; // @[Switch.scala 33:19:@300.4]
  assign _GEN_44 = 5'hc == select_1 ? io_inData_12 : _GEN_43; // @[Switch.scala 33:19:@300.4]
  assign _GEN_45 = 5'hd == select_1 ? io_inData_13 : _GEN_44; // @[Switch.scala 33:19:@300.4]
  assign _GEN_46 = 5'he == select_1 ? io_inData_14 : _GEN_45; // @[Switch.scala 33:19:@300.4]
  assign _GEN_47 = 5'hf == select_1 ? io_inData_15 : _GEN_46; // @[Switch.scala 33:19:@300.4]
  assign _GEN_48 = 5'h10 == select_1 ? io_inData_16 : _GEN_47; // @[Switch.scala 33:19:@300.4]
  assign _GEN_49 = 5'h11 == select_1 ? io_inData_17 : _GEN_48; // @[Switch.scala 33:19:@300.4]
  assign _GEN_50 = 5'h12 == select_1 ? io_inData_18 : _GEN_49; // @[Switch.scala 33:19:@300.4]
  assign _GEN_51 = 5'h13 == select_1 ? io_inData_19 : _GEN_50; // @[Switch.scala 33:19:@300.4]
  assign _GEN_52 = 5'h14 == select_1 ? io_inData_20 : _GEN_51; // @[Switch.scala 33:19:@300.4]
  assign _GEN_53 = 5'h15 == select_1 ? io_inData_21 : _GEN_52; // @[Switch.scala 33:19:@300.4]
  assign _GEN_54 = 5'h16 == select_1 ? io_inData_22 : _GEN_53; // @[Switch.scala 33:19:@300.4]
  assign _GEN_55 = 5'h17 == select_1 ? io_inData_23 : _GEN_54; // @[Switch.scala 33:19:@300.4]
  assign _GEN_56 = 5'h18 == select_1 ? io_inData_24 : _GEN_55; // @[Switch.scala 33:19:@300.4]
  assign _GEN_57 = 5'h19 == select_1 ? io_inData_25 : _GEN_56; // @[Switch.scala 33:19:@300.4]
  assign _GEN_58 = 5'h1a == select_1 ? io_inData_26 : _GEN_57; // @[Switch.scala 33:19:@300.4]
  assign _GEN_59 = 5'h1b == select_1 ? io_inData_27 : _GEN_58; // @[Switch.scala 33:19:@300.4]
  assign _GEN_60 = 5'h1c == select_1 ? io_inData_28 : _GEN_59; // @[Switch.scala 33:19:@300.4]
  assign _GEN_61 = 5'h1d == select_1 ? io_inData_29 : _GEN_60; // @[Switch.scala 33:19:@300.4]
  assign _GEN_62 = 5'h1e == select_1 ? io_inData_30 : _GEN_61; // @[Switch.scala 33:19:@300.4]
  assign _T_5116 = {valid_1_7,valid_1_6,valid_1_5,valid_1_4,valid_1_3,valid_1_2,valid_1_1,valid_1_0}; // @[Switch.scala 34:32:@307.4]
  assign _T_5124 = {valid_1_15,valid_1_14,valid_1_13,valid_1_12,valid_1_11,valid_1_10,valid_1_9,valid_1_8,_T_5116}; // @[Switch.scala 34:32:@315.4]
  assign _T_5131 = {valid_1_23,valid_1_22,valid_1_21,valid_1_20,valid_1_19,valid_1_18,valid_1_17,valid_1_16}; // @[Switch.scala 34:32:@322.4]
  assign _T_5140 = {valid_1_31,valid_1_30,valid_1_29,valid_1_28,valid_1_27,valid_1_26,valid_1_25,valid_1_24,_T_5131,_T_5124}; // @[Switch.scala 34:32:@331.4]
  assign _T_5144 = io_inAddr_0 == 5'h2; // @[Switch.scala 30:53:@334.4]
  assign valid_2_0 = io_inValid_0 & _T_5144; // @[Switch.scala 30:36:@335.4]
  assign _T_5147 = io_inAddr_1 == 5'h2; // @[Switch.scala 30:53:@337.4]
  assign valid_2_1 = io_inValid_1 & _T_5147; // @[Switch.scala 30:36:@338.4]
  assign _T_5150 = io_inAddr_2 == 5'h2; // @[Switch.scala 30:53:@340.4]
  assign valid_2_2 = io_inValid_2 & _T_5150; // @[Switch.scala 30:36:@341.4]
  assign _T_5153 = io_inAddr_3 == 5'h2; // @[Switch.scala 30:53:@343.4]
  assign valid_2_3 = io_inValid_3 & _T_5153; // @[Switch.scala 30:36:@344.4]
  assign _T_5156 = io_inAddr_4 == 5'h2; // @[Switch.scala 30:53:@346.4]
  assign valid_2_4 = io_inValid_4 & _T_5156; // @[Switch.scala 30:36:@347.4]
  assign _T_5159 = io_inAddr_5 == 5'h2; // @[Switch.scala 30:53:@349.4]
  assign valid_2_5 = io_inValid_5 & _T_5159; // @[Switch.scala 30:36:@350.4]
  assign _T_5162 = io_inAddr_6 == 5'h2; // @[Switch.scala 30:53:@352.4]
  assign valid_2_6 = io_inValid_6 & _T_5162; // @[Switch.scala 30:36:@353.4]
  assign _T_5165 = io_inAddr_7 == 5'h2; // @[Switch.scala 30:53:@355.4]
  assign valid_2_7 = io_inValid_7 & _T_5165; // @[Switch.scala 30:36:@356.4]
  assign _T_5168 = io_inAddr_8 == 5'h2; // @[Switch.scala 30:53:@358.4]
  assign valid_2_8 = io_inValid_8 & _T_5168; // @[Switch.scala 30:36:@359.4]
  assign _T_5171 = io_inAddr_9 == 5'h2; // @[Switch.scala 30:53:@361.4]
  assign valid_2_9 = io_inValid_9 & _T_5171; // @[Switch.scala 30:36:@362.4]
  assign _T_5174 = io_inAddr_10 == 5'h2; // @[Switch.scala 30:53:@364.4]
  assign valid_2_10 = io_inValid_10 & _T_5174; // @[Switch.scala 30:36:@365.4]
  assign _T_5177 = io_inAddr_11 == 5'h2; // @[Switch.scala 30:53:@367.4]
  assign valid_2_11 = io_inValid_11 & _T_5177; // @[Switch.scala 30:36:@368.4]
  assign _T_5180 = io_inAddr_12 == 5'h2; // @[Switch.scala 30:53:@370.4]
  assign valid_2_12 = io_inValid_12 & _T_5180; // @[Switch.scala 30:36:@371.4]
  assign _T_5183 = io_inAddr_13 == 5'h2; // @[Switch.scala 30:53:@373.4]
  assign valid_2_13 = io_inValid_13 & _T_5183; // @[Switch.scala 30:36:@374.4]
  assign _T_5186 = io_inAddr_14 == 5'h2; // @[Switch.scala 30:53:@376.4]
  assign valid_2_14 = io_inValid_14 & _T_5186; // @[Switch.scala 30:36:@377.4]
  assign _T_5189 = io_inAddr_15 == 5'h2; // @[Switch.scala 30:53:@379.4]
  assign valid_2_15 = io_inValid_15 & _T_5189; // @[Switch.scala 30:36:@380.4]
  assign _T_5192 = io_inAddr_16 == 5'h2; // @[Switch.scala 30:53:@382.4]
  assign valid_2_16 = io_inValid_16 & _T_5192; // @[Switch.scala 30:36:@383.4]
  assign _T_5195 = io_inAddr_17 == 5'h2; // @[Switch.scala 30:53:@385.4]
  assign valid_2_17 = io_inValid_17 & _T_5195; // @[Switch.scala 30:36:@386.4]
  assign _T_5198 = io_inAddr_18 == 5'h2; // @[Switch.scala 30:53:@388.4]
  assign valid_2_18 = io_inValid_18 & _T_5198; // @[Switch.scala 30:36:@389.4]
  assign _T_5201 = io_inAddr_19 == 5'h2; // @[Switch.scala 30:53:@391.4]
  assign valid_2_19 = io_inValid_19 & _T_5201; // @[Switch.scala 30:36:@392.4]
  assign _T_5204 = io_inAddr_20 == 5'h2; // @[Switch.scala 30:53:@394.4]
  assign valid_2_20 = io_inValid_20 & _T_5204; // @[Switch.scala 30:36:@395.4]
  assign _T_5207 = io_inAddr_21 == 5'h2; // @[Switch.scala 30:53:@397.4]
  assign valid_2_21 = io_inValid_21 & _T_5207; // @[Switch.scala 30:36:@398.4]
  assign _T_5210 = io_inAddr_22 == 5'h2; // @[Switch.scala 30:53:@400.4]
  assign valid_2_22 = io_inValid_22 & _T_5210; // @[Switch.scala 30:36:@401.4]
  assign _T_5213 = io_inAddr_23 == 5'h2; // @[Switch.scala 30:53:@403.4]
  assign valid_2_23 = io_inValid_23 & _T_5213; // @[Switch.scala 30:36:@404.4]
  assign _T_5216 = io_inAddr_24 == 5'h2; // @[Switch.scala 30:53:@406.4]
  assign valid_2_24 = io_inValid_24 & _T_5216; // @[Switch.scala 30:36:@407.4]
  assign _T_5219 = io_inAddr_25 == 5'h2; // @[Switch.scala 30:53:@409.4]
  assign valid_2_25 = io_inValid_25 & _T_5219; // @[Switch.scala 30:36:@410.4]
  assign _T_5222 = io_inAddr_26 == 5'h2; // @[Switch.scala 30:53:@412.4]
  assign valid_2_26 = io_inValid_26 & _T_5222; // @[Switch.scala 30:36:@413.4]
  assign _T_5225 = io_inAddr_27 == 5'h2; // @[Switch.scala 30:53:@415.4]
  assign valid_2_27 = io_inValid_27 & _T_5225; // @[Switch.scala 30:36:@416.4]
  assign _T_5228 = io_inAddr_28 == 5'h2; // @[Switch.scala 30:53:@418.4]
  assign valid_2_28 = io_inValid_28 & _T_5228; // @[Switch.scala 30:36:@419.4]
  assign _T_5231 = io_inAddr_29 == 5'h2; // @[Switch.scala 30:53:@421.4]
  assign valid_2_29 = io_inValid_29 & _T_5231; // @[Switch.scala 30:36:@422.4]
  assign _T_5234 = io_inAddr_30 == 5'h2; // @[Switch.scala 30:53:@424.4]
  assign valid_2_30 = io_inValid_30 & _T_5234; // @[Switch.scala 30:36:@425.4]
  assign _T_5237 = io_inAddr_31 == 5'h2; // @[Switch.scala 30:53:@427.4]
  assign valid_2_31 = io_inValid_31 & _T_5237; // @[Switch.scala 30:36:@428.4]
  assign _T_5271 = valid_2_30 ? 5'h1e : 5'h1f; // @[Mux.scala 31:69:@430.4]
  assign _T_5272 = valid_2_29 ? 5'h1d : _T_5271; // @[Mux.scala 31:69:@431.4]
  assign _T_5273 = valid_2_28 ? 5'h1c : _T_5272; // @[Mux.scala 31:69:@432.4]
  assign _T_5274 = valid_2_27 ? 5'h1b : _T_5273; // @[Mux.scala 31:69:@433.4]
  assign _T_5275 = valid_2_26 ? 5'h1a : _T_5274; // @[Mux.scala 31:69:@434.4]
  assign _T_5276 = valid_2_25 ? 5'h19 : _T_5275; // @[Mux.scala 31:69:@435.4]
  assign _T_5277 = valid_2_24 ? 5'h18 : _T_5276; // @[Mux.scala 31:69:@436.4]
  assign _T_5278 = valid_2_23 ? 5'h17 : _T_5277; // @[Mux.scala 31:69:@437.4]
  assign _T_5279 = valid_2_22 ? 5'h16 : _T_5278; // @[Mux.scala 31:69:@438.4]
  assign _T_5280 = valid_2_21 ? 5'h15 : _T_5279; // @[Mux.scala 31:69:@439.4]
  assign _T_5281 = valid_2_20 ? 5'h14 : _T_5280; // @[Mux.scala 31:69:@440.4]
  assign _T_5282 = valid_2_19 ? 5'h13 : _T_5281; // @[Mux.scala 31:69:@441.4]
  assign _T_5283 = valid_2_18 ? 5'h12 : _T_5282; // @[Mux.scala 31:69:@442.4]
  assign _T_5284 = valid_2_17 ? 5'h11 : _T_5283; // @[Mux.scala 31:69:@443.4]
  assign _T_5285 = valid_2_16 ? 5'h10 : _T_5284; // @[Mux.scala 31:69:@444.4]
  assign _T_5286 = valid_2_15 ? 5'hf : _T_5285; // @[Mux.scala 31:69:@445.4]
  assign _T_5287 = valid_2_14 ? 5'he : _T_5286; // @[Mux.scala 31:69:@446.4]
  assign _T_5288 = valid_2_13 ? 5'hd : _T_5287; // @[Mux.scala 31:69:@447.4]
  assign _T_5289 = valid_2_12 ? 5'hc : _T_5288; // @[Mux.scala 31:69:@448.4]
  assign _T_5290 = valid_2_11 ? 5'hb : _T_5289; // @[Mux.scala 31:69:@449.4]
  assign _T_5291 = valid_2_10 ? 5'ha : _T_5290; // @[Mux.scala 31:69:@450.4]
  assign _T_5292 = valid_2_9 ? 5'h9 : _T_5291; // @[Mux.scala 31:69:@451.4]
  assign _T_5293 = valid_2_8 ? 5'h8 : _T_5292; // @[Mux.scala 31:69:@452.4]
  assign _T_5294 = valid_2_7 ? 5'h7 : _T_5293; // @[Mux.scala 31:69:@453.4]
  assign _T_5295 = valid_2_6 ? 5'h6 : _T_5294; // @[Mux.scala 31:69:@454.4]
  assign _T_5296 = valid_2_5 ? 5'h5 : _T_5295; // @[Mux.scala 31:69:@455.4]
  assign _T_5297 = valid_2_4 ? 5'h4 : _T_5296; // @[Mux.scala 31:69:@456.4]
  assign _T_5298 = valid_2_3 ? 5'h3 : _T_5297; // @[Mux.scala 31:69:@457.4]
  assign _T_5299 = valid_2_2 ? 5'h2 : _T_5298; // @[Mux.scala 31:69:@458.4]
  assign _T_5300 = valid_2_1 ? 5'h1 : _T_5299; // @[Mux.scala 31:69:@459.4]
  assign select_2 = valid_2_0 ? 5'h0 : _T_5300; // @[Mux.scala 31:69:@460.4]
  assign _GEN_65 = 5'h1 == select_2 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@462.4]
  assign _GEN_66 = 5'h2 == select_2 ? io_inData_2 : _GEN_65; // @[Switch.scala 33:19:@462.4]
  assign _GEN_67 = 5'h3 == select_2 ? io_inData_3 : _GEN_66; // @[Switch.scala 33:19:@462.4]
  assign _GEN_68 = 5'h4 == select_2 ? io_inData_4 : _GEN_67; // @[Switch.scala 33:19:@462.4]
  assign _GEN_69 = 5'h5 == select_2 ? io_inData_5 : _GEN_68; // @[Switch.scala 33:19:@462.4]
  assign _GEN_70 = 5'h6 == select_2 ? io_inData_6 : _GEN_69; // @[Switch.scala 33:19:@462.4]
  assign _GEN_71 = 5'h7 == select_2 ? io_inData_7 : _GEN_70; // @[Switch.scala 33:19:@462.4]
  assign _GEN_72 = 5'h8 == select_2 ? io_inData_8 : _GEN_71; // @[Switch.scala 33:19:@462.4]
  assign _GEN_73 = 5'h9 == select_2 ? io_inData_9 : _GEN_72; // @[Switch.scala 33:19:@462.4]
  assign _GEN_74 = 5'ha == select_2 ? io_inData_10 : _GEN_73; // @[Switch.scala 33:19:@462.4]
  assign _GEN_75 = 5'hb == select_2 ? io_inData_11 : _GEN_74; // @[Switch.scala 33:19:@462.4]
  assign _GEN_76 = 5'hc == select_2 ? io_inData_12 : _GEN_75; // @[Switch.scala 33:19:@462.4]
  assign _GEN_77 = 5'hd == select_2 ? io_inData_13 : _GEN_76; // @[Switch.scala 33:19:@462.4]
  assign _GEN_78 = 5'he == select_2 ? io_inData_14 : _GEN_77; // @[Switch.scala 33:19:@462.4]
  assign _GEN_79 = 5'hf == select_2 ? io_inData_15 : _GEN_78; // @[Switch.scala 33:19:@462.4]
  assign _GEN_80 = 5'h10 == select_2 ? io_inData_16 : _GEN_79; // @[Switch.scala 33:19:@462.4]
  assign _GEN_81 = 5'h11 == select_2 ? io_inData_17 : _GEN_80; // @[Switch.scala 33:19:@462.4]
  assign _GEN_82 = 5'h12 == select_2 ? io_inData_18 : _GEN_81; // @[Switch.scala 33:19:@462.4]
  assign _GEN_83 = 5'h13 == select_2 ? io_inData_19 : _GEN_82; // @[Switch.scala 33:19:@462.4]
  assign _GEN_84 = 5'h14 == select_2 ? io_inData_20 : _GEN_83; // @[Switch.scala 33:19:@462.4]
  assign _GEN_85 = 5'h15 == select_2 ? io_inData_21 : _GEN_84; // @[Switch.scala 33:19:@462.4]
  assign _GEN_86 = 5'h16 == select_2 ? io_inData_22 : _GEN_85; // @[Switch.scala 33:19:@462.4]
  assign _GEN_87 = 5'h17 == select_2 ? io_inData_23 : _GEN_86; // @[Switch.scala 33:19:@462.4]
  assign _GEN_88 = 5'h18 == select_2 ? io_inData_24 : _GEN_87; // @[Switch.scala 33:19:@462.4]
  assign _GEN_89 = 5'h19 == select_2 ? io_inData_25 : _GEN_88; // @[Switch.scala 33:19:@462.4]
  assign _GEN_90 = 5'h1a == select_2 ? io_inData_26 : _GEN_89; // @[Switch.scala 33:19:@462.4]
  assign _GEN_91 = 5'h1b == select_2 ? io_inData_27 : _GEN_90; // @[Switch.scala 33:19:@462.4]
  assign _GEN_92 = 5'h1c == select_2 ? io_inData_28 : _GEN_91; // @[Switch.scala 33:19:@462.4]
  assign _GEN_93 = 5'h1d == select_2 ? io_inData_29 : _GEN_92; // @[Switch.scala 33:19:@462.4]
  assign _GEN_94 = 5'h1e == select_2 ? io_inData_30 : _GEN_93; // @[Switch.scala 33:19:@462.4]
  assign _T_5309 = {valid_2_7,valid_2_6,valid_2_5,valid_2_4,valid_2_3,valid_2_2,valid_2_1,valid_2_0}; // @[Switch.scala 34:32:@469.4]
  assign _T_5317 = {valid_2_15,valid_2_14,valid_2_13,valid_2_12,valid_2_11,valid_2_10,valid_2_9,valid_2_8,_T_5309}; // @[Switch.scala 34:32:@477.4]
  assign _T_5324 = {valid_2_23,valid_2_22,valid_2_21,valid_2_20,valid_2_19,valid_2_18,valid_2_17,valid_2_16}; // @[Switch.scala 34:32:@484.4]
  assign _T_5333 = {valid_2_31,valid_2_30,valid_2_29,valid_2_28,valid_2_27,valid_2_26,valid_2_25,valid_2_24,_T_5324,_T_5317}; // @[Switch.scala 34:32:@493.4]
  assign _T_5337 = io_inAddr_0 == 5'h3; // @[Switch.scala 30:53:@496.4]
  assign valid_3_0 = io_inValid_0 & _T_5337; // @[Switch.scala 30:36:@497.4]
  assign _T_5340 = io_inAddr_1 == 5'h3; // @[Switch.scala 30:53:@499.4]
  assign valid_3_1 = io_inValid_1 & _T_5340; // @[Switch.scala 30:36:@500.4]
  assign _T_5343 = io_inAddr_2 == 5'h3; // @[Switch.scala 30:53:@502.4]
  assign valid_3_2 = io_inValid_2 & _T_5343; // @[Switch.scala 30:36:@503.4]
  assign _T_5346 = io_inAddr_3 == 5'h3; // @[Switch.scala 30:53:@505.4]
  assign valid_3_3 = io_inValid_3 & _T_5346; // @[Switch.scala 30:36:@506.4]
  assign _T_5349 = io_inAddr_4 == 5'h3; // @[Switch.scala 30:53:@508.4]
  assign valid_3_4 = io_inValid_4 & _T_5349; // @[Switch.scala 30:36:@509.4]
  assign _T_5352 = io_inAddr_5 == 5'h3; // @[Switch.scala 30:53:@511.4]
  assign valid_3_5 = io_inValid_5 & _T_5352; // @[Switch.scala 30:36:@512.4]
  assign _T_5355 = io_inAddr_6 == 5'h3; // @[Switch.scala 30:53:@514.4]
  assign valid_3_6 = io_inValid_6 & _T_5355; // @[Switch.scala 30:36:@515.4]
  assign _T_5358 = io_inAddr_7 == 5'h3; // @[Switch.scala 30:53:@517.4]
  assign valid_3_7 = io_inValid_7 & _T_5358; // @[Switch.scala 30:36:@518.4]
  assign _T_5361 = io_inAddr_8 == 5'h3; // @[Switch.scala 30:53:@520.4]
  assign valid_3_8 = io_inValid_8 & _T_5361; // @[Switch.scala 30:36:@521.4]
  assign _T_5364 = io_inAddr_9 == 5'h3; // @[Switch.scala 30:53:@523.4]
  assign valid_3_9 = io_inValid_9 & _T_5364; // @[Switch.scala 30:36:@524.4]
  assign _T_5367 = io_inAddr_10 == 5'h3; // @[Switch.scala 30:53:@526.4]
  assign valid_3_10 = io_inValid_10 & _T_5367; // @[Switch.scala 30:36:@527.4]
  assign _T_5370 = io_inAddr_11 == 5'h3; // @[Switch.scala 30:53:@529.4]
  assign valid_3_11 = io_inValid_11 & _T_5370; // @[Switch.scala 30:36:@530.4]
  assign _T_5373 = io_inAddr_12 == 5'h3; // @[Switch.scala 30:53:@532.4]
  assign valid_3_12 = io_inValid_12 & _T_5373; // @[Switch.scala 30:36:@533.4]
  assign _T_5376 = io_inAddr_13 == 5'h3; // @[Switch.scala 30:53:@535.4]
  assign valid_3_13 = io_inValid_13 & _T_5376; // @[Switch.scala 30:36:@536.4]
  assign _T_5379 = io_inAddr_14 == 5'h3; // @[Switch.scala 30:53:@538.4]
  assign valid_3_14 = io_inValid_14 & _T_5379; // @[Switch.scala 30:36:@539.4]
  assign _T_5382 = io_inAddr_15 == 5'h3; // @[Switch.scala 30:53:@541.4]
  assign valid_3_15 = io_inValid_15 & _T_5382; // @[Switch.scala 30:36:@542.4]
  assign _T_5385 = io_inAddr_16 == 5'h3; // @[Switch.scala 30:53:@544.4]
  assign valid_3_16 = io_inValid_16 & _T_5385; // @[Switch.scala 30:36:@545.4]
  assign _T_5388 = io_inAddr_17 == 5'h3; // @[Switch.scala 30:53:@547.4]
  assign valid_3_17 = io_inValid_17 & _T_5388; // @[Switch.scala 30:36:@548.4]
  assign _T_5391 = io_inAddr_18 == 5'h3; // @[Switch.scala 30:53:@550.4]
  assign valid_3_18 = io_inValid_18 & _T_5391; // @[Switch.scala 30:36:@551.4]
  assign _T_5394 = io_inAddr_19 == 5'h3; // @[Switch.scala 30:53:@553.4]
  assign valid_3_19 = io_inValid_19 & _T_5394; // @[Switch.scala 30:36:@554.4]
  assign _T_5397 = io_inAddr_20 == 5'h3; // @[Switch.scala 30:53:@556.4]
  assign valid_3_20 = io_inValid_20 & _T_5397; // @[Switch.scala 30:36:@557.4]
  assign _T_5400 = io_inAddr_21 == 5'h3; // @[Switch.scala 30:53:@559.4]
  assign valid_3_21 = io_inValid_21 & _T_5400; // @[Switch.scala 30:36:@560.4]
  assign _T_5403 = io_inAddr_22 == 5'h3; // @[Switch.scala 30:53:@562.4]
  assign valid_3_22 = io_inValid_22 & _T_5403; // @[Switch.scala 30:36:@563.4]
  assign _T_5406 = io_inAddr_23 == 5'h3; // @[Switch.scala 30:53:@565.4]
  assign valid_3_23 = io_inValid_23 & _T_5406; // @[Switch.scala 30:36:@566.4]
  assign _T_5409 = io_inAddr_24 == 5'h3; // @[Switch.scala 30:53:@568.4]
  assign valid_3_24 = io_inValid_24 & _T_5409; // @[Switch.scala 30:36:@569.4]
  assign _T_5412 = io_inAddr_25 == 5'h3; // @[Switch.scala 30:53:@571.4]
  assign valid_3_25 = io_inValid_25 & _T_5412; // @[Switch.scala 30:36:@572.4]
  assign _T_5415 = io_inAddr_26 == 5'h3; // @[Switch.scala 30:53:@574.4]
  assign valid_3_26 = io_inValid_26 & _T_5415; // @[Switch.scala 30:36:@575.4]
  assign _T_5418 = io_inAddr_27 == 5'h3; // @[Switch.scala 30:53:@577.4]
  assign valid_3_27 = io_inValid_27 & _T_5418; // @[Switch.scala 30:36:@578.4]
  assign _T_5421 = io_inAddr_28 == 5'h3; // @[Switch.scala 30:53:@580.4]
  assign valid_3_28 = io_inValid_28 & _T_5421; // @[Switch.scala 30:36:@581.4]
  assign _T_5424 = io_inAddr_29 == 5'h3; // @[Switch.scala 30:53:@583.4]
  assign valid_3_29 = io_inValid_29 & _T_5424; // @[Switch.scala 30:36:@584.4]
  assign _T_5427 = io_inAddr_30 == 5'h3; // @[Switch.scala 30:53:@586.4]
  assign valid_3_30 = io_inValid_30 & _T_5427; // @[Switch.scala 30:36:@587.4]
  assign _T_5430 = io_inAddr_31 == 5'h3; // @[Switch.scala 30:53:@589.4]
  assign valid_3_31 = io_inValid_31 & _T_5430; // @[Switch.scala 30:36:@590.4]
  assign _T_5464 = valid_3_30 ? 5'h1e : 5'h1f; // @[Mux.scala 31:69:@592.4]
  assign _T_5465 = valid_3_29 ? 5'h1d : _T_5464; // @[Mux.scala 31:69:@593.4]
  assign _T_5466 = valid_3_28 ? 5'h1c : _T_5465; // @[Mux.scala 31:69:@594.4]
  assign _T_5467 = valid_3_27 ? 5'h1b : _T_5466; // @[Mux.scala 31:69:@595.4]
  assign _T_5468 = valid_3_26 ? 5'h1a : _T_5467; // @[Mux.scala 31:69:@596.4]
  assign _T_5469 = valid_3_25 ? 5'h19 : _T_5468; // @[Mux.scala 31:69:@597.4]
  assign _T_5470 = valid_3_24 ? 5'h18 : _T_5469; // @[Mux.scala 31:69:@598.4]
  assign _T_5471 = valid_3_23 ? 5'h17 : _T_5470; // @[Mux.scala 31:69:@599.4]
  assign _T_5472 = valid_3_22 ? 5'h16 : _T_5471; // @[Mux.scala 31:69:@600.4]
  assign _T_5473 = valid_3_21 ? 5'h15 : _T_5472; // @[Mux.scala 31:69:@601.4]
  assign _T_5474 = valid_3_20 ? 5'h14 : _T_5473; // @[Mux.scala 31:69:@602.4]
  assign _T_5475 = valid_3_19 ? 5'h13 : _T_5474; // @[Mux.scala 31:69:@603.4]
  assign _T_5476 = valid_3_18 ? 5'h12 : _T_5475; // @[Mux.scala 31:69:@604.4]
  assign _T_5477 = valid_3_17 ? 5'h11 : _T_5476; // @[Mux.scala 31:69:@605.4]
  assign _T_5478 = valid_3_16 ? 5'h10 : _T_5477; // @[Mux.scala 31:69:@606.4]
  assign _T_5479 = valid_3_15 ? 5'hf : _T_5478; // @[Mux.scala 31:69:@607.4]
  assign _T_5480 = valid_3_14 ? 5'he : _T_5479; // @[Mux.scala 31:69:@608.4]
  assign _T_5481 = valid_3_13 ? 5'hd : _T_5480; // @[Mux.scala 31:69:@609.4]
  assign _T_5482 = valid_3_12 ? 5'hc : _T_5481; // @[Mux.scala 31:69:@610.4]
  assign _T_5483 = valid_3_11 ? 5'hb : _T_5482; // @[Mux.scala 31:69:@611.4]
  assign _T_5484 = valid_3_10 ? 5'ha : _T_5483; // @[Mux.scala 31:69:@612.4]
  assign _T_5485 = valid_3_9 ? 5'h9 : _T_5484; // @[Mux.scala 31:69:@613.4]
  assign _T_5486 = valid_3_8 ? 5'h8 : _T_5485; // @[Mux.scala 31:69:@614.4]
  assign _T_5487 = valid_3_7 ? 5'h7 : _T_5486; // @[Mux.scala 31:69:@615.4]
  assign _T_5488 = valid_3_6 ? 5'h6 : _T_5487; // @[Mux.scala 31:69:@616.4]
  assign _T_5489 = valid_3_5 ? 5'h5 : _T_5488; // @[Mux.scala 31:69:@617.4]
  assign _T_5490 = valid_3_4 ? 5'h4 : _T_5489; // @[Mux.scala 31:69:@618.4]
  assign _T_5491 = valid_3_3 ? 5'h3 : _T_5490; // @[Mux.scala 31:69:@619.4]
  assign _T_5492 = valid_3_2 ? 5'h2 : _T_5491; // @[Mux.scala 31:69:@620.4]
  assign _T_5493 = valid_3_1 ? 5'h1 : _T_5492; // @[Mux.scala 31:69:@621.4]
  assign select_3 = valid_3_0 ? 5'h0 : _T_5493; // @[Mux.scala 31:69:@622.4]
  assign _GEN_97 = 5'h1 == select_3 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@624.4]
  assign _GEN_98 = 5'h2 == select_3 ? io_inData_2 : _GEN_97; // @[Switch.scala 33:19:@624.4]
  assign _GEN_99 = 5'h3 == select_3 ? io_inData_3 : _GEN_98; // @[Switch.scala 33:19:@624.4]
  assign _GEN_100 = 5'h4 == select_3 ? io_inData_4 : _GEN_99; // @[Switch.scala 33:19:@624.4]
  assign _GEN_101 = 5'h5 == select_3 ? io_inData_5 : _GEN_100; // @[Switch.scala 33:19:@624.4]
  assign _GEN_102 = 5'h6 == select_3 ? io_inData_6 : _GEN_101; // @[Switch.scala 33:19:@624.4]
  assign _GEN_103 = 5'h7 == select_3 ? io_inData_7 : _GEN_102; // @[Switch.scala 33:19:@624.4]
  assign _GEN_104 = 5'h8 == select_3 ? io_inData_8 : _GEN_103; // @[Switch.scala 33:19:@624.4]
  assign _GEN_105 = 5'h9 == select_3 ? io_inData_9 : _GEN_104; // @[Switch.scala 33:19:@624.4]
  assign _GEN_106 = 5'ha == select_3 ? io_inData_10 : _GEN_105; // @[Switch.scala 33:19:@624.4]
  assign _GEN_107 = 5'hb == select_3 ? io_inData_11 : _GEN_106; // @[Switch.scala 33:19:@624.4]
  assign _GEN_108 = 5'hc == select_3 ? io_inData_12 : _GEN_107; // @[Switch.scala 33:19:@624.4]
  assign _GEN_109 = 5'hd == select_3 ? io_inData_13 : _GEN_108; // @[Switch.scala 33:19:@624.4]
  assign _GEN_110 = 5'he == select_3 ? io_inData_14 : _GEN_109; // @[Switch.scala 33:19:@624.4]
  assign _GEN_111 = 5'hf == select_3 ? io_inData_15 : _GEN_110; // @[Switch.scala 33:19:@624.4]
  assign _GEN_112 = 5'h10 == select_3 ? io_inData_16 : _GEN_111; // @[Switch.scala 33:19:@624.4]
  assign _GEN_113 = 5'h11 == select_3 ? io_inData_17 : _GEN_112; // @[Switch.scala 33:19:@624.4]
  assign _GEN_114 = 5'h12 == select_3 ? io_inData_18 : _GEN_113; // @[Switch.scala 33:19:@624.4]
  assign _GEN_115 = 5'h13 == select_3 ? io_inData_19 : _GEN_114; // @[Switch.scala 33:19:@624.4]
  assign _GEN_116 = 5'h14 == select_3 ? io_inData_20 : _GEN_115; // @[Switch.scala 33:19:@624.4]
  assign _GEN_117 = 5'h15 == select_3 ? io_inData_21 : _GEN_116; // @[Switch.scala 33:19:@624.4]
  assign _GEN_118 = 5'h16 == select_3 ? io_inData_22 : _GEN_117; // @[Switch.scala 33:19:@624.4]
  assign _GEN_119 = 5'h17 == select_3 ? io_inData_23 : _GEN_118; // @[Switch.scala 33:19:@624.4]
  assign _GEN_120 = 5'h18 == select_3 ? io_inData_24 : _GEN_119; // @[Switch.scala 33:19:@624.4]
  assign _GEN_121 = 5'h19 == select_3 ? io_inData_25 : _GEN_120; // @[Switch.scala 33:19:@624.4]
  assign _GEN_122 = 5'h1a == select_3 ? io_inData_26 : _GEN_121; // @[Switch.scala 33:19:@624.4]
  assign _GEN_123 = 5'h1b == select_3 ? io_inData_27 : _GEN_122; // @[Switch.scala 33:19:@624.4]
  assign _GEN_124 = 5'h1c == select_3 ? io_inData_28 : _GEN_123; // @[Switch.scala 33:19:@624.4]
  assign _GEN_125 = 5'h1d == select_3 ? io_inData_29 : _GEN_124; // @[Switch.scala 33:19:@624.4]
  assign _GEN_126 = 5'h1e == select_3 ? io_inData_30 : _GEN_125; // @[Switch.scala 33:19:@624.4]
  assign _T_5502 = {valid_3_7,valid_3_6,valid_3_5,valid_3_4,valid_3_3,valid_3_2,valid_3_1,valid_3_0}; // @[Switch.scala 34:32:@631.4]
  assign _T_5510 = {valid_3_15,valid_3_14,valid_3_13,valid_3_12,valid_3_11,valid_3_10,valid_3_9,valid_3_8,_T_5502}; // @[Switch.scala 34:32:@639.4]
  assign _T_5517 = {valid_3_23,valid_3_22,valid_3_21,valid_3_20,valid_3_19,valid_3_18,valid_3_17,valid_3_16}; // @[Switch.scala 34:32:@646.4]
  assign _T_5526 = {valid_3_31,valid_3_30,valid_3_29,valid_3_28,valid_3_27,valid_3_26,valid_3_25,valid_3_24,_T_5517,_T_5510}; // @[Switch.scala 34:32:@655.4]
  assign _T_5530 = io_inAddr_0 == 5'h4; // @[Switch.scala 30:53:@658.4]
  assign valid_4_0 = io_inValid_0 & _T_5530; // @[Switch.scala 30:36:@659.4]
  assign _T_5533 = io_inAddr_1 == 5'h4; // @[Switch.scala 30:53:@661.4]
  assign valid_4_1 = io_inValid_1 & _T_5533; // @[Switch.scala 30:36:@662.4]
  assign _T_5536 = io_inAddr_2 == 5'h4; // @[Switch.scala 30:53:@664.4]
  assign valid_4_2 = io_inValid_2 & _T_5536; // @[Switch.scala 30:36:@665.4]
  assign _T_5539 = io_inAddr_3 == 5'h4; // @[Switch.scala 30:53:@667.4]
  assign valid_4_3 = io_inValid_3 & _T_5539; // @[Switch.scala 30:36:@668.4]
  assign _T_5542 = io_inAddr_4 == 5'h4; // @[Switch.scala 30:53:@670.4]
  assign valid_4_4 = io_inValid_4 & _T_5542; // @[Switch.scala 30:36:@671.4]
  assign _T_5545 = io_inAddr_5 == 5'h4; // @[Switch.scala 30:53:@673.4]
  assign valid_4_5 = io_inValid_5 & _T_5545; // @[Switch.scala 30:36:@674.4]
  assign _T_5548 = io_inAddr_6 == 5'h4; // @[Switch.scala 30:53:@676.4]
  assign valid_4_6 = io_inValid_6 & _T_5548; // @[Switch.scala 30:36:@677.4]
  assign _T_5551 = io_inAddr_7 == 5'h4; // @[Switch.scala 30:53:@679.4]
  assign valid_4_7 = io_inValid_7 & _T_5551; // @[Switch.scala 30:36:@680.4]
  assign _T_5554 = io_inAddr_8 == 5'h4; // @[Switch.scala 30:53:@682.4]
  assign valid_4_8 = io_inValid_8 & _T_5554; // @[Switch.scala 30:36:@683.4]
  assign _T_5557 = io_inAddr_9 == 5'h4; // @[Switch.scala 30:53:@685.4]
  assign valid_4_9 = io_inValid_9 & _T_5557; // @[Switch.scala 30:36:@686.4]
  assign _T_5560 = io_inAddr_10 == 5'h4; // @[Switch.scala 30:53:@688.4]
  assign valid_4_10 = io_inValid_10 & _T_5560; // @[Switch.scala 30:36:@689.4]
  assign _T_5563 = io_inAddr_11 == 5'h4; // @[Switch.scala 30:53:@691.4]
  assign valid_4_11 = io_inValid_11 & _T_5563; // @[Switch.scala 30:36:@692.4]
  assign _T_5566 = io_inAddr_12 == 5'h4; // @[Switch.scala 30:53:@694.4]
  assign valid_4_12 = io_inValid_12 & _T_5566; // @[Switch.scala 30:36:@695.4]
  assign _T_5569 = io_inAddr_13 == 5'h4; // @[Switch.scala 30:53:@697.4]
  assign valid_4_13 = io_inValid_13 & _T_5569; // @[Switch.scala 30:36:@698.4]
  assign _T_5572 = io_inAddr_14 == 5'h4; // @[Switch.scala 30:53:@700.4]
  assign valid_4_14 = io_inValid_14 & _T_5572; // @[Switch.scala 30:36:@701.4]
  assign _T_5575 = io_inAddr_15 == 5'h4; // @[Switch.scala 30:53:@703.4]
  assign valid_4_15 = io_inValid_15 & _T_5575; // @[Switch.scala 30:36:@704.4]
  assign _T_5578 = io_inAddr_16 == 5'h4; // @[Switch.scala 30:53:@706.4]
  assign valid_4_16 = io_inValid_16 & _T_5578; // @[Switch.scala 30:36:@707.4]
  assign _T_5581 = io_inAddr_17 == 5'h4; // @[Switch.scala 30:53:@709.4]
  assign valid_4_17 = io_inValid_17 & _T_5581; // @[Switch.scala 30:36:@710.4]
  assign _T_5584 = io_inAddr_18 == 5'h4; // @[Switch.scala 30:53:@712.4]
  assign valid_4_18 = io_inValid_18 & _T_5584; // @[Switch.scala 30:36:@713.4]
  assign _T_5587 = io_inAddr_19 == 5'h4; // @[Switch.scala 30:53:@715.4]
  assign valid_4_19 = io_inValid_19 & _T_5587; // @[Switch.scala 30:36:@716.4]
  assign _T_5590 = io_inAddr_20 == 5'h4; // @[Switch.scala 30:53:@718.4]
  assign valid_4_20 = io_inValid_20 & _T_5590; // @[Switch.scala 30:36:@719.4]
  assign _T_5593 = io_inAddr_21 == 5'h4; // @[Switch.scala 30:53:@721.4]
  assign valid_4_21 = io_inValid_21 & _T_5593; // @[Switch.scala 30:36:@722.4]
  assign _T_5596 = io_inAddr_22 == 5'h4; // @[Switch.scala 30:53:@724.4]
  assign valid_4_22 = io_inValid_22 & _T_5596; // @[Switch.scala 30:36:@725.4]
  assign _T_5599 = io_inAddr_23 == 5'h4; // @[Switch.scala 30:53:@727.4]
  assign valid_4_23 = io_inValid_23 & _T_5599; // @[Switch.scala 30:36:@728.4]
  assign _T_5602 = io_inAddr_24 == 5'h4; // @[Switch.scala 30:53:@730.4]
  assign valid_4_24 = io_inValid_24 & _T_5602; // @[Switch.scala 30:36:@731.4]
  assign _T_5605 = io_inAddr_25 == 5'h4; // @[Switch.scala 30:53:@733.4]
  assign valid_4_25 = io_inValid_25 & _T_5605; // @[Switch.scala 30:36:@734.4]
  assign _T_5608 = io_inAddr_26 == 5'h4; // @[Switch.scala 30:53:@736.4]
  assign valid_4_26 = io_inValid_26 & _T_5608; // @[Switch.scala 30:36:@737.4]
  assign _T_5611 = io_inAddr_27 == 5'h4; // @[Switch.scala 30:53:@739.4]
  assign valid_4_27 = io_inValid_27 & _T_5611; // @[Switch.scala 30:36:@740.4]
  assign _T_5614 = io_inAddr_28 == 5'h4; // @[Switch.scala 30:53:@742.4]
  assign valid_4_28 = io_inValid_28 & _T_5614; // @[Switch.scala 30:36:@743.4]
  assign _T_5617 = io_inAddr_29 == 5'h4; // @[Switch.scala 30:53:@745.4]
  assign valid_4_29 = io_inValid_29 & _T_5617; // @[Switch.scala 30:36:@746.4]
  assign _T_5620 = io_inAddr_30 == 5'h4; // @[Switch.scala 30:53:@748.4]
  assign valid_4_30 = io_inValid_30 & _T_5620; // @[Switch.scala 30:36:@749.4]
  assign _T_5623 = io_inAddr_31 == 5'h4; // @[Switch.scala 30:53:@751.4]
  assign valid_4_31 = io_inValid_31 & _T_5623; // @[Switch.scala 30:36:@752.4]
  assign _T_5657 = valid_4_30 ? 5'h1e : 5'h1f; // @[Mux.scala 31:69:@754.4]
  assign _T_5658 = valid_4_29 ? 5'h1d : _T_5657; // @[Mux.scala 31:69:@755.4]
  assign _T_5659 = valid_4_28 ? 5'h1c : _T_5658; // @[Mux.scala 31:69:@756.4]
  assign _T_5660 = valid_4_27 ? 5'h1b : _T_5659; // @[Mux.scala 31:69:@757.4]
  assign _T_5661 = valid_4_26 ? 5'h1a : _T_5660; // @[Mux.scala 31:69:@758.4]
  assign _T_5662 = valid_4_25 ? 5'h19 : _T_5661; // @[Mux.scala 31:69:@759.4]
  assign _T_5663 = valid_4_24 ? 5'h18 : _T_5662; // @[Mux.scala 31:69:@760.4]
  assign _T_5664 = valid_4_23 ? 5'h17 : _T_5663; // @[Mux.scala 31:69:@761.4]
  assign _T_5665 = valid_4_22 ? 5'h16 : _T_5664; // @[Mux.scala 31:69:@762.4]
  assign _T_5666 = valid_4_21 ? 5'h15 : _T_5665; // @[Mux.scala 31:69:@763.4]
  assign _T_5667 = valid_4_20 ? 5'h14 : _T_5666; // @[Mux.scala 31:69:@764.4]
  assign _T_5668 = valid_4_19 ? 5'h13 : _T_5667; // @[Mux.scala 31:69:@765.4]
  assign _T_5669 = valid_4_18 ? 5'h12 : _T_5668; // @[Mux.scala 31:69:@766.4]
  assign _T_5670 = valid_4_17 ? 5'h11 : _T_5669; // @[Mux.scala 31:69:@767.4]
  assign _T_5671 = valid_4_16 ? 5'h10 : _T_5670; // @[Mux.scala 31:69:@768.4]
  assign _T_5672 = valid_4_15 ? 5'hf : _T_5671; // @[Mux.scala 31:69:@769.4]
  assign _T_5673 = valid_4_14 ? 5'he : _T_5672; // @[Mux.scala 31:69:@770.4]
  assign _T_5674 = valid_4_13 ? 5'hd : _T_5673; // @[Mux.scala 31:69:@771.4]
  assign _T_5675 = valid_4_12 ? 5'hc : _T_5674; // @[Mux.scala 31:69:@772.4]
  assign _T_5676 = valid_4_11 ? 5'hb : _T_5675; // @[Mux.scala 31:69:@773.4]
  assign _T_5677 = valid_4_10 ? 5'ha : _T_5676; // @[Mux.scala 31:69:@774.4]
  assign _T_5678 = valid_4_9 ? 5'h9 : _T_5677; // @[Mux.scala 31:69:@775.4]
  assign _T_5679 = valid_4_8 ? 5'h8 : _T_5678; // @[Mux.scala 31:69:@776.4]
  assign _T_5680 = valid_4_7 ? 5'h7 : _T_5679; // @[Mux.scala 31:69:@777.4]
  assign _T_5681 = valid_4_6 ? 5'h6 : _T_5680; // @[Mux.scala 31:69:@778.4]
  assign _T_5682 = valid_4_5 ? 5'h5 : _T_5681; // @[Mux.scala 31:69:@779.4]
  assign _T_5683 = valid_4_4 ? 5'h4 : _T_5682; // @[Mux.scala 31:69:@780.4]
  assign _T_5684 = valid_4_3 ? 5'h3 : _T_5683; // @[Mux.scala 31:69:@781.4]
  assign _T_5685 = valid_4_2 ? 5'h2 : _T_5684; // @[Mux.scala 31:69:@782.4]
  assign _T_5686 = valid_4_1 ? 5'h1 : _T_5685; // @[Mux.scala 31:69:@783.4]
  assign select_4 = valid_4_0 ? 5'h0 : _T_5686; // @[Mux.scala 31:69:@784.4]
  assign _GEN_129 = 5'h1 == select_4 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@786.4]
  assign _GEN_130 = 5'h2 == select_4 ? io_inData_2 : _GEN_129; // @[Switch.scala 33:19:@786.4]
  assign _GEN_131 = 5'h3 == select_4 ? io_inData_3 : _GEN_130; // @[Switch.scala 33:19:@786.4]
  assign _GEN_132 = 5'h4 == select_4 ? io_inData_4 : _GEN_131; // @[Switch.scala 33:19:@786.4]
  assign _GEN_133 = 5'h5 == select_4 ? io_inData_5 : _GEN_132; // @[Switch.scala 33:19:@786.4]
  assign _GEN_134 = 5'h6 == select_4 ? io_inData_6 : _GEN_133; // @[Switch.scala 33:19:@786.4]
  assign _GEN_135 = 5'h7 == select_4 ? io_inData_7 : _GEN_134; // @[Switch.scala 33:19:@786.4]
  assign _GEN_136 = 5'h8 == select_4 ? io_inData_8 : _GEN_135; // @[Switch.scala 33:19:@786.4]
  assign _GEN_137 = 5'h9 == select_4 ? io_inData_9 : _GEN_136; // @[Switch.scala 33:19:@786.4]
  assign _GEN_138 = 5'ha == select_4 ? io_inData_10 : _GEN_137; // @[Switch.scala 33:19:@786.4]
  assign _GEN_139 = 5'hb == select_4 ? io_inData_11 : _GEN_138; // @[Switch.scala 33:19:@786.4]
  assign _GEN_140 = 5'hc == select_4 ? io_inData_12 : _GEN_139; // @[Switch.scala 33:19:@786.4]
  assign _GEN_141 = 5'hd == select_4 ? io_inData_13 : _GEN_140; // @[Switch.scala 33:19:@786.4]
  assign _GEN_142 = 5'he == select_4 ? io_inData_14 : _GEN_141; // @[Switch.scala 33:19:@786.4]
  assign _GEN_143 = 5'hf == select_4 ? io_inData_15 : _GEN_142; // @[Switch.scala 33:19:@786.4]
  assign _GEN_144 = 5'h10 == select_4 ? io_inData_16 : _GEN_143; // @[Switch.scala 33:19:@786.4]
  assign _GEN_145 = 5'h11 == select_4 ? io_inData_17 : _GEN_144; // @[Switch.scala 33:19:@786.4]
  assign _GEN_146 = 5'h12 == select_4 ? io_inData_18 : _GEN_145; // @[Switch.scala 33:19:@786.4]
  assign _GEN_147 = 5'h13 == select_4 ? io_inData_19 : _GEN_146; // @[Switch.scala 33:19:@786.4]
  assign _GEN_148 = 5'h14 == select_4 ? io_inData_20 : _GEN_147; // @[Switch.scala 33:19:@786.4]
  assign _GEN_149 = 5'h15 == select_4 ? io_inData_21 : _GEN_148; // @[Switch.scala 33:19:@786.4]
  assign _GEN_150 = 5'h16 == select_4 ? io_inData_22 : _GEN_149; // @[Switch.scala 33:19:@786.4]
  assign _GEN_151 = 5'h17 == select_4 ? io_inData_23 : _GEN_150; // @[Switch.scala 33:19:@786.4]
  assign _GEN_152 = 5'h18 == select_4 ? io_inData_24 : _GEN_151; // @[Switch.scala 33:19:@786.4]
  assign _GEN_153 = 5'h19 == select_4 ? io_inData_25 : _GEN_152; // @[Switch.scala 33:19:@786.4]
  assign _GEN_154 = 5'h1a == select_4 ? io_inData_26 : _GEN_153; // @[Switch.scala 33:19:@786.4]
  assign _GEN_155 = 5'h1b == select_4 ? io_inData_27 : _GEN_154; // @[Switch.scala 33:19:@786.4]
  assign _GEN_156 = 5'h1c == select_4 ? io_inData_28 : _GEN_155; // @[Switch.scala 33:19:@786.4]
  assign _GEN_157 = 5'h1d == select_4 ? io_inData_29 : _GEN_156; // @[Switch.scala 33:19:@786.4]
  assign _GEN_158 = 5'h1e == select_4 ? io_inData_30 : _GEN_157; // @[Switch.scala 33:19:@786.4]
  assign _T_5695 = {valid_4_7,valid_4_6,valid_4_5,valid_4_4,valid_4_3,valid_4_2,valid_4_1,valid_4_0}; // @[Switch.scala 34:32:@793.4]
  assign _T_5703 = {valid_4_15,valid_4_14,valid_4_13,valid_4_12,valid_4_11,valid_4_10,valid_4_9,valid_4_8,_T_5695}; // @[Switch.scala 34:32:@801.4]
  assign _T_5710 = {valid_4_23,valid_4_22,valid_4_21,valid_4_20,valid_4_19,valid_4_18,valid_4_17,valid_4_16}; // @[Switch.scala 34:32:@808.4]
  assign _T_5719 = {valid_4_31,valid_4_30,valid_4_29,valid_4_28,valid_4_27,valid_4_26,valid_4_25,valid_4_24,_T_5710,_T_5703}; // @[Switch.scala 34:32:@817.4]
  assign _T_5723 = io_inAddr_0 == 5'h5; // @[Switch.scala 30:53:@820.4]
  assign valid_5_0 = io_inValid_0 & _T_5723; // @[Switch.scala 30:36:@821.4]
  assign _T_5726 = io_inAddr_1 == 5'h5; // @[Switch.scala 30:53:@823.4]
  assign valid_5_1 = io_inValid_1 & _T_5726; // @[Switch.scala 30:36:@824.4]
  assign _T_5729 = io_inAddr_2 == 5'h5; // @[Switch.scala 30:53:@826.4]
  assign valid_5_2 = io_inValid_2 & _T_5729; // @[Switch.scala 30:36:@827.4]
  assign _T_5732 = io_inAddr_3 == 5'h5; // @[Switch.scala 30:53:@829.4]
  assign valid_5_3 = io_inValid_3 & _T_5732; // @[Switch.scala 30:36:@830.4]
  assign _T_5735 = io_inAddr_4 == 5'h5; // @[Switch.scala 30:53:@832.4]
  assign valid_5_4 = io_inValid_4 & _T_5735; // @[Switch.scala 30:36:@833.4]
  assign _T_5738 = io_inAddr_5 == 5'h5; // @[Switch.scala 30:53:@835.4]
  assign valid_5_5 = io_inValid_5 & _T_5738; // @[Switch.scala 30:36:@836.4]
  assign _T_5741 = io_inAddr_6 == 5'h5; // @[Switch.scala 30:53:@838.4]
  assign valid_5_6 = io_inValid_6 & _T_5741; // @[Switch.scala 30:36:@839.4]
  assign _T_5744 = io_inAddr_7 == 5'h5; // @[Switch.scala 30:53:@841.4]
  assign valid_5_7 = io_inValid_7 & _T_5744; // @[Switch.scala 30:36:@842.4]
  assign _T_5747 = io_inAddr_8 == 5'h5; // @[Switch.scala 30:53:@844.4]
  assign valid_5_8 = io_inValid_8 & _T_5747; // @[Switch.scala 30:36:@845.4]
  assign _T_5750 = io_inAddr_9 == 5'h5; // @[Switch.scala 30:53:@847.4]
  assign valid_5_9 = io_inValid_9 & _T_5750; // @[Switch.scala 30:36:@848.4]
  assign _T_5753 = io_inAddr_10 == 5'h5; // @[Switch.scala 30:53:@850.4]
  assign valid_5_10 = io_inValid_10 & _T_5753; // @[Switch.scala 30:36:@851.4]
  assign _T_5756 = io_inAddr_11 == 5'h5; // @[Switch.scala 30:53:@853.4]
  assign valid_5_11 = io_inValid_11 & _T_5756; // @[Switch.scala 30:36:@854.4]
  assign _T_5759 = io_inAddr_12 == 5'h5; // @[Switch.scala 30:53:@856.4]
  assign valid_5_12 = io_inValid_12 & _T_5759; // @[Switch.scala 30:36:@857.4]
  assign _T_5762 = io_inAddr_13 == 5'h5; // @[Switch.scala 30:53:@859.4]
  assign valid_5_13 = io_inValid_13 & _T_5762; // @[Switch.scala 30:36:@860.4]
  assign _T_5765 = io_inAddr_14 == 5'h5; // @[Switch.scala 30:53:@862.4]
  assign valid_5_14 = io_inValid_14 & _T_5765; // @[Switch.scala 30:36:@863.4]
  assign _T_5768 = io_inAddr_15 == 5'h5; // @[Switch.scala 30:53:@865.4]
  assign valid_5_15 = io_inValid_15 & _T_5768; // @[Switch.scala 30:36:@866.4]
  assign _T_5771 = io_inAddr_16 == 5'h5; // @[Switch.scala 30:53:@868.4]
  assign valid_5_16 = io_inValid_16 & _T_5771; // @[Switch.scala 30:36:@869.4]
  assign _T_5774 = io_inAddr_17 == 5'h5; // @[Switch.scala 30:53:@871.4]
  assign valid_5_17 = io_inValid_17 & _T_5774; // @[Switch.scala 30:36:@872.4]
  assign _T_5777 = io_inAddr_18 == 5'h5; // @[Switch.scala 30:53:@874.4]
  assign valid_5_18 = io_inValid_18 & _T_5777; // @[Switch.scala 30:36:@875.4]
  assign _T_5780 = io_inAddr_19 == 5'h5; // @[Switch.scala 30:53:@877.4]
  assign valid_5_19 = io_inValid_19 & _T_5780; // @[Switch.scala 30:36:@878.4]
  assign _T_5783 = io_inAddr_20 == 5'h5; // @[Switch.scala 30:53:@880.4]
  assign valid_5_20 = io_inValid_20 & _T_5783; // @[Switch.scala 30:36:@881.4]
  assign _T_5786 = io_inAddr_21 == 5'h5; // @[Switch.scala 30:53:@883.4]
  assign valid_5_21 = io_inValid_21 & _T_5786; // @[Switch.scala 30:36:@884.4]
  assign _T_5789 = io_inAddr_22 == 5'h5; // @[Switch.scala 30:53:@886.4]
  assign valid_5_22 = io_inValid_22 & _T_5789; // @[Switch.scala 30:36:@887.4]
  assign _T_5792 = io_inAddr_23 == 5'h5; // @[Switch.scala 30:53:@889.4]
  assign valid_5_23 = io_inValid_23 & _T_5792; // @[Switch.scala 30:36:@890.4]
  assign _T_5795 = io_inAddr_24 == 5'h5; // @[Switch.scala 30:53:@892.4]
  assign valid_5_24 = io_inValid_24 & _T_5795; // @[Switch.scala 30:36:@893.4]
  assign _T_5798 = io_inAddr_25 == 5'h5; // @[Switch.scala 30:53:@895.4]
  assign valid_5_25 = io_inValid_25 & _T_5798; // @[Switch.scala 30:36:@896.4]
  assign _T_5801 = io_inAddr_26 == 5'h5; // @[Switch.scala 30:53:@898.4]
  assign valid_5_26 = io_inValid_26 & _T_5801; // @[Switch.scala 30:36:@899.4]
  assign _T_5804 = io_inAddr_27 == 5'h5; // @[Switch.scala 30:53:@901.4]
  assign valid_5_27 = io_inValid_27 & _T_5804; // @[Switch.scala 30:36:@902.4]
  assign _T_5807 = io_inAddr_28 == 5'h5; // @[Switch.scala 30:53:@904.4]
  assign valid_5_28 = io_inValid_28 & _T_5807; // @[Switch.scala 30:36:@905.4]
  assign _T_5810 = io_inAddr_29 == 5'h5; // @[Switch.scala 30:53:@907.4]
  assign valid_5_29 = io_inValid_29 & _T_5810; // @[Switch.scala 30:36:@908.4]
  assign _T_5813 = io_inAddr_30 == 5'h5; // @[Switch.scala 30:53:@910.4]
  assign valid_5_30 = io_inValid_30 & _T_5813; // @[Switch.scala 30:36:@911.4]
  assign _T_5816 = io_inAddr_31 == 5'h5; // @[Switch.scala 30:53:@913.4]
  assign valid_5_31 = io_inValid_31 & _T_5816; // @[Switch.scala 30:36:@914.4]
  assign _T_5850 = valid_5_30 ? 5'h1e : 5'h1f; // @[Mux.scala 31:69:@916.4]
  assign _T_5851 = valid_5_29 ? 5'h1d : _T_5850; // @[Mux.scala 31:69:@917.4]
  assign _T_5852 = valid_5_28 ? 5'h1c : _T_5851; // @[Mux.scala 31:69:@918.4]
  assign _T_5853 = valid_5_27 ? 5'h1b : _T_5852; // @[Mux.scala 31:69:@919.4]
  assign _T_5854 = valid_5_26 ? 5'h1a : _T_5853; // @[Mux.scala 31:69:@920.4]
  assign _T_5855 = valid_5_25 ? 5'h19 : _T_5854; // @[Mux.scala 31:69:@921.4]
  assign _T_5856 = valid_5_24 ? 5'h18 : _T_5855; // @[Mux.scala 31:69:@922.4]
  assign _T_5857 = valid_5_23 ? 5'h17 : _T_5856; // @[Mux.scala 31:69:@923.4]
  assign _T_5858 = valid_5_22 ? 5'h16 : _T_5857; // @[Mux.scala 31:69:@924.4]
  assign _T_5859 = valid_5_21 ? 5'h15 : _T_5858; // @[Mux.scala 31:69:@925.4]
  assign _T_5860 = valid_5_20 ? 5'h14 : _T_5859; // @[Mux.scala 31:69:@926.4]
  assign _T_5861 = valid_5_19 ? 5'h13 : _T_5860; // @[Mux.scala 31:69:@927.4]
  assign _T_5862 = valid_5_18 ? 5'h12 : _T_5861; // @[Mux.scala 31:69:@928.4]
  assign _T_5863 = valid_5_17 ? 5'h11 : _T_5862; // @[Mux.scala 31:69:@929.4]
  assign _T_5864 = valid_5_16 ? 5'h10 : _T_5863; // @[Mux.scala 31:69:@930.4]
  assign _T_5865 = valid_5_15 ? 5'hf : _T_5864; // @[Mux.scala 31:69:@931.4]
  assign _T_5866 = valid_5_14 ? 5'he : _T_5865; // @[Mux.scala 31:69:@932.4]
  assign _T_5867 = valid_5_13 ? 5'hd : _T_5866; // @[Mux.scala 31:69:@933.4]
  assign _T_5868 = valid_5_12 ? 5'hc : _T_5867; // @[Mux.scala 31:69:@934.4]
  assign _T_5869 = valid_5_11 ? 5'hb : _T_5868; // @[Mux.scala 31:69:@935.4]
  assign _T_5870 = valid_5_10 ? 5'ha : _T_5869; // @[Mux.scala 31:69:@936.4]
  assign _T_5871 = valid_5_9 ? 5'h9 : _T_5870; // @[Mux.scala 31:69:@937.4]
  assign _T_5872 = valid_5_8 ? 5'h8 : _T_5871; // @[Mux.scala 31:69:@938.4]
  assign _T_5873 = valid_5_7 ? 5'h7 : _T_5872; // @[Mux.scala 31:69:@939.4]
  assign _T_5874 = valid_5_6 ? 5'h6 : _T_5873; // @[Mux.scala 31:69:@940.4]
  assign _T_5875 = valid_5_5 ? 5'h5 : _T_5874; // @[Mux.scala 31:69:@941.4]
  assign _T_5876 = valid_5_4 ? 5'h4 : _T_5875; // @[Mux.scala 31:69:@942.4]
  assign _T_5877 = valid_5_3 ? 5'h3 : _T_5876; // @[Mux.scala 31:69:@943.4]
  assign _T_5878 = valid_5_2 ? 5'h2 : _T_5877; // @[Mux.scala 31:69:@944.4]
  assign _T_5879 = valid_5_1 ? 5'h1 : _T_5878; // @[Mux.scala 31:69:@945.4]
  assign select_5 = valid_5_0 ? 5'h0 : _T_5879; // @[Mux.scala 31:69:@946.4]
  assign _GEN_161 = 5'h1 == select_5 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@948.4]
  assign _GEN_162 = 5'h2 == select_5 ? io_inData_2 : _GEN_161; // @[Switch.scala 33:19:@948.4]
  assign _GEN_163 = 5'h3 == select_5 ? io_inData_3 : _GEN_162; // @[Switch.scala 33:19:@948.4]
  assign _GEN_164 = 5'h4 == select_5 ? io_inData_4 : _GEN_163; // @[Switch.scala 33:19:@948.4]
  assign _GEN_165 = 5'h5 == select_5 ? io_inData_5 : _GEN_164; // @[Switch.scala 33:19:@948.4]
  assign _GEN_166 = 5'h6 == select_5 ? io_inData_6 : _GEN_165; // @[Switch.scala 33:19:@948.4]
  assign _GEN_167 = 5'h7 == select_5 ? io_inData_7 : _GEN_166; // @[Switch.scala 33:19:@948.4]
  assign _GEN_168 = 5'h8 == select_5 ? io_inData_8 : _GEN_167; // @[Switch.scala 33:19:@948.4]
  assign _GEN_169 = 5'h9 == select_5 ? io_inData_9 : _GEN_168; // @[Switch.scala 33:19:@948.4]
  assign _GEN_170 = 5'ha == select_5 ? io_inData_10 : _GEN_169; // @[Switch.scala 33:19:@948.4]
  assign _GEN_171 = 5'hb == select_5 ? io_inData_11 : _GEN_170; // @[Switch.scala 33:19:@948.4]
  assign _GEN_172 = 5'hc == select_5 ? io_inData_12 : _GEN_171; // @[Switch.scala 33:19:@948.4]
  assign _GEN_173 = 5'hd == select_5 ? io_inData_13 : _GEN_172; // @[Switch.scala 33:19:@948.4]
  assign _GEN_174 = 5'he == select_5 ? io_inData_14 : _GEN_173; // @[Switch.scala 33:19:@948.4]
  assign _GEN_175 = 5'hf == select_5 ? io_inData_15 : _GEN_174; // @[Switch.scala 33:19:@948.4]
  assign _GEN_176 = 5'h10 == select_5 ? io_inData_16 : _GEN_175; // @[Switch.scala 33:19:@948.4]
  assign _GEN_177 = 5'h11 == select_5 ? io_inData_17 : _GEN_176; // @[Switch.scala 33:19:@948.4]
  assign _GEN_178 = 5'h12 == select_5 ? io_inData_18 : _GEN_177; // @[Switch.scala 33:19:@948.4]
  assign _GEN_179 = 5'h13 == select_5 ? io_inData_19 : _GEN_178; // @[Switch.scala 33:19:@948.4]
  assign _GEN_180 = 5'h14 == select_5 ? io_inData_20 : _GEN_179; // @[Switch.scala 33:19:@948.4]
  assign _GEN_181 = 5'h15 == select_5 ? io_inData_21 : _GEN_180; // @[Switch.scala 33:19:@948.4]
  assign _GEN_182 = 5'h16 == select_5 ? io_inData_22 : _GEN_181; // @[Switch.scala 33:19:@948.4]
  assign _GEN_183 = 5'h17 == select_5 ? io_inData_23 : _GEN_182; // @[Switch.scala 33:19:@948.4]
  assign _GEN_184 = 5'h18 == select_5 ? io_inData_24 : _GEN_183; // @[Switch.scala 33:19:@948.4]
  assign _GEN_185 = 5'h19 == select_5 ? io_inData_25 : _GEN_184; // @[Switch.scala 33:19:@948.4]
  assign _GEN_186 = 5'h1a == select_5 ? io_inData_26 : _GEN_185; // @[Switch.scala 33:19:@948.4]
  assign _GEN_187 = 5'h1b == select_5 ? io_inData_27 : _GEN_186; // @[Switch.scala 33:19:@948.4]
  assign _GEN_188 = 5'h1c == select_5 ? io_inData_28 : _GEN_187; // @[Switch.scala 33:19:@948.4]
  assign _GEN_189 = 5'h1d == select_5 ? io_inData_29 : _GEN_188; // @[Switch.scala 33:19:@948.4]
  assign _GEN_190 = 5'h1e == select_5 ? io_inData_30 : _GEN_189; // @[Switch.scala 33:19:@948.4]
  assign _T_5888 = {valid_5_7,valid_5_6,valid_5_5,valid_5_4,valid_5_3,valid_5_2,valid_5_1,valid_5_0}; // @[Switch.scala 34:32:@955.4]
  assign _T_5896 = {valid_5_15,valid_5_14,valid_5_13,valid_5_12,valid_5_11,valid_5_10,valid_5_9,valid_5_8,_T_5888}; // @[Switch.scala 34:32:@963.4]
  assign _T_5903 = {valid_5_23,valid_5_22,valid_5_21,valid_5_20,valid_5_19,valid_5_18,valid_5_17,valid_5_16}; // @[Switch.scala 34:32:@970.4]
  assign _T_5912 = {valid_5_31,valid_5_30,valid_5_29,valid_5_28,valid_5_27,valid_5_26,valid_5_25,valid_5_24,_T_5903,_T_5896}; // @[Switch.scala 34:32:@979.4]
  assign _T_5916 = io_inAddr_0 == 5'h6; // @[Switch.scala 30:53:@982.4]
  assign valid_6_0 = io_inValid_0 & _T_5916; // @[Switch.scala 30:36:@983.4]
  assign _T_5919 = io_inAddr_1 == 5'h6; // @[Switch.scala 30:53:@985.4]
  assign valid_6_1 = io_inValid_1 & _T_5919; // @[Switch.scala 30:36:@986.4]
  assign _T_5922 = io_inAddr_2 == 5'h6; // @[Switch.scala 30:53:@988.4]
  assign valid_6_2 = io_inValid_2 & _T_5922; // @[Switch.scala 30:36:@989.4]
  assign _T_5925 = io_inAddr_3 == 5'h6; // @[Switch.scala 30:53:@991.4]
  assign valid_6_3 = io_inValid_3 & _T_5925; // @[Switch.scala 30:36:@992.4]
  assign _T_5928 = io_inAddr_4 == 5'h6; // @[Switch.scala 30:53:@994.4]
  assign valid_6_4 = io_inValid_4 & _T_5928; // @[Switch.scala 30:36:@995.4]
  assign _T_5931 = io_inAddr_5 == 5'h6; // @[Switch.scala 30:53:@997.4]
  assign valid_6_5 = io_inValid_5 & _T_5931; // @[Switch.scala 30:36:@998.4]
  assign _T_5934 = io_inAddr_6 == 5'h6; // @[Switch.scala 30:53:@1000.4]
  assign valid_6_6 = io_inValid_6 & _T_5934; // @[Switch.scala 30:36:@1001.4]
  assign _T_5937 = io_inAddr_7 == 5'h6; // @[Switch.scala 30:53:@1003.4]
  assign valid_6_7 = io_inValid_7 & _T_5937; // @[Switch.scala 30:36:@1004.4]
  assign _T_5940 = io_inAddr_8 == 5'h6; // @[Switch.scala 30:53:@1006.4]
  assign valid_6_8 = io_inValid_8 & _T_5940; // @[Switch.scala 30:36:@1007.4]
  assign _T_5943 = io_inAddr_9 == 5'h6; // @[Switch.scala 30:53:@1009.4]
  assign valid_6_9 = io_inValid_9 & _T_5943; // @[Switch.scala 30:36:@1010.4]
  assign _T_5946 = io_inAddr_10 == 5'h6; // @[Switch.scala 30:53:@1012.4]
  assign valid_6_10 = io_inValid_10 & _T_5946; // @[Switch.scala 30:36:@1013.4]
  assign _T_5949 = io_inAddr_11 == 5'h6; // @[Switch.scala 30:53:@1015.4]
  assign valid_6_11 = io_inValid_11 & _T_5949; // @[Switch.scala 30:36:@1016.4]
  assign _T_5952 = io_inAddr_12 == 5'h6; // @[Switch.scala 30:53:@1018.4]
  assign valid_6_12 = io_inValid_12 & _T_5952; // @[Switch.scala 30:36:@1019.4]
  assign _T_5955 = io_inAddr_13 == 5'h6; // @[Switch.scala 30:53:@1021.4]
  assign valid_6_13 = io_inValid_13 & _T_5955; // @[Switch.scala 30:36:@1022.4]
  assign _T_5958 = io_inAddr_14 == 5'h6; // @[Switch.scala 30:53:@1024.4]
  assign valid_6_14 = io_inValid_14 & _T_5958; // @[Switch.scala 30:36:@1025.4]
  assign _T_5961 = io_inAddr_15 == 5'h6; // @[Switch.scala 30:53:@1027.4]
  assign valid_6_15 = io_inValid_15 & _T_5961; // @[Switch.scala 30:36:@1028.4]
  assign _T_5964 = io_inAddr_16 == 5'h6; // @[Switch.scala 30:53:@1030.4]
  assign valid_6_16 = io_inValid_16 & _T_5964; // @[Switch.scala 30:36:@1031.4]
  assign _T_5967 = io_inAddr_17 == 5'h6; // @[Switch.scala 30:53:@1033.4]
  assign valid_6_17 = io_inValid_17 & _T_5967; // @[Switch.scala 30:36:@1034.4]
  assign _T_5970 = io_inAddr_18 == 5'h6; // @[Switch.scala 30:53:@1036.4]
  assign valid_6_18 = io_inValid_18 & _T_5970; // @[Switch.scala 30:36:@1037.4]
  assign _T_5973 = io_inAddr_19 == 5'h6; // @[Switch.scala 30:53:@1039.4]
  assign valid_6_19 = io_inValid_19 & _T_5973; // @[Switch.scala 30:36:@1040.4]
  assign _T_5976 = io_inAddr_20 == 5'h6; // @[Switch.scala 30:53:@1042.4]
  assign valid_6_20 = io_inValid_20 & _T_5976; // @[Switch.scala 30:36:@1043.4]
  assign _T_5979 = io_inAddr_21 == 5'h6; // @[Switch.scala 30:53:@1045.4]
  assign valid_6_21 = io_inValid_21 & _T_5979; // @[Switch.scala 30:36:@1046.4]
  assign _T_5982 = io_inAddr_22 == 5'h6; // @[Switch.scala 30:53:@1048.4]
  assign valid_6_22 = io_inValid_22 & _T_5982; // @[Switch.scala 30:36:@1049.4]
  assign _T_5985 = io_inAddr_23 == 5'h6; // @[Switch.scala 30:53:@1051.4]
  assign valid_6_23 = io_inValid_23 & _T_5985; // @[Switch.scala 30:36:@1052.4]
  assign _T_5988 = io_inAddr_24 == 5'h6; // @[Switch.scala 30:53:@1054.4]
  assign valid_6_24 = io_inValid_24 & _T_5988; // @[Switch.scala 30:36:@1055.4]
  assign _T_5991 = io_inAddr_25 == 5'h6; // @[Switch.scala 30:53:@1057.4]
  assign valid_6_25 = io_inValid_25 & _T_5991; // @[Switch.scala 30:36:@1058.4]
  assign _T_5994 = io_inAddr_26 == 5'h6; // @[Switch.scala 30:53:@1060.4]
  assign valid_6_26 = io_inValid_26 & _T_5994; // @[Switch.scala 30:36:@1061.4]
  assign _T_5997 = io_inAddr_27 == 5'h6; // @[Switch.scala 30:53:@1063.4]
  assign valid_6_27 = io_inValid_27 & _T_5997; // @[Switch.scala 30:36:@1064.4]
  assign _T_6000 = io_inAddr_28 == 5'h6; // @[Switch.scala 30:53:@1066.4]
  assign valid_6_28 = io_inValid_28 & _T_6000; // @[Switch.scala 30:36:@1067.4]
  assign _T_6003 = io_inAddr_29 == 5'h6; // @[Switch.scala 30:53:@1069.4]
  assign valid_6_29 = io_inValid_29 & _T_6003; // @[Switch.scala 30:36:@1070.4]
  assign _T_6006 = io_inAddr_30 == 5'h6; // @[Switch.scala 30:53:@1072.4]
  assign valid_6_30 = io_inValid_30 & _T_6006; // @[Switch.scala 30:36:@1073.4]
  assign _T_6009 = io_inAddr_31 == 5'h6; // @[Switch.scala 30:53:@1075.4]
  assign valid_6_31 = io_inValid_31 & _T_6009; // @[Switch.scala 30:36:@1076.4]
  assign _T_6043 = valid_6_30 ? 5'h1e : 5'h1f; // @[Mux.scala 31:69:@1078.4]
  assign _T_6044 = valid_6_29 ? 5'h1d : _T_6043; // @[Mux.scala 31:69:@1079.4]
  assign _T_6045 = valid_6_28 ? 5'h1c : _T_6044; // @[Mux.scala 31:69:@1080.4]
  assign _T_6046 = valid_6_27 ? 5'h1b : _T_6045; // @[Mux.scala 31:69:@1081.4]
  assign _T_6047 = valid_6_26 ? 5'h1a : _T_6046; // @[Mux.scala 31:69:@1082.4]
  assign _T_6048 = valid_6_25 ? 5'h19 : _T_6047; // @[Mux.scala 31:69:@1083.4]
  assign _T_6049 = valid_6_24 ? 5'h18 : _T_6048; // @[Mux.scala 31:69:@1084.4]
  assign _T_6050 = valid_6_23 ? 5'h17 : _T_6049; // @[Mux.scala 31:69:@1085.4]
  assign _T_6051 = valid_6_22 ? 5'h16 : _T_6050; // @[Mux.scala 31:69:@1086.4]
  assign _T_6052 = valid_6_21 ? 5'h15 : _T_6051; // @[Mux.scala 31:69:@1087.4]
  assign _T_6053 = valid_6_20 ? 5'h14 : _T_6052; // @[Mux.scala 31:69:@1088.4]
  assign _T_6054 = valid_6_19 ? 5'h13 : _T_6053; // @[Mux.scala 31:69:@1089.4]
  assign _T_6055 = valid_6_18 ? 5'h12 : _T_6054; // @[Mux.scala 31:69:@1090.4]
  assign _T_6056 = valid_6_17 ? 5'h11 : _T_6055; // @[Mux.scala 31:69:@1091.4]
  assign _T_6057 = valid_6_16 ? 5'h10 : _T_6056; // @[Mux.scala 31:69:@1092.4]
  assign _T_6058 = valid_6_15 ? 5'hf : _T_6057; // @[Mux.scala 31:69:@1093.4]
  assign _T_6059 = valid_6_14 ? 5'he : _T_6058; // @[Mux.scala 31:69:@1094.4]
  assign _T_6060 = valid_6_13 ? 5'hd : _T_6059; // @[Mux.scala 31:69:@1095.4]
  assign _T_6061 = valid_6_12 ? 5'hc : _T_6060; // @[Mux.scala 31:69:@1096.4]
  assign _T_6062 = valid_6_11 ? 5'hb : _T_6061; // @[Mux.scala 31:69:@1097.4]
  assign _T_6063 = valid_6_10 ? 5'ha : _T_6062; // @[Mux.scala 31:69:@1098.4]
  assign _T_6064 = valid_6_9 ? 5'h9 : _T_6063; // @[Mux.scala 31:69:@1099.4]
  assign _T_6065 = valid_6_8 ? 5'h8 : _T_6064; // @[Mux.scala 31:69:@1100.4]
  assign _T_6066 = valid_6_7 ? 5'h7 : _T_6065; // @[Mux.scala 31:69:@1101.4]
  assign _T_6067 = valid_6_6 ? 5'h6 : _T_6066; // @[Mux.scala 31:69:@1102.4]
  assign _T_6068 = valid_6_5 ? 5'h5 : _T_6067; // @[Mux.scala 31:69:@1103.4]
  assign _T_6069 = valid_6_4 ? 5'h4 : _T_6068; // @[Mux.scala 31:69:@1104.4]
  assign _T_6070 = valid_6_3 ? 5'h3 : _T_6069; // @[Mux.scala 31:69:@1105.4]
  assign _T_6071 = valid_6_2 ? 5'h2 : _T_6070; // @[Mux.scala 31:69:@1106.4]
  assign _T_6072 = valid_6_1 ? 5'h1 : _T_6071; // @[Mux.scala 31:69:@1107.4]
  assign select_6 = valid_6_0 ? 5'h0 : _T_6072; // @[Mux.scala 31:69:@1108.4]
  assign _GEN_193 = 5'h1 == select_6 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@1110.4]
  assign _GEN_194 = 5'h2 == select_6 ? io_inData_2 : _GEN_193; // @[Switch.scala 33:19:@1110.4]
  assign _GEN_195 = 5'h3 == select_6 ? io_inData_3 : _GEN_194; // @[Switch.scala 33:19:@1110.4]
  assign _GEN_196 = 5'h4 == select_6 ? io_inData_4 : _GEN_195; // @[Switch.scala 33:19:@1110.4]
  assign _GEN_197 = 5'h5 == select_6 ? io_inData_5 : _GEN_196; // @[Switch.scala 33:19:@1110.4]
  assign _GEN_198 = 5'h6 == select_6 ? io_inData_6 : _GEN_197; // @[Switch.scala 33:19:@1110.4]
  assign _GEN_199 = 5'h7 == select_6 ? io_inData_7 : _GEN_198; // @[Switch.scala 33:19:@1110.4]
  assign _GEN_200 = 5'h8 == select_6 ? io_inData_8 : _GEN_199; // @[Switch.scala 33:19:@1110.4]
  assign _GEN_201 = 5'h9 == select_6 ? io_inData_9 : _GEN_200; // @[Switch.scala 33:19:@1110.4]
  assign _GEN_202 = 5'ha == select_6 ? io_inData_10 : _GEN_201; // @[Switch.scala 33:19:@1110.4]
  assign _GEN_203 = 5'hb == select_6 ? io_inData_11 : _GEN_202; // @[Switch.scala 33:19:@1110.4]
  assign _GEN_204 = 5'hc == select_6 ? io_inData_12 : _GEN_203; // @[Switch.scala 33:19:@1110.4]
  assign _GEN_205 = 5'hd == select_6 ? io_inData_13 : _GEN_204; // @[Switch.scala 33:19:@1110.4]
  assign _GEN_206 = 5'he == select_6 ? io_inData_14 : _GEN_205; // @[Switch.scala 33:19:@1110.4]
  assign _GEN_207 = 5'hf == select_6 ? io_inData_15 : _GEN_206; // @[Switch.scala 33:19:@1110.4]
  assign _GEN_208 = 5'h10 == select_6 ? io_inData_16 : _GEN_207; // @[Switch.scala 33:19:@1110.4]
  assign _GEN_209 = 5'h11 == select_6 ? io_inData_17 : _GEN_208; // @[Switch.scala 33:19:@1110.4]
  assign _GEN_210 = 5'h12 == select_6 ? io_inData_18 : _GEN_209; // @[Switch.scala 33:19:@1110.4]
  assign _GEN_211 = 5'h13 == select_6 ? io_inData_19 : _GEN_210; // @[Switch.scala 33:19:@1110.4]
  assign _GEN_212 = 5'h14 == select_6 ? io_inData_20 : _GEN_211; // @[Switch.scala 33:19:@1110.4]
  assign _GEN_213 = 5'h15 == select_6 ? io_inData_21 : _GEN_212; // @[Switch.scala 33:19:@1110.4]
  assign _GEN_214 = 5'h16 == select_6 ? io_inData_22 : _GEN_213; // @[Switch.scala 33:19:@1110.4]
  assign _GEN_215 = 5'h17 == select_6 ? io_inData_23 : _GEN_214; // @[Switch.scala 33:19:@1110.4]
  assign _GEN_216 = 5'h18 == select_6 ? io_inData_24 : _GEN_215; // @[Switch.scala 33:19:@1110.4]
  assign _GEN_217 = 5'h19 == select_6 ? io_inData_25 : _GEN_216; // @[Switch.scala 33:19:@1110.4]
  assign _GEN_218 = 5'h1a == select_6 ? io_inData_26 : _GEN_217; // @[Switch.scala 33:19:@1110.4]
  assign _GEN_219 = 5'h1b == select_6 ? io_inData_27 : _GEN_218; // @[Switch.scala 33:19:@1110.4]
  assign _GEN_220 = 5'h1c == select_6 ? io_inData_28 : _GEN_219; // @[Switch.scala 33:19:@1110.4]
  assign _GEN_221 = 5'h1d == select_6 ? io_inData_29 : _GEN_220; // @[Switch.scala 33:19:@1110.4]
  assign _GEN_222 = 5'h1e == select_6 ? io_inData_30 : _GEN_221; // @[Switch.scala 33:19:@1110.4]
  assign _T_6081 = {valid_6_7,valid_6_6,valid_6_5,valid_6_4,valid_6_3,valid_6_2,valid_6_1,valid_6_0}; // @[Switch.scala 34:32:@1117.4]
  assign _T_6089 = {valid_6_15,valid_6_14,valid_6_13,valid_6_12,valid_6_11,valid_6_10,valid_6_9,valid_6_8,_T_6081}; // @[Switch.scala 34:32:@1125.4]
  assign _T_6096 = {valid_6_23,valid_6_22,valid_6_21,valid_6_20,valid_6_19,valid_6_18,valid_6_17,valid_6_16}; // @[Switch.scala 34:32:@1132.4]
  assign _T_6105 = {valid_6_31,valid_6_30,valid_6_29,valid_6_28,valid_6_27,valid_6_26,valid_6_25,valid_6_24,_T_6096,_T_6089}; // @[Switch.scala 34:32:@1141.4]
  assign _T_6109 = io_inAddr_0 == 5'h7; // @[Switch.scala 30:53:@1144.4]
  assign valid_7_0 = io_inValid_0 & _T_6109; // @[Switch.scala 30:36:@1145.4]
  assign _T_6112 = io_inAddr_1 == 5'h7; // @[Switch.scala 30:53:@1147.4]
  assign valid_7_1 = io_inValid_1 & _T_6112; // @[Switch.scala 30:36:@1148.4]
  assign _T_6115 = io_inAddr_2 == 5'h7; // @[Switch.scala 30:53:@1150.4]
  assign valid_7_2 = io_inValid_2 & _T_6115; // @[Switch.scala 30:36:@1151.4]
  assign _T_6118 = io_inAddr_3 == 5'h7; // @[Switch.scala 30:53:@1153.4]
  assign valid_7_3 = io_inValid_3 & _T_6118; // @[Switch.scala 30:36:@1154.4]
  assign _T_6121 = io_inAddr_4 == 5'h7; // @[Switch.scala 30:53:@1156.4]
  assign valid_7_4 = io_inValid_4 & _T_6121; // @[Switch.scala 30:36:@1157.4]
  assign _T_6124 = io_inAddr_5 == 5'h7; // @[Switch.scala 30:53:@1159.4]
  assign valid_7_5 = io_inValid_5 & _T_6124; // @[Switch.scala 30:36:@1160.4]
  assign _T_6127 = io_inAddr_6 == 5'h7; // @[Switch.scala 30:53:@1162.4]
  assign valid_7_6 = io_inValid_6 & _T_6127; // @[Switch.scala 30:36:@1163.4]
  assign _T_6130 = io_inAddr_7 == 5'h7; // @[Switch.scala 30:53:@1165.4]
  assign valid_7_7 = io_inValid_7 & _T_6130; // @[Switch.scala 30:36:@1166.4]
  assign _T_6133 = io_inAddr_8 == 5'h7; // @[Switch.scala 30:53:@1168.4]
  assign valid_7_8 = io_inValid_8 & _T_6133; // @[Switch.scala 30:36:@1169.4]
  assign _T_6136 = io_inAddr_9 == 5'h7; // @[Switch.scala 30:53:@1171.4]
  assign valid_7_9 = io_inValid_9 & _T_6136; // @[Switch.scala 30:36:@1172.4]
  assign _T_6139 = io_inAddr_10 == 5'h7; // @[Switch.scala 30:53:@1174.4]
  assign valid_7_10 = io_inValid_10 & _T_6139; // @[Switch.scala 30:36:@1175.4]
  assign _T_6142 = io_inAddr_11 == 5'h7; // @[Switch.scala 30:53:@1177.4]
  assign valid_7_11 = io_inValid_11 & _T_6142; // @[Switch.scala 30:36:@1178.4]
  assign _T_6145 = io_inAddr_12 == 5'h7; // @[Switch.scala 30:53:@1180.4]
  assign valid_7_12 = io_inValid_12 & _T_6145; // @[Switch.scala 30:36:@1181.4]
  assign _T_6148 = io_inAddr_13 == 5'h7; // @[Switch.scala 30:53:@1183.4]
  assign valid_7_13 = io_inValid_13 & _T_6148; // @[Switch.scala 30:36:@1184.4]
  assign _T_6151 = io_inAddr_14 == 5'h7; // @[Switch.scala 30:53:@1186.4]
  assign valid_7_14 = io_inValid_14 & _T_6151; // @[Switch.scala 30:36:@1187.4]
  assign _T_6154 = io_inAddr_15 == 5'h7; // @[Switch.scala 30:53:@1189.4]
  assign valid_7_15 = io_inValid_15 & _T_6154; // @[Switch.scala 30:36:@1190.4]
  assign _T_6157 = io_inAddr_16 == 5'h7; // @[Switch.scala 30:53:@1192.4]
  assign valid_7_16 = io_inValid_16 & _T_6157; // @[Switch.scala 30:36:@1193.4]
  assign _T_6160 = io_inAddr_17 == 5'h7; // @[Switch.scala 30:53:@1195.4]
  assign valid_7_17 = io_inValid_17 & _T_6160; // @[Switch.scala 30:36:@1196.4]
  assign _T_6163 = io_inAddr_18 == 5'h7; // @[Switch.scala 30:53:@1198.4]
  assign valid_7_18 = io_inValid_18 & _T_6163; // @[Switch.scala 30:36:@1199.4]
  assign _T_6166 = io_inAddr_19 == 5'h7; // @[Switch.scala 30:53:@1201.4]
  assign valid_7_19 = io_inValid_19 & _T_6166; // @[Switch.scala 30:36:@1202.4]
  assign _T_6169 = io_inAddr_20 == 5'h7; // @[Switch.scala 30:53:@1204.4]
  assign valid_7_20 = io_inValid_20 & _T_6169; // @[Switch.scala 30:36:@1205.4]
  assign _T_6172 = io_inAddr_21 == 5'h7; // @[Switch.scala 30:53:@1207.4]
  assign valid_7_21 = io_inValid_21 & _T_6172; // @[Switch.scala 30:36:@1208.4]
  assign _T_6175 = io_inAddr_22 == 5'h7; // @[Switch.scala 30:53:@1210.4]
  assign valid_7_22 = io_inValid_22 & _T_6175; // @[Switch.scala 30:36:@1211.4]
  assign _T_6178 = io_inAddr_23 == 5'h7; // @[Switch.scala 30:53:@1213.4]
  assign valid_7_23 = io_inValid_23 & _T_6178; // @[Switch.scala 30:36:@1214.4]
  assign _T_6181 = io_inAddr_24 == 5'h7; // @[Switch.scala 30:53:@1216.4]
  assign valid_7_24 = io_inValid_24 & _T_6181; // @[Switch.scala 30:36:@1217.4]
  assign _T_6184 = io_inAddr_25 == 5'h7; // @[Switch.scala 30:53:@1219.4]
  assign valid_7_25 = io_inValid_25 & _T_6184; // @[Switch.scala 30:36:@1220.4]
  assign _T_6187 = io_inAddr_26 == 5'h7; // @[Switch.scala 30:53:@1222.4]
  assign valid_7_26 = io_inValid_26 & _T_6187; // @[Switch.scala 30:36:@1223.4]
  assign _T_6190 = io_inAddr_27 == 5'h7; // @[Switch.scala 30:53:@1225.4]
  assign valid_7_27 = io_inValid_27 & _T_6190; // @[Switch.scala 30:36:@1226.4]
  assign _T_6193 = io_inAddr_28 == 5'h7; // @[Switch.scala 30:53:@1228.4]
  assign valid_7_28 = io_inValid_28 & _T_6193; // @[Switch.scala 30:36:@1229.4]
  assign _T_6196 = io_inAddr_29 == 5'h7; // @[Switch.scala 30:53:@1231.4]
  assign valid_7_29 = io_inValid_29 & _T_6196; // @[Switch.scala 30:36:@1232.4]
  assign _T_6199 = io_inAddr_30 == 5'h7; // @[Switch.scala 30:53:@1234.4]
  assign valid_7_30 = io_inValid_30 & _T_6199; // @[Switch.scala 30:36:@1235.4]
  assign _T_6202 = io_inAddr_31 == 5'h7; // @[Switch.scala 30:53:@1237.4]
  assign valid_7_31 = io_inValid_31 & _T_6202; // @[Switch.scala 30:36:@1238.4]
  assign _T_6236 = valid_7_30 ? 5'h1e : 5'h1f; // @[Mux.scala 31:69:@1240.4]
  assign _T_6237 = valid_7_29 ? 5'h1d : _T_6236; // @[Mux.scala 31:69:@1241.4]
  assign _T_6238 = valid_7_28 ? 5'h1c : _T_6237; // @[Mux.scala 31:69:@1242.4]
  assign _T_6239 = valid_7_27 ? 5'h1b : _T_6238; // @[Mux.scala 31:69:@1243.4]
  assign _T_6240 = valid_7_26 ? 5'h1a : _T_6239; // @[Mux.scala 31:69:@1244.4]
  assign _T_6241 = valid_7_25 ? 5'h19 : _T_6240; // @[Mux.scala 31:69:@1245.4]
  assign _T_6242 = valid_7_24 ? 5'h18 : _T_6241; // @[Mux.scala 31:69:@1246.4]
  assign _T_6243 = valid_7_23 ? 5'h17 : _T_6242; // @[Mux.scala 31:69:@1247.4]
  assign _T_6244 = valid_7_22 ? 5'h16 : _T_6243; // @[Mux.scala 31:69:@1248.4]
  assign _T_6245 = valid_7_21 ? 5'h15 : _T_6244; // @[Mux.scala 31:69:@1249.4]
  assign _T_6246 = valid_7_20 ? 5'h14 : _T_6245; // @[Mux.scala 31:69:@1250.4]
  assign _T_6247 = valid_7_19 ? 5'h13 : _T_6246; // @[Mux.scala 31:69:@1251.4]
  assign _T_6248 = valid_7_18 ? 5'h12 : _T_6247; // @[Mux.scala 31:69:@1252.4]
  assign _T_6249 = valid_7_17 ? 5'h11 : _T_6248; // @[Mux.scala 31:69:@1253.4]
  assign _T_6250 = valid_7_16 ? 5'h10 : _T_6249; // @[Mux.scala 31:69:@1254.4]
  assign _T_6251 = valid_7_15 ? 5'hf : _T_6250; // @[Mux.scala 31:69:@1255.4]
  assign _T_6252 = valid_7_14 ? 5'he : _T_6251; // @[Mux.scala 31:69:@1256.4]
  assign _T_6253 = valid_7_13 ? 5'hd : _T_6252; // @[Mux.scala 31:69:@1257.4]
  assign _T_6254 = valid_7_12 ? 5'hc : _T_6253; // @[Mux.scala 31:69:@1258.4]
  assign _T_6255 = valid_7_11 ? 5'hb : _T_6254; // @[Mux.scala 31:69:@1259.4]
  assign _T_6256 = valid_7_10 ? 5'ha : _T_6255; // @[Mux.scala 31:69:@1260.4]
  assign _T_6257 = valid_7_9 ? 5'h9 : _T_6256; // @[Mux.scala 31:69:@1261.4]
  assign _T_6258 = valid_7_8 ? 5'h8 : _T_6257; // @[Mux.scala 31:69:@1262.4]
  assign _T_6259 = valid_7_7 ? 5'h7 : _T_6258; // @[Mux.scala 31:69:@1263.4]
  assign _T_6260 = valid_7_6 ? 5'h6 : _T_6259; // @[Mux.scala 31:69:@1264.4]
  assign _T_6261 = valid_7_5 ? 5'h5 : _T_6260; // @[Mux.scala 31:69:@1265.4]
  assign _T_6262 = valid_7_4 ? 5'h4 : _T_6261; // @[Mux.scala 31:69:@1266.4]
  assign _T_6263 = valid_7_3 ? 5'h3 : _T_6262; // @[Mux.scala 31:69:@1267.4]
  assign _T_6264 = valid_7_2 ? 5'h2 : _T_6263; // @[Mux.scala 31:69:@1268.4]
  assign _T_6265 = valid_7_1 ? 5'h1 : _T_6264; // @[Mux.scala 31:69:@1269.4]
  assign select_7 = valid_7_0 ? 5'h0 : _T_6265; // @[Mux.scala 31:69:@1270.4]
  assign _GEN_225 = 5'h1 == select_7 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@1272.4]
  assign _GEN_226 = 5'h2 == select_7 ? io_inData_2 : _GEN_225; // @[Switch.scala 33:19:@1272.4]
  assign _GEN_227 = 5'h3 == select_7 ? io_inData_3 : _GEN_226; // @[Switch.scala 33:19:@1272.4]
  assign _GEN_228 = 5'h4 == select_7 ? io_inData_4 : _GEN_227; // @[Switch.scala 33:19:@1272.4]
  assign _GEN_229 = 5'h5 == select_7 ? io_inData_5 : _GEN_228; // @[Switch.scala 33:19:@1272.4]
  assign _GEN_230 = 5'h6 == select_7 ? io_inData_6 : _GEN_229; // @[Switch.scala 33:19:@1272.4]
  assign _GEN_231 = 5'h7 == select_7 ? io_inData_7 : _GEN_230; // @[Switch.scala 33:19:@1272.4]
  assign _GEN_232 = 5'h8 == select_7 ? io_inData_8 : _GEN_231; // @[Switch.scala 33:19:@1272.4]
  assign _GEN_233 = 5'h9 == select_7 ? io_inData_9 : _GEN_232; // @[Switch.scala 33:19:@1272.4]
  assign _GEN_234 = 5'ha == select_7 ? io_inData_10 : _GEN_233; // @[Switch.scala 33:19:@1272.4]
  assign _GEN_235 = 5'hb == select_7 ? io_inData_11 : _GEN_234; // @[Switch.scala 33:19:@1272.4]
  assign _GEN_236 = 5'hc == select_7 ? io_inData_12 : _GEN_235; // @[Switch.scala 33:19:@1272.4]
  assign _GEN_237 = 5'hd == select_7 ? io_inData_13 : _GEN_236; // @[Switch.scala 33:19:@1272.4]
  assign _GEN_238 = 5'he == select_7 ? io_inData_14 : _GEN_237; // @[Switch.scala 33:19:@1272.4]
  assign _GEN_239 = 5'hf == select_7 ? io_inData_15 : _GEN_238; // @[Switch.scala 33:19:@1272.4]
  assign _GEN_240 = 5'h10 == select_7 ? io_inData_16 : _GEN_239; // @[Switch.scala 33:19:@1272.4]
  assign _GEN_241 = 5'h11 == select_7 ? io_inData_17 : _GEN_240; // @[Switch.scala 33:19:@1272.4]
  assign _GEN_242 = 5'h12 == select_7 ? io_inData_18 : _GEN_241; // @[Switch.scala 33:19:@1272.4]
  assign _GEN_243 = 5'h13 == select_7 ? io_inData_19 : _GEN_242; // @[Switch.scala 33:19:@1272.4]
  assign _GEN_244 = 5'h14 == select_7 ? io_inData_20 : _GEN_243; // @[Switch.scala 33:19:@1272.4]
  assign _GEN_245 = 5'h15 == select_7 ? io_inData_21 : _GEN_244; // @[Switch.scala 33:19:@1272.4]
  assign _GEN_246 = 5'h16 == select_7 ? io_inData_22 : _GEN_245; // @[Switch.scala 33:19:@1272.4]
  assign _GEN_247 = 5'h17 == select_7 ? io_inData_23 : _GEN_246; // @[Switch.scala 33:19:@1272.4]
  assign _GEN_248 = 5'h18 == select_7 ? io_inData_24 : _GEN_247; // @[Switch.scala 33:19:@1272.4]
  assign _GEN_249 = 5'h19 == select_7 ? io_inData_25 : _GEN_248; // @[Switch.scala 33:19:@1272.4]
  assign _GEN_250 = 5'h1a == select_7 ? io_inData_26 : _GEN_249; // @[Switch.scala 33:19:@1272.4]
  assign _GEN_251 = 5'h1b == select_7 ? io_inData_27 : _GEN_250; // @[Switch.scala 33:19:@1272.4]
  assign _GEN_252 = 5'h1c == select_7 ? io_inData_28 : _GEN_251; // @[Switch.scala 33:19:@1272.4]
  assign _GEN_253 = 5'h1d == select_7 ? io_inData_29 : _GEN_252; // @[Switch.scala 33:19:@1272.4]
  assign _GEN_254 = 5'h1e == select_7 ? io_inData_30 : _GEN_253; // @[Switch.scala 33:19:@1272.4]
  assign _T_6274 = {valid_7_7,valid_7_6,valid_7_5,valid_7_4,valid_7_3,valid_7_2,valid_7_1,valid_7_0}; // @[Switch.scala 34:32:@1279.4]
  assign _T_6282 = {valid_7_15,valid_7_14,valid_7_13,valid_7_12,valid_7_11,valid_7_10,valid_7_9,valid_7_8,_T_6274}; // @[Switch.scala 34:32:@1287.4]
  assign _T_6289 = {valid_7_23,valid_7_22,valid_7_21,valid_7_20,valid_7_19,valid_7_18,valid_7_17,valid_7_16}; // @[Switch.scala 34:32:@1294.4]
  assign _T_6298 = {valid_7_31,valid_7_30,valid_7_29,valid_7_28,valid_7_27,valid_7_26,valid_7_25,valid_7_24,_T_6289,_T_6282}; // @[Switch.scala 34:32:@1303.4]
  assign _T_6302 = io_inAddr_0 == 5'h8; // @[Switch.scala 30:53:@1306.4]
  assign valid_8_0 = io_inValid_0 & _T_6302; // @[Switch.scala 30:36:@1307.4]
  assign _T_6305 = io_inAddr_1 == 5'h8; // @[Switch.scala 30:53:@1309.4]
  assign valid_8_1 = io_inValid_1 & _T_6305; // @[Switch.scala 30:36:@1310.4]
  assign _T_6308 = io_inAddr_2 == 5'h8; // @[Switch.scala 30:53:@1312.4]
  assign valid_8_2 = io_inValid_2 & _T_6308; // @[Switch.scala 30:36:@1313.4]
  assign _T_6311 = io_inAddr_3 == 5'h8; // @[Switch.scala 30:53:@1315.4]
  assign valid_8_3 = io_inValid_3 & _T_6311; // @[Switch.scala 30:36:@1316.4]
  assign _T_6314 = io_inAddr_4 == 5'h8; // @[Switch.scala 30:53:@1318.4]
  assign valid_8_4 = io_inValid_4 & _T_6314; // @[Switch.scala 30:36:@1319.4]
  assign _T_6317 = io_inAddr_5 == 5'h8; // @[Switch.scala 30:53:@1321.4]
  assign valid_8_5 = io_inValid_5 & _T_6317; // @[Switch.scala 30:36:@1322.4]
  assign _T_6320 = io_inAddr_6 == 5'h8; // @[Switch.scala 30:53:@1324.4]
  assign valid_8_6 = io_inValid_6 & _T_6320; // @[Switch.scala 30:36:@1325.4]
  assign _T_6323 = io_inAddr_7 == 5'h8; // @[Switch.scala 30:53:@1327.4]
  assign valid_8_7 = io_inValid_7 & _T_6323; // @[Switch.scala 30:36:@1328.4]
  assign _T_6326 = io_inAddr_8 == 5'h8; // @[Switch.scala 30:53:@1330.4]
  assign valid_8_8 = io_inValid_8 & _T_6326; // @[Switch.scala 30:36:@1331.4]
  assign _T_6329 = io_inAddr_9 == 5'h8; // @[Switch.scala 30:53:@1333.4]
  assign valid_8_9 = io_inValid_9 & _T_6329; // @[Switch.scala 30:36:@1334.4]
  assign _T_6332 = io_inAddr_10 == 5'h8; // @[Switch.scala 30:53:@1336.4]
  assign valid_8_10 = io_inValid_10 & _T_6332; // @[Switch.scala 30:36:@1337.4]
  assign _T_6335 = io_inAddr_11 == 5'h8; // @[Switch.scala 30:53:@1339.4]
  assign valid_8_11 = io_inValid_11 & _T_6335; // @[Switch.scala 30:36:@1340.4]
  assign _T_6338 = io_inAddr_12 == 5'h8; // @[Switch.scala 30:53:@1342.4]
  assign valid_8_12 = io_inValid_12 & _T_6338; // @[Switch.scala 30:36:@1343.4]
  assign _T_6341 = io_inAddr_13 == 5'h8; // @[Switch.scala 30:53:@1345.4]
  assign valid_8_13 = io_inValid_13 & _T_6341; // @[Switch.scala 30:36:@1346.4]
  assign _T_6344 = io_inAddr_14 == 5'h8; // @[Switch.scala 30:53:@1348.4]
  assign valid_8_14 = io_inValid_14 & _T_6344; // @[Switch.scala 30:36:@1349.4]
  assign _T_6347 = io_inAddr_15 == 5'h8; // @[Switch.scala 30:53:@1351.4]
  assign valid_8_15 = io_inValid_15 & _T_6347; // @[Switch.scala 30:36:@1352.4]
  assign _T_6350 = io_inAddr_16 == 5'h8; // @[Switch.scala 30:53:@1354.4]
  assign valid_8_16 = io_inValid_16 & _T_6350; // @[Switch.scala 30:36:@1355.4]
  assign _T_6353 = io_inAddr_17 == 5'h8; // @[Switch.scala 30:53:@1357.4]
  assign valid_8_17 = io_inValid_17 & _T_6353; // @[Switch.scala 30:36:@1358.4]
  assign _T_6356 = io_inAddr_18 == 5'h8; // @[Switch.scala 30:53:@1360.4]
  assign valid_8_18 = io_inValid_18 & _T_6356; // @[Switch.scala 30:36:@1361.4]
  assign _T_6359 = io_inAddr_19 == 5'h8; // @[Switch.scala 30:53:@1363.4]
  assign valid_8_19 = io_inValid_19 & _T_6359; // @[Switch.scala 30:36:@1364.4]
  assign _T_6362 = io_inAddr_20 == 5'h8; // @[Switch.scala 30:53:@1366.4]
  assign valid_8_20 = io_inValid_20 & _T_6362; // @[Switch.scala 30:36:@1367.4]
  assign _T_6365 = io_inAddr_21 == 5'h8; // @[Switch.scala 30:53:@1369.4]
  assign valid_8_21 = io_inValid_21 & _T_6365; // @[Switch.scala 30:36:@1370.4]
  assign _T_6368 = io_inAddr_22 == 5'h8; // @[Switch.scala 30:53:@1372.4]
  assign valid_8_22 = io_inValid_22 & _T_6368; // @[Switch.scala 30:36:@1373.4]
  assign _T_6371 = io_inAddr_23 == 5'h8; // @[Switch.scala 30:53:@1375.4]
  assign valid_8_23 = io_inValid_23 & _T_6371; // @[Switch.scala 30:36:@1376.4]
  assign _T_6374 = io_inAddr_24 == 5'h8; // @[Switch.scala 30:53:@1378.4]
  assign valid_8_24 = io_inValid_24 & _T_6374; // @[Switch.scala 30:36:@1379.4]
  assign _T_6377 = io_inAddr_25 == 5'h8; // @[Switch.scala 30:53:@1381.4]
  assign valid_8_25 = io_inValid_25 & _T_6377; // @[Switch.scala 30:36:@1382.4]
  assign _T_6380 = io_inAddr_26 == 5'h8; // @[Switch.scala 30:53:@1384.4]
  assign valid_8_26 = io_inValid_26 & _T_6380; // @[Switch.scala 30:36:@1385.4]
  assign _T_6383 = io_inAddr_27 == 5'h8; // @[Switch.scala 30:53:@1387.4]
  assign valid_8_27 = io_inValid_27 & _T_6383; // @[Switch.scala 30:36:@1388.4]
  assign _T_6386 = io_inAddr_28 == 5'h8; // @[Switch.scala 30:53:@1390.4]
  assign valid_8_28 = io_inValid_28 & _T_6386; // @[Switch.scala 30:36:@1391.4]
  assign _T_6389 = io_inAddr_29 == 5'h8; // @[Switch.scala 30:53:@1393.4]
  assign valid_8_29 = io_inValid_29 & _T_6389; // @[Switch.scala 30:36:@1394.4]
  assign _T_6392 = io_inAddr_30 == 5'h8; // @[Switch.scala 30:53:@1396.4]
  assign valid_8_30 = io_inValid_30 & _T_6392; // @[Switch.scala 30:36:@1397.4]
  assign _T_6395 = io_inAddr_31 == 5'h8; // @[Switch.scala 30:53:@1399.4]
  assign valid_8_31 = io_inValid_31 & _T_6395; // @[Switch.scala 30:36:@1400.4]
  assign _T_6429 = valid_8_30 ? 5'h1e : 5'h1f; // @[Mux.scala 31:69:@1402.4]
  assign _T_6430 = valid_8_29 ? 5'h1d : _T_6429; // @[Mux.scala 31:69:@1403.4]
  assign _T_6431 = valid_8_28 ? 5'h1c : _T_6430; // @[Mux.scala 31:69:@1404.4]
  assign _T_6432 = valid_8_27 ? 5'h1b : _T_6431; // @[Mux.scala 31:69:@1405.4]
  assign _T_6433 = valid_8_26 ? 5'h1a : _T_6432; // @[Mux.scala 31:69:@1406.4]
  assign _T_6434 = valid_8_25 ? 5'h19 : _T_6433; // @[Mux.scala 31:69:@1407.4]
  assign _T_6435 = valid_8_24 ? 5'h18 : _T_6434; // @[Mux.scala 31:69:@1408.4]
  assign _T_6436 = valid_8_23 ? 5'h17 : _T_6435; // @[Mux.scala 31:69:@1409.4]
  assign _T_6437 = valid_8_22 ? 5'h16 : _T_6436; // @[Mux.scala 31:69:@1410.4]
  assign _T_6438 = valid_8_21 ? 5'h15 : _T_6437; // @[Mux.scala 31:69:@1411.4]
  assign _T_6439 = valid_8_20 ? 5'h14 : _T_6438; // @[Mux.scala 31:69:@1412.4]
  assign _T_6440 = valid_8_19 ? 5'h13 : _T_6439; // @[Mux.scala 31:69:@1413.4]
  assign _T_6441 = valid_8_18 ? 5'h12 : _T_6440; // @[Mux.scala 31:69:@1414.4]
  assign _T_6442 = valid_8_17 ? 5'h11 : _T_6441; // @[Mux.scala 31:69:@1415.4]
  assign _T_6443 = valid_8_16 ? 5'h10 : _T_6442; // @[Mux.scala 31:69:@1416.4]
  assign _T_6444 = valid_8_15 ? 5'hf : _T_6443; // @[Mux.scala 31:69:@1417.4]
  assign _T_6445 = valid_8_14 ? 5'he : _T_6444; // @[Mux.scala 31:69:@1418.4]
  assign _T_6446 = valid_8_13 ? 5'hd : _T_6445; // @[Mux.scala 31:69:@1419.4]
  assign _T_6447 = valid_8_12 ? 5'hc : _T_6446; // @[Mux.scala 31:69:@1420.4]
  assign _T_6448 = valid_8_11 ? 5'hb : _T_6447; // @[Mux.scala 31:69:@1421.4]
  assign _T_6449 = valid_8_10 ? 5'ha : _T_6448; // @[Mux.scala 31:69:@1422.4]
  assign _T_6450 = valid_8_9 ? 5'h9 : _T_6449; // @[Mux.scala 31:69:@1423.4]
  assign _T_6451 = valid_8_8 ? 5'h8 : _T_6450; // @[Mux.scala 31:69:@1424.4]
  assign _T_6452 = valid_8_7 ? 5'h7 : _T_6451; // @[Mux.scala 31:69:@1425.4]
  assign _T_6453 = valid_8_6 ? 5'h6 : _T_6452; // @[Mux.scala 31:69:@1426.4]
  assign _T_6454 = valid_8_5 ? 5'h5 : _T_6453; // @[Mux.scala 31:69:@1427.4]
  assign _T_6455 = valid_8_4 ? 5'h4 : _T_6454; // @[Mux.scala 31:69:@1428.4]
  assign _T_6456 = valid_8_3 ? 5'h3 : _T_6455; // @[Mux.scala 31:69:@1429.4]
  assign _T_6457 = valid_8_2 ? 5'h2 : _T_6456; // @[Mux.scala 31:69:@1430.4]
  assign _T_6458 = valid_8_1 ? 5'h1 : _T_6457; // @[Mux.scala 31:69:@1431.4]
  assign select_8 = valid_8_0 ? 5'h0 : _T_6458; // @[Mux.scala 31:69:@1432.4]
  assign _GEN_257 = 5'h1 == select_8 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@1434.4]
  assign _GEN_258 = 5'h2 == select_8 ? io_inData_2 : _GEN_257; // @[Switch.scala 33:19:@1434.4]
  assign _GEN_259 = 5'h3 == select_8 ? io_inData_3 : _GEN_258; // @[Switch.scala 33:19:@1434.4]
  assign _GEN_260 = 5'h4 == select_8 ? io_inData_4 : _GEN_259; // @[Switch.scala 33:19:@1434.4]
  assign _GEN_261 = 5'h5 == select_8 ? io_inData_5 : _GEN_260; // @[Switch.scala 33:19:@1434.4]
  assign _GEN_262 = 5'h6 == select_8 ? io_inData_6 : _GEN_261; // @[Switch.scala 33:19:@1434.4]
  assign _GEN_263 = 5'h7 == select_8 ? io_inData_7 : _GEN_262; // @[Switch.scala 33:19:@1434.4]
  assign _GEN_264 = 5'h8 == select_8 ? io_inData_8 : _GEN_263; // @[Switch.scala 33:19:@1434.4]
  assign _GEN_265 = 5'h9 == select_8 ? io_inData_9 : _GEN_264; // @[Switch.scala 33:19:@1434.4]
  assign _GEN_266 = 5'ha == select_8 ? io_inData_10 : _GEN_265; // @[Switch.scala 33:19:@1434.4]
  assign _GEN_267 = 5'hb == select_8 ? io_inData_11 : _GEN_266; // @[Switch.scala 33:19:@1434.4]
  assign _GEN_268 = 5'hc == select_8 ? io_inData_12 : _GEN_267; // @[Switch.scala 33:19:@1434.4]
  assign _GEN_269 = 5'hd == select_8 ? io_inData_13 : _GEN_268; // @[Switch.scala 33:19:@1434.4]
  assign _GEN_270 = 5'he == select_8 ? io_inData_14 : _GEN_269; // @[Switch.scala 33:19:@1434.4]
  assign _GEN_271 = 5'hf == select_8 ? io_inData_15 : _GEN_270; // @[Switch.scala 33:19:@1434.4]
  assign _GEN_272 = 5'h10 == select_8 ? io_inData_16 : _GEN_271; // @[Switch.scala 33:19:@1434.4]
  assign _GEN_273 = 5'h11 == select_8 ? io_inData_17 : _GEN_272; // @[Switch.scala 33:19:@1434.4]
  assign _GEN_274 = 5'h12 == select_8 ? io_inData_18 : _GEN_273; // @[Switch.scala 33:19:@1434.4]
  assign _GEN_275 = 5'h13 == select_8 ? io_inData_19 : _GEN_274; // @[Switch.scala 33:19:@1434.4]
  assign _GEN_276 = 5'h14 == select_8 ? io_inData_20 : _GEN_275; // @[Switch.scala 33:19:@1434.4]
  assign _GEN_277 = 5'h15 == select_8 ? io_inData_21 : _GEN_276; // @[Switch.scala 33:19:@1434.4]
  assign _GEN_278 = 5'h16 == select_8 ? io_inData_22 : _GEN_277; // @[Switch.scala 33:19:@1434.4]
  assign _GEN_279 = 5'h17 == select_8 ? io_inData_23 : _GEN_278; // @[Switch.scala 33:19:@1434.4]
  assign _GEN_280 = 5'h18 == select_8 ? io_inData_24 : _GEN_279; // @[Switch.scala 33:19:@1434.4]
  assign _GEN_281 = 5'h19 == select_8 ? io_inData_25 : _GEN_280; // @[Switch.scala 33:19:@1434.4]
  assign _GEN_282 = 5'h1a == select_8 ? io_inData_26 : _GEN_281; // @[Switch.scala 33:19:@1434.4]
  assign _GEN_283 = 5'h1b == select_8 ? io_inData_27 : _GEN_282; // @[Switch.scala 33:19:@1434.4]
  assign _GEN_284 = 5'h1c == select_8 ? io_inData_28 : _GEN_283; // @[Switch.scala 33:19:@1434.4]
  assign _GEN_285 = 5'h1d == select_8 ? io_inData_29 : _GEN_284; // @[Switch.scala 33:19:@1434.4]
  assign _GEN_286 = 5'h1e == select_8 ? io_inData_30 : _GEN_285; // @[Switch.scala 33:19:@1434.4]
  assign _T_6467 = {valid_8_7,valid_8_6,valid_8_5,valid_8_4,valid_8_3,valid_8_2,valid_8_1,valid_8_0}; // @[Switch.scala 34:32:@1441.4]
  assign _T_6475 = {valid_8_15,valid_8_14,valid_8_13,valid_8_12,valid_8_11,valid_8_10,valid_8_9,valid_8_8,_T_6467}; // @[Switch.scala 34:32:@1449.4]
  assign _T_6482 = {valid_8_23,valid_8_22,valid_8_21,valid_8_20,valid_8_19,valid_8_18,valid_8_17,valid_8_16}; // @[Switch.scala 34:32:@1456.4]
  assign _T_6491 = {valid_8_31,valid_8_30,valid_8_29,valid_8_28,valid_8_27,valid_8_26,valid_8_25,valid_8_24,_T_6482,_T_6475}; // @[Switch.scala 34:32:@1465.4]
  assign _T_6495 = io_inAddr_0 == 5'h9; // @[Switch.scala 30:53:@1468.4]
  assign valid_9_0 = io_inValid_0 & _T_6495; // @[Switch.scala 30:36:@1469.4]
  assign _T_6498 = io_inAddr_1 == 5'h9; // @[Switch.scala 30:53:@1471.4]
  assign valid_9_1 = io_inValid_1 & _T_6498; // @[Switch.scala 30:36:@1472.4]
  assign _T_6501 = io_inAddr_2 == 5'h9; // @[Switch.scala 30:53:@1474.4]
  assign valid_9_2 = io_inValid_2 & _T_6501; // @[Switch.scala 30:36:@1475.4]
  assign _T_6504 = io_inAddr_3 == 5'h9; // @[Switch.scala 30:53:@1477.4]
  assign valid_9_3 = io_inValid_3 & _T_6504; // @[Switch.scala 30:36:@1478.4]
  assign _T_6507 = io_inAddr_4 == 5'h9; // @[Switch.scala 30:53:@1480.4]
  assign valid_9_4 = io_inValid_4 & _T_6507; // @[Switch.scala 30:36:@1481.4]
  assign _T_6510 = io_inAddr_5 == 5'h9; // @[Switch.scala 30:53:@1483.4]
  assign valid_9_5 = io_inValid_5 & _T_6510; // @[Switch.scala 30:36:@1484.4]
  assign _T_6513 = io_inAddr_6 == 5'h9; // @[Switch.scala 30:53:@1486.4]
  assign valid_9_6 = io_inValid_6 & _T_6513; // @[Switch.scala 30:36:@1487.4]
  assign _T_6516 = io_inAddr_7 == 5'h9; // @[Switch.scala 30:53:@1489.4]
  assign valid_9_7 = io_inValid_7 & _T_6516; // @[Switch.scala 30:36:@1490.4]
  assign _T_6519 = io_inAddr_8 == 5'h9; // @[Switch.scala 30:53:@1492.4]
  assign valid_9_8 = io_inValid_8 & _T_6519; // @[Switch.scala 30:36:@1493.4]
  assign _T_6522 = io_inAddr_9 == 5'h9; // @[Switch.scala 30:53:@1495.4]
  assign valid_9_9 = io_inValid_9 & _T_6522; // @[Switch.scala 30:36:@1496.4]
  assign _T_6525 = io_inAddr_10 == 5'h9; // @[Switch.scala 30:53:@1498.4]
  assign valid_9_10 = io_inValid_10 & _T_6525; // @[Switch.scala 30:36:@1499.4]
  assign _T_6528 = io_inAddr_11 == 5'h9; // @[Switch.scala 30:53:@1501.4]
  assign valid_9_11 = io_inValid_11 & _T_6528; // @[Switch.scala 30:36:@1502.4]
  assign _T_6531 = io_inAddr_12 == 5'h9; // @[Switch.scala 30:53:@1504.4]
  assign valid_9_12 = io_inValid_12 & _T_6531; // @[Switch.scala 30:36:@1505.4]
  assign _T_6534 = io_inAddr_13 == 5'h9; // @[Switch.scala 30:53:@1507.4]
  assign valid_9_13 = io_inValid_13 & _T_6534; // @[Switch.scala 30:36:@1508.4]
  assign _T_6537 = io_inAddr_14 == 5'h9; // @[Switch.scala 30:53:@1510.4]
  assign valid_9_14 = io_inValid_14 & _T_6537; // @[Switch.scala 30:36:@1511.4]
  assign _T_6540 = io_inAddr_15 == 5'h9; // @[Switch.scala 30:53:@1513.4]
  assign valid_9_15 = io_inValid_15 & _T_6540; // @[Switch.scala 30:36:@1514.4]
  assign _T_6543 = io_inAddr_16 == 5'h9; // @[Switch.scala 30:53:@1516.4]
  assign valid_9_16 = io_inValid_16 & _T_6543; // @[Switch.scala 30:36:@1517.4]
  assign _T_6546 = io_inAddr_17 == 5'h9; // @[Switch.scala 30:53:@1519.4]
  assign valid_9_17 = io_inValid_17 & _T_6546; // @[Switch.scala 30:36:@1520.4]
  assign _T_6549 = io_inAddr_18 == 5'h9; // @[Switch.scala 30:53:@1522.4]
  assign valid_9_18 = io_inValid_18 & _T_6549; // @[Switch.scala 30:36:@1523.4]
  assign _T_6552 = io_inAddr_19 == 5'h9; // @[Switch.scala 30:53:@1525.4]
  assign valid_9_19 = io_inValid_19 & _T_6552; // @[Switch.scala 30:36:@1526.4]
  assign _T_6555 = io_inAddr_20 == 5'h9; // @[Switch.scala 30:53:@1528.4]
  assign valid_9_20 = io_inValid_20 & _T_6555; // @[Switch.scala 30:36:@1529.4]
  assign _T_6558 = io_inAddr_21 == 5'h9; // @[Switch.scala 30:53:@1531.4]
  assign valid_9_21 = io_inValid_21 & _T_6558; // @[Switch.scala 30:36:@1532.4]
  assign _T_6561 = io_inAddr_22 == 5'h9; // @[Switch.scala 30:53:@1534.4]
  assign valid_9_22 = io_inValid_22 & _T_6561; // @[Switch.scala 30:36:@1535.4]
  assign _T_6564 = io_inAddr_23 == 5'h9; // @[Switch.scala 30:53:@1537.4]
  assign valid_9_23 = io_inValid_23 & _T_6564; // @[Switch.scala 30:36:@1538.4]
  assign _T_6567 = io_inAddr_24 == 5'h9; // @[Switch.scala 30:53:@1540.4]
  assign valid_9_24 = io_inValid_24 & _T_6567; // @[Switch.scala 30:36:@1541.4]
  assign _T_6570 = io_inAddr_25 == 5'h9; // @[Switch.scala 30:53:@1543.4]
  assign valid_9_25 = io_inValid_25 & _T_6570; // @[Switch.scala 30:36:@1544.4]
  assign _T_6573 = io_inAddr_26 == 5'h9; // @[Switch.scala 30:53:@1546.4]
  assign valid_9_26 = io_inValid_26 & _T_6573; // @[Switch.scala 30:36:@1547.4]
  assign _T_6576 = io_inAddr_27 == 5'h9; // @[Switch.scala 30:53:@1549.4]
  assign valid_9_27 = io_inValid_27 & _T_6576; // @[Switch.scala 30:36:@1550.4]
  assign _T_6579 = io_inAddr_28 == 5'h9; // @[Switch.scala 30:53:@1552.4]
  assign valid_9_28 = io_inValid_28 & _T_6579; // @[Switch.scala 30:36:@1553.4]
  assign _T_6582 = io_inAddr_29 == 5'h9; // @[Switch.scala 30:53:@1555.4]
  assign valid_9_29 = io_inValid_29 & _T_6582; // @[Switch.scala 30:36:@1556.4]
  assign _T_6585 = io_inAddr_30 == 5'h9; // @[Switch.scala 30:53:@1558.4]
  assign valid_9_30 = io_inValid_30 & _T_6585; // @[Switch.scala 30:36:@1559.4]
  assign _T_6588 = io_inAddr_31 == 5'h9; // @[Switch.scala 30:53:@1561.4]
  assign valid_9_31 = io_inValid_31 & _T_6588; // @[Switch.scala 30:36:@1562.4]
  assign _T_6622 = valid_9_30 ? 5'h1e : 5'h1f; // @[Mux.scala 31:69:@1564.4]
  assign _T_6623 = valid_9_29 ? 5'h1d : _T_6622; // @[Mux.scala 31:69:@1565.4]
  assign _T_6624 = valid_9_28 ? 5'h1c : _T_6623; // @[Mux.scala 31:69:@1566.4]
  assign _T_6625 = valid_9_27 ? 5'h1b : _T_6624; // @[Mux.scala 31:69:@1567.4]
  assign _T_6626 = valid_9_26 ? 5'h1a : _T_6625; // @[Mux.scala 31:69:@1568.4]
  assign _T_6627 = valid_9_25 ? 5'h19 : _T_6626; // @[Mux.scala 31:69:@1569.4]
  assign _T_6628 = valid_9_24 ? 5'h18 : _T_6627; // @[Mux.scala 31:69:@1570.4]
  assign _T_6629 = valid_9_23 ? 5'h17 : _T_6628; // @[Mux.scala 31:69:@1571.4]
  assign _T_6630 = valid_9_22 ? 5'h16 : _T_6629; // @[Mux.scala 31:69:@1572.4]
  assign _T_6631 = valid_9_21 ? 5'h15 : _T_6630; // @[Mux.scala 31:69:@1573.4]
  assign _T_6632 = valid_9_20 ? 5'h14 : _T_6631; // @[Mux.scala 31:69:@1574.4]
  assign _T_6633 = valid_9_19 ? 5'h13 : _T_6632; // @[Mux.scala 31:69:@1575.4]
  assign _T_6634 = valid_9_18 ? 5'h12 : _T_6633; // @[Mux.scala 31:69:@1576.4]
  assign _T_6635 = valid_9_17 ? 5'h11 : _T_6634; // @[Mux.scala 31:69:@1577.4]
  assign _T_6636 = valid_9_16 ? 5'h10 : _T_6635; // @[Mux.scala 31:69:@1578.4]
  assign _T_6637 = valid_9_15 ? 5'hf : _T_6636; // @[Mux.scala 31:69:@1579.4]
  assign _T_6638 = valid_9_14 ? 5'he : _T_6637; // @[Mux.scala 31:69:@1580.4]
  assign _T_6639 = valid_9_13 ? 5'hd : _T_6638; // @[Mux.scala 31:69:@1581.4]
  assign _T_6640 = valid_9_12 ? 5'hc : _T_6639; // @[Mux.scala 31:69:@1582.4]
  assign _T_6641 = valid_9_11 ? 5'hb : _T_6640; // @[Mux.scala 31:69:@1583.4]
  assign _T_6642 = valid_9_10 ? 5'ha : _T_6641; // @[Mux.scala 31:69:@1584.4]
  assign _T_6643 = valid_9_9 ? 5'h9 : _T_6642; // @[Mux.scala 31:69:@1585.4]
  assign _T_6644 = valid_9_8 ? 5'h8 : _T_6643; // @[Mux.scala 31:69:@1586.4]
  assign _T_6645 = valid_9_7 ? 5'h7 : _T_6644; // @[Mux.scala 31:69:@1587.4]
  assign _T_6646 = valid_9_6 ? 5'h6 : _T_6645; // @[Mux.scala 31:69:@1588.4]
  assign _T_6647 = valid_9_5 ? 5'h5 : _T_6646; // @[Mux.scala 31:69:@1589.4]
  assign _T_6648 = valid_9_4 ? 5'h4 : _T_6647; // @[Mux.scala 31:69:@1590.4]
  assign _T_6649 = valid_9_3 ? 5'h3 : _T_6648; // @[Mux.scala 31:69:@1591.4]
  assign _T_6650 = valid_9_2 ? 5'h2 : _T_6649; // @[Mux.scala 31:69:@1592.4]
  assign _T_6651 = valid_9_1 ? 5'h1 : _T_6650; // @[Mux.scala 31:69:@1593.4]
  assign select_9 = valid_9_0 ? 5'h0 : _T_6651; // @[Mux.scala 31:69:@1594.4]
  assign _GEN_289 = 5'h1 == select_9 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@1596.4]
  assign _GEN_290 = 5'h2 == select_9 ? io_inData_2 : _GEN_289; // @[Switch.scala 33:19:@1596.4]
  assign _GEN_291 = 5'h3 == select_9 ? io_inData_3 : _GEN_290; // @[Switch.scala 33:19:@1596.4]
  assign _GEN_292 = 5'h4 == select_9 ? io_inData_4 : _GEN_291; // @[Switch.scala 33:19:@1596.4]
  assign _GEN_293 = 5'h5 == select_9 ? io_inData_5 : _GEN_292; // @[Switch.scala 33:19:@1596.4]
  assign _GEN_294 = 5'h6 == select_9 ? io_inData_6 : _GEN_293; // @[Switch.scala 33:19:@1596.4]
  assign _GEN_295 = 5'h7 == select_9 ? io_inData_7 : _GEN_294; // @[Switch.scala 33:19:@1596.4]
  assign _GEN_296 = 5'h8 == select_9 ? io_inData_8 : _GEN_295; // @[Switch.scala 33:19:@1596.4]
  assign _GEN_297 = 5'h9 == select_9 ? io_inData_9 : _GEN_296; // @[Switch.scala 33:19:@1596.4]
  assign _GEN_298 = 5'ha == select_9 ? io_inData_10 : _GEN_297; // @[Switch.scala 33:19:@1596.4]
  assign _GEN_299 = 5'hb == select_9 ? io_inData_11 : _GEN_298; // @[Switch.scala 33:19:@1596.4]
  assign _GEN_300 = 5'hc == select_9 ? io_inData_12 : _GEN_299; // @[Switch.scala 33:19:@1596.4]
  assign _GEN_301 = 5'hd == select_9 ? io_inData_13 : _GEN_300; // @[Switch.scala 33:19:@1596.4]
  assign _GEN_302 = 5'he == select_9 ? io_inData_14 : _GEN_301; // @[Switch.scala 33:19:@1596.4]
  assign _GEN_303 = 5'hf == select_9 ? io_inData_15 : _GEN_302; // @[Switch.scala 33:19:@1596.4]
  assign _GEN_304 = 5'h10 == select_9 ? io_inData_16 : _GEN_303; // @[Switch.scala 33:19:@1596.4]
  assign _GEN_305 = 5'h11 == select_9 ? io_inData_17 : _GEN_304; // @[Switch.scala 33:19:@1596.4]
  assign _GEN_306 = 5'h12 == select_9 ? io_inData_18 : _GEN_305; // @[Switch.scala 33:19:@1596.4]
  assign _GEN_307 = 5'h13 == select_9 ? io_inData_19 : _GEN_306; // @[Switch.scala 33:19:@1596.4]
  assign _GEN_308 = 5'h14 == select_9 ? io_inData_20 : _GEN_307; // @[Switch.scala 33:19:@1596.4]
  assign _GEN_309 = 5'h15 == select_9 ? io_inData_21 : _GEN_308; // @[Switch.scala 33:19:@1596.4]
  assign _GEN_310 = 5'h16 == select_9 ? io_inData_22 : _GEN_309; // @[Switch.scala 33:19:@1596.4]
  assign _GEN_311 = 5'h17 == select_9 ? io_inData_23 : _GEN_310; // @[Switch.scala 33:19:@1596.4]
  assign _GEN_312 = 5'h18 == select_9 ? io_inData_24 : _GEN_311; // @[Switch.scala 33:19:@1596.4]
  assign _GEN_313 = 5'h19 == select_9 ? io_inData_25 : _GEN_312; // @[Switch.scala 33:19:@1596.4]
  assign _GEN_314 = 5'h1a == select_9 ? io_inData_26 : _GEN_313; // @[Switch.scala 33:19:@1596.4]
  assign _GEN_315 = 5'h1b == select_9 ? io_inData_27 : _GEN_314; // @[Switch.scala 33:19:@1596.4]
  assign _GEN_316 = 5'h1c == select_9 ? io_inData_28 : _GEN_315; // @[Switch.scala 33:19:@1596.4]
  assign _GEN_317 = 5'h1d == select_9 ? io_inData_29 : _GEN_316; // @[Switch.scala 33:19:@1596.4]
  assign _GEN_318 = 5'h1e == select_9 ? io_inData_30 : _GEN_317; // @[Switch.scala 33:19:@1596.4]
  assign _T_6660 = {valid_9_7,valid_9_6,valid_9_5,valid_9_4,valid_9_3,valid_9_2,valid_9_1,valid_9_0}; // @[Switch.scala 34:32:@1603.4]
  assign _T_6668 = {valid_9_15,valid_9_14,valid_9_13,valid_9_12,valid_9_11,valid_9_10,valid_9_9,valid_9_8,_T_6660}; // @[Switch.scala 34:32:@1611.4]
  assign _T_6675 = {valid_9_23,valid_9_22,valid_9_21,valid_9_20,valid_9_19,valid_9_18,valid_9_17,valid_9_16}; // @[Switch.scala 34:32:@1618.4]
  assign _T_6684 = {valid_9_31,valid_9_30,valid_9_29,valid_9_28,valid_9_27,valid_9_26,valid_9_25,valid_9_24,_T_6675,_T_6668}; // @[Switch.scala 34:32:@1627.4]
  assign _T_6688 = io_inAddr_0 == 5'ha; // @[Switch.scala 30:53:@1630.4]
  assign valid_10_0 = io_inValid_0 & _T_6688; // @[Switch.scala 30:36:@1631.4]
  assign _T_6691 = io_inAddr_1 == 5'ha; // @[Switch.scala 30:53:@1633.4]
  assign valid_10_1 = io_inValid_1 & _T_6691; // @[Switch.scala 30:36:@1634.4]
  assign _T_6694 = io_inAddr_2 == 5'ha; // @[Switch.scala 30:53:@1636.4]
  assign valid_10_2 = io_inValid_2 & _T_6694; // @[Switch.scala 30:36:@1637.4]
  assign _T_6697 = io_inAddr_3 == 5'ha; // @[Switch.scala 30:53:@1639.4]
  assign valid_10_3 = io_inValid_3 & _T_6697; // @[Switch.scala 30:36:@1640.4]
  assign _T_6700 = io_inAddr_4 == 5'ha; // @[Switch.scala 30:53:@1642.4]
  assign valid_10_4 = io_inValid_4 & _T_6700; // @[Switch.scala 30:36:@1643.4]
  assign _T_6703 = io_inAddr_5 == 5'ha; // @[Switch.scala 30:53:@1645.4]
  assign valid_10_5 = io_inValid_5 & _T_6703; // @[Switch.scala 30:36:@1646.4]
  assign _T_6706 = io_inAddr_6 == 5'ha; // @[Switch.scala 30:53:@1648.4]
  assign valid_10_6 = io_inValid_6 & _T_6706; // @[Switch.scala 30:36:@1649.4]
  assign _T_6709 = io_inAddr_7 == 5'ha; // @[Switch.scala 30:53:@1651.4]
  assign valid_10_7 = io_inValid_7 & _T_6709; // @[Switch.scala 30:36:@1652.4]
  assign _T_6712 = io_inAddr_8 == 5'ha; // @[Switch.scala 30:53:@1654.4]
  assign valid_10_8 = io_inValid_8 & _T_6712; // @[Switch.scala 30:36:@1655.4]
  assign _T_6715 = io_inAddr_9 == 5'ha; // @[Switch.scala 30:53:@1657.4]
  assign valid_10_9 = io_inValid_9 & _T_6715; // @[Switch.scala 30:36:@1658.4]
  assign _T_6718 = io_inAddr_10 == 5'ha; // @[Switch.scala 30:53:@1660.4]
  assign valid_10_10 = io_inValid_10 & _T_6718; // @[Switch.scala 30:36:@1661.4]
  assign _T_6721 = io_inAddr_11 == 5'ha; // @[Switch.scala 30:53:@1663.4]
  assign valid_10_11 = io_inValid_11 & _T_6721; // @[Switch.scala 30:36:@1664.4]
  assign _T_6724 = io_inAddr_12 == 5'ha; // @[Switch.scala 30:53:@1666.4]
  assign valid_10_12 = io_inValid_12 & _T_6724; // @[Switch.scala 30:36:@1667.4]
  assign _T_6727 = io_inAddr_13 == 5'ha; // @[Switch.scala 30:53:@1669.4]
  assign valid_10_13 = io_inValid_13 & _T_6727; // @[Switch.scala 30:36:@1670.4]
  assign _T_6730 = io_inAddr_14 == 5'ha; // @[Switch.scala 30:53:@1672.4]
  assign valid_10_14 = io_inValid_14 & _T_6730; // @[Switch.scala 30:36:@1673.4]
  assign _T_6733 = io_inAddr_15 == 5'ha; // @[Switch.scala 30:53:@1675.4]
  assign valid_10_15 = io_inValid_15 & _T_6733; // @[Switch.scala 30:36:@1676.4]
  assign _T_6736 = io_inAddr_16 == 5'ha; // @[Switch.scala 30:53:@1678.4]
  assign valid_10_16 = io_inValid_16 & _T_6736; // @[Switch.scala 30:36:@1679.4]
  assign _T_6739 = io_inAddr_17 == 5'ha; // @[Switch.scala 30:53:@1681.4]
  assign valid_10_17 = io_inValid_17 & _T_6739; // @[Switch.scala 30:36:@1682.4]
  assign _T_6742 = io_inAddr_18 == 5'ha; // @[Switch.scala 30:53:@1684.4]
  assign valid_10_18 = io_inValid_18 & _T_6742; // @[Switch.scala 30:36:@1685.4]
  assign _T_6745 = io_inAddr_19 == 5'ha; // @[Switch.scala 30:53:@1687.4]
  assign valid_10_19 = io_inValid_19 & _T_6745; // @[Switch.scala 30:36:@1688.4]
  assign _T_6748 = io_inAddr_20 == 5'ha; // @[Switch.scala 30:53:@1690.4]
  assign valid_10_20 = io_inValid_20 & _T_6748; // @[Switch.scala 30:36:@1691.4]
  assign _T_6751 = io_inAddr_21 == 5'ha; // @[Switch.scala 30:53:@1693.4]
  assign valid_10_21 = io_inValid_21 & _T_6751; // @[Switch.scala 30:36:@1694.4]
  assign _T_6754 = io_inAddr_22 == 5'ha; // @[Switch.scala 30:53:@1696.4]
  assign valid_10_22 = io_inValid_22 & _T_6754; // @[Switch.scala 30:36:@1697.4]
  assign _T_6757 = io_inAddr_23 == 5'ha; // @[Switch.scala 30:53:@1699.4]
  assign valid_10_23 = io_inValid_23 & _T_6757; // @[Switch.scala 30:36:@1700.4]
  assign _T_6760 = io_inAddr_24 == 5'ha; // @[Switch.scala 30:53:@1702.4]
  assign valid_10_24 = io_inValid_24 & _T_6760; // @[Switch.scala 30:36:@1703.4]
  assign _T_6763 = io_inAddr_25 == 5'ha; // @[Switch.scala 30:53:@1705.4]
  assign valid_10_25 = io_inValid_25 & _T_6763; // @[Switch.scala 30:36:@1706.4]
  assign _T_6766 = io_inAddr_26 == 5'ha; // @[Switch.scala 30:53:@1708.4]
  assign valid_10_26 = io_inValid_26 & _T_6766; // @[Switch.scala 30:36:@1709.4]
  assign _T_6769 = io_inAddr_27 == 5'ha; // @[Switch.scala 30:53:@1711.4]
  assign valid_10_27 = io_inValid_27 & _T_6769; // @[Switch.scala 30:36:@1712.4]
  assign _T_6772 = io_inAddr_28 == 5'ha; // @[Switch.scala 30:53:@1714.4]
  assign valid_10_28 = io_inValid_28 & _T_6772; // @[Switch.scala 30:36:@1715.4]
  assign _T_6775 = io_inAddr_29 == 5'ha; // @[Switch.scala 30:53:@1717.4]
  assign valid_10_29 = io_inValid_29 & _T_6775; // @[Switch.scala 30:36:@1718.4]
  assign _T_6778 = io_inAddr_30 == 5'ha; // @[Switch.scala 30:53:@1720.4]
  assign valid_10_30 = io_inValid_30 & _T_6778; // @[Switch.scala 30:36:@1721.4]
  assign _T_6781 = io_inAddr_31 == 5'ha; // @[Switch.scala 30:53:@1723.4]
  assign valid_10_31 = io_inValid_31 & _T_6781; // @[Switch.scala 30:36:@1724.4]
  assign _T_6815 = valid_10_30 ? 5'h1e : 5'h1f; // @[Mux.scala 31:69:@1726.4]
  assign _T_6816 = valid_10_29 ? 5'h1d : _T_6815; // @[Mux.scala 31:69:@1727.4]
  assign _T_6817 = valid_10_28 ? 5'h1c : _T_6816; // @[Mux.scala 31:69:@1728.4]
  assign _T_6818 = valid_10_27 ? 5'h1b : _T_6817; // @[Mux.scala 31:69:@1729.4]
  assign _T_6819 = valid_10_26 ? 5'h1a : _T_6818; // @[Mux.scala 31:69:@1730.4]
  assign _T_6820 = valid_10_25 ? 5'h19 : _T_6819; // @[Mux.scala 31:69:@1731.4]
  assign _T_6821 = valid_10_24 ? 5'h18 : _T_6820; // @[Mux.scala 31:69:@1732.4]
  assign _T_6822 = valid_10_23 ? 5'h17 : _T_6821; // @[Mux.scala 31:69:@1733.4]
  assign _T_6823 = valid_10_22 ? 5'h16 : _T_6822; // @[Mux.scala 31:69:@1734.4]
  assign _T_6824 = valid_10_21 ? 5'h15 : _T_6823; // @[Mux.scala 31:69:@1735.4]
  assign _T_6825 = valid_10_20 ? 5'h14 : _T_6824; // @[Mux.scala 31:69:@1736.4]
  assign _T_6826 = valid_10_19 ? 5'h13 : _T_6825; // @[Mux.scala 31:69:@1737.4]
  assign _T_6827 = valid_10_18 ? 5'h12 : _T_6826; // @[Mux.scala 31:69:@1738.4]
  assign _T_6828 = valid_10_17 ? 5'h11 : _T_6827; // @[Mux.scala 31:69:@1739.4]
  assign _T_6829 = valid_10_16 ? 5'h10 : _T_6828; // @[Mux.scala 31:69:@1740.4]
  assign _T_6830 = valid_10_15 ? 5'hf : _T_6829; // @[Mux.scala 31:69:@1741.4]
  assign _T_6831 = valid_10_14 ? 5'he : _T_6830; // @[Mux.scala 31:69:@1742.4]
  assign _T_6832 = valid_10_13 ? 5'hd : _T_6831; // @[Mux.scala 31:69:@1743.4]
  assign _T_6833 = valid_10_12 ? 5'hc : _T_6832; // @[Mux.scala 31:69:@1744.4]
  assign _T_6834 = valid_10_11 ? 5'hb : _T_6833; // @[Mux.scala 31:69:@1745.4]
  assign _T_6835 = valid_10_10 ? 5'ha : _T_6834; // @[Mux.scala 31:69:@1746.4]
  assign _T_6836 = valid_10_9 ? 5'h9 : _T_6835; // @[Mux.scala 31:69:@1747.4]
  assign _T_6837 = valid_10_8 ? 5'h8 : _T_6836; // @[Mux.scala 31:69:@1748.4]
  assign _T_6838 = valid_10_7 ? 5'h7 : _T_6837; // @[Mux.scala 31:69:@1749.4]
  assign _T_6839 = valid_10_6 ? 5'h6 : _T_6838; // @[Mux.scala 31:69:@1750.4]
  assign _T_6840 = valid_10_5 ? 5'h5 : _T_6839; // @[Mux.scala 31:69:@1751.4]
  assign _T_6841 = valid_10_4 ? 5'h4 : _T_6840; // @[Mux.scala 31:69:@1752.4]
  assign _T_6842 = valid_10_3 ? 5'h3 : _T_6841; // @[Mux.scala 31:69:@1753.4]
  assign _T_6843 = valid_10_2 ? 5'h2 : _T_6842; // @[Mux.scala 31:69:@1754.4]
  assign _T_6844 = valid_10_1 ? 5'h1 : _T_6843; // @[Mux.scala 31:69:@1755.4]
  assign select_10 = valid_10_0 ? 5'h0 : _T_6844; // @[Mux.scala 31:69:@1756.4]
  assign _GEN_321 = 5'h1 == select_10 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@1758.4]
  assign _GEN_322 = 5'h2 == select_10 ? io_inData_2 : _GEN_321; // @[Switch.scala 33:19:@1758.4]
  assign _GEN_323 = 5'h3 == select_10 ? io_inData_3 : _GEN_322; // @[Switch.scala 33:19:@1758.4]
  assign _GEN_324 = 5'h4 == select_10 ? io_inData_4 : _GEN_323; // @[Switch.scala 33:19:@1758.4]
  assign _GEN_325 = 5'h5 == select_10 ? io_inData_5 : _GEN_324; // @[Switch.scala 33:19:@1758.4]
  assign _GEN_326 = 5'h6 == select_10 ? io_inData_6 : _GEN_325; // @[Switch.scala 33:19:@1758.4]
  assign _GEN_327 = 5'h7 == select_10 ? io_inData_7 : _GEN_326; // @[Switch.scala 33:19:@1758.4]
  assign _GEN_328 = 5'h8 == select_10 ? io_inData_8 : _GEN_327; // @[Switch.scala 33:19:@1758.4]
  assign _GEN_329 = 5'h9 == select_10 ? io_inData_9 : _GEN_328; // @[Switch.scala 33:19:@1758.4]
  assign _GEN_330 = 5'ha == select_10 ? io_inData_10 : _GEN_329; // @[Switch.scala 33:19:@1758.4]
  assign _GEN_331 = 5'hb == select_10 ? io_inData_11 : _GEN_330; // @[Switch.scala 33:19:@1758.4]
  assign _GEN_332 = 5'hc == select_10 ? io_inData_12 : _GEN_331; // @[Switch.scala 33:19:@1758.4]
  assign _GEN_333 = 5'hd == select_10 ? io_inData_13 : _GEN_332; // @[Switch.scala 33:19:@1758.4]
  assign _GEN_334 = 5'he == select_10 ? io_inData_14 : _GEN_333; // @[Switch.scala 33:19:@1758.4]
  assign _GEN_335 = 5'hf == select_10 ? io_inData_15 : _GEN_334; // @[Switch.scala 33:19:@1758.4]
  assign _GEN_336 = 5'h10 == select_10 ? io_inData_16 : _GEN_335; // @[Switch.scala 33:19:@1758.4]
  assign _GEN_337 = 5'h11 == select_10 ? io_inData_17 : _GEN_336; // @[Switch.scala 33:19:@1758.4]
  assign _GEN_338 = 5'h12 == select_10 ? io_inData_18 : _GEN_337; // @[Switch.scala 33:19:@1758.4]
  assign _GEN_339 = 5'h13 == select_10 ? io_inData_19 : _GEN_338; // @[Switch.scala 33:19:@1758.4]
  assign _GEN_340 = 5'h14 == select_10 ? io_inData_20 : _GEN_339; // @[Switch.scala 33:19:@1758.4]
  assign _GEN_341 = 5'h15 == select_10 ? io_inData_21 : _GEN_340; // @[Switch.scala 33:19:@1758.4]
  assign _GEN_342 = 5'h16 == select_10 ? io_inData_22 : _GEN_341; // @[Switch.scala 33:19:@1758.4]
  assign _GEN_343 = 5'h17 == select_10 ? io_inData_23 : _GEN_342; // @[Switch.scala 33:19:@1758.4]
  assign _GEN_344 = 5'h18 == select_10 ? io_inData_24 : _GEN_343; // @[Switch.scala 33:19:@1758.4]
  assign _GEN_345 = 5'h19 == select_10 ? io_inData_25 : _GEN_344; // @[Switch.scala 33:19:@1758.4]
  assign _GEN_346 = 5'h1a == select_10 ? io_inData_26 : _GEN_345; // @[Switch.scala 33:19:@1758.4]
  assign _GEN_347 = 5'h1b == select_10 ? io_inData_27 : _GEN_346; // @[Switch.scala 33:19:@1758.4]
  assign _GEN_348 = 5'h1c == select_10 ? io_inData_28 : _GEN_347; // @[Switch.scala 33:19:@1758.4]
  assign _GEN_349 = 5'h1d == select_10 ? io_inData_29 : _GEN_348; // @[Switch.scala 33:19:@1758.4]
  assign _GEN_350 = 5'h1e == select_10 ? io_inData_30 : _GEN_349; // @[Switch.scala 33:19:@1758.4]
  assign _T_6853 = {valid_10_7,valid_10_6,valid_10_5,valid_10_4,valid_10_3,valid_10_2,valid_10_1,valid_10_0}; // @[Switch.scala 34:32:@1765.4]
  assign _T_6861 = {valid_10_15,valid_10_14,valid_10_13,valid_10_12,valid_10_11,valid_10_10,valid_10_9,valid_10_8,_T_6853}; // @[Switch.scala 34:32:@1773.4]
  assign _T_6868 = {valid_10_23,valid_10_22,valid_10_21,valid_10_20,valid_10_19,valid_10_18,valid_10_17,valid_10_16}; // @[Switch.scala 34:32:@1780.4]
  assign _T_6877 = {valid_10_31,valid_10_30,valid_10_29,valid_10_28,valid_10_27,valid_10_26,valid_10_25,valid_10_24,_T_6868,_T_6861}; // @[Switch.scala 34:32:@1789.4]
  assign _T_6881 = io_inAddr_0 == 5'hb; // @[Switch.scala 30:53:@1792.4]
  assign valid_11_0 = io_inValid_0 & _T_6881; // @[Switch.scala 30:36:@1793.4]
  assign _T_6884 = io_inAddr_1 == 5'hb; // @[Switch.scala 30:53:@1795.4]
  assign valid_11_1 = io_inValid_1 & _T_6884; // @[Switch.scala 30:36:@1796.4]
  assign _T_6887 = io_inAddr_2 == 5'hb; // @[Switch.scala 30:53:@1798.4]
  assign valid_11_2 = io_inValid_2 & _T_6887; // @[Switch.scala 30:36:@1799.4]
  assign _T_6890 = io_inAddr_3 == 5'hb; // @[Switch.scala 30:53:@1801.4]
  assign valid_11_3 = io_inValid_3 & _T_6890; // @[Switch.scala 30:36:@1802.4]
  assign _T_6893 = io_inAddr_4 == 5'hb; // @[Switch.scala 30:53:@1804.4]
  assign valid_11_4 = io_inValid_4 & _T_6893; // @[Switch.scala 30:36:@1805.4]
  assign _T_6896 = io_inAddr_5 == 5'hb; // @[Switch.scala 30:53:@1807.4]
  assign valid_11_5 = io_inValid_5 & _T_6896; // @[Switch.scala 30:36:@1808.4]
  assign _T_6899 = io_inAddr_6 == 5'hb; // @[Switch.scala 30:53:@1810.4]
  assign valid_11_6 = io_inValid_6 & _T_6899; // @[Switch.scala 30:36:@1811.4]
  assign _T_6902 = io_inAddr_7 == 5'hb; // @[Switch.scala 30:53:@1813.4]
  assign valid_11_7 = io_inValid_7 & _T_6902; // @[Switch.scala 30:36:@1814.4]
  assign _T_6905 = io_inAddr_8 == 5'hb; // @[Switch.scala 30:53:@1816.4]
  assign valid_11_8 = io_inValid_8 & _T_6905; // @[Switch.scala 30:36:@1817.4]
  assign _T_6908 = io_inAddr_9 == 5'hb; // @[Switch.scala 30:53:@1819.4]
  assign valid_11_9 = io_inValid_9 & _T_6908; // @[Switch.scala 30:36:@1820.4]
  assign _T_6911 = io_inAddr_10 == 5'hb; // @[Switch.scala 30:53:@1822.4]
  assign valid_11_10 = io_inValid_10 & _T_6911; // @[Switch.scala 30:36:@1823.4]
  assign _T_6914 = io_inAddr_11 == 5'hb; // @[Switch.scala 30:53:@1825.4]
  assign valid_11_11 = io_inValid_11 & _T_6914; // @[Switch.scala 30:36:@1826.4]
  assign _T_6917 = io_inAddr_12 == 5'hb; // @[Switch.scala 30:53:@1828.4]
  assign valid_11_12 = io_inValid_12 & _T_6917; // @[Switch.scala 30:36:@1829.4]
  assign _T_6920 = io_inAddr_13 == 5'hb; // @[Switch.scala 30:53:@1831.4]
  assign valid_11_13 = io_inValid_13 & _T_6920; // @[Switch.scala 30:36:@1832.4]
  assign _T_6923 = io_inAddr_14 == 5'hb; // @[Switch.scala 30:53:@1834.4]
  assign valid_11_14 = io_inValid_14 & _T_6923; // @[Switch.scala 30:36:@1835.4]
  assign _T_6926 = io_inAddr_15 == 5'hb; // @[Switch.scala 30:53:@1837.4]
  assign valid_11_15 = io_inValid_15 & _T_6926; // @[Switch.scala 30:36:@1838.4]
  assign _T_6929 = io_inAddr_16 == 5'hb; // @[Switch.scala 30:53:@1840.4]
  assign valid_11_16 = io_inValid_16 & _T_6929; // @[Switch.scala 30:36:@1841.4]
  assign _T_6932 = io_inAddr_17 == 5'hb; // @[Switch.scala 30:53:@1843.4]
  assign valid_11_17 = io_inValid_17 & _T_6932; // @[Switch.scala 30:36:@1844.4]
  assign _T_6935 = io_inAddr_18 == 5'hb; // @[Switch.scala 30:53:@1846.4]
  assign valid_11_18 = io_inValid_18 & _T_6935; // @[Switch.scala 30:36:@1847.4]
  assign _T_6938 = io_inAddr_19 == 5'hb; // @[Switch.scala 30:53:@1849.4]
  assign valid_11_19 = io_inValid_19 & _T_6938; // @[Switch.scala 30:36:@1850.4]
  assign _T_6941 = io_inAddr_20 == 5'hb; // @[Switch.scala 30:53:@1852.4]
  assign valid_11_20 = io_inValid_20 & _T_6941; // @[Switch.scala 30:36:@1853.4]
  assign _T_6944 = io_inAddr_21 == 5'hb; // @[Switch.scala 30:53:@1855.4]
  assign valid_11_21 = io_inValid_21 & _T_6944; // @[Switch.scala 30:36:@1856.4]
  assign _T_6947 = io_inAddr_22 == 5'hb; // @[Switch.scala 30:53:@1858.4]
  assign valid_11_22 = io_inValid_22 & _T_6947; // @[Switch.scala 30:36:@1859.4]
  assign _T_6950 = io_inAddr_23 == 5'hb; // @[Switch.scala 30:53:@1861.4]
  assign valid_11_23 = io_inValid_23 & _T_6950; // @[Switch.scala 30:36:@1862.4]
  assign _T_6953 = io_inAddr_24 == 5'hb; // @[Switch.scala 30:53:@1864.4]
  assign valid_11_24 = io_inValid_24 & _T_6953; // @[Switch.scala 30:36:@1865.4]
  assign _T_6956 = io_inAddr_25 == 5'hb; // @[Switch.scala 30:53:@1867.4]
  assign valid_11_25 = io_inValid_25 & _T_6956; // @[Switch.scala 30:36:@1868.4]
  assign _T_6959 = io_inAddr_26 == 5'hb; // @[Switch.scala 30:53:@1870.4]
  assign valid_11_26 = io_inValid_26 & _T_6959; // @[Switch.scala 30:36:@1871.4]
  assign _T_6962 = io_inAddr_27 == 5'hb; // @[Switch.scala 30:53:@1873.4]
  assign valid_11_27 = io_inValid_27 & _T_6962; // @[Switch.scala 30:36:@1874.4]
  assign _T_6965 = io_inAddr_28 == 5'hb; // @[Switch.scala 30:53:@1876.4]
  assign valid_11_28 = io_inValid_28 & _T_6965; // @[Switch.scala 30:36:@1877.4]
  assign _T_6968 = io_inAddr_29 == 5'hb; // @[Switch.scala 30:53:@1879.4]
  assign valid_11_29 = io_inValid_29 & _T_6968; // @[Switch.scala 30:36:@1880.4]
  assign _T_6971 = io_inAddr_30 == 5'hb; // @[Switch.scala 30:53:@1882.4]
  assign valid_11_30 = io_inValid_30 & _T_6971; // @[Switch.scala 30:36:@1883.4]
  assign _T_6974 = io_inAddr_31 == 5'hb; // @[Switch.scala 30:53:@1885.4]
  assign valid_11_31 = io_inValid_31 & _T_6974; // @[Switch.scala 30:36:@1886.4]
  assign _T_7008 = valid_11_30 ? 5'h1e : 5'h1f; // @[Mux.scala 31:69:@1888.4]
  assign _T_7009 = valid_11_29 ? 5'h1d : _T_7008; // @[Mux.scala 31:69:@1889.4]
  assign _T_7010 = valid_11_28 ? 5'h1c : _T_7009; // @[Mux.scala 31:69:@1890.4]
  assign _T_7011 = valid_11_27 ? 5'h1b : _T_7010; // @[Mux.scala 31:69:@1891.4]
  assign _T_7012 = valid_11_26 ? 5'h1a : _T_7011; // @[Mux.scala 31:69:@1892.4]
  assign _T_7013 = valid_11_25 ? 5'h19 : _T_7012; // @[Mux.scala 31:69:@1893.4]
  assign _T_7014 = valid_11_24 ? 5'h18 : _T_7013; // @[Mux.scala 31:69:@1894.4]
  assign _T_7015 = valid_11_23 ? 5'h17 : _T_7014; // @[Mux.scala 31:69:@1895.4]
  assign _T_7016 = valid_11_22 ? 5'h16 : _T_7015; // @[Mux.scala 31:69:@1896.4]
  assign _T_7017 = valid_11_21 ? 5'h15 : _T_7016; // @[Mux.scala 31:69:@1897.4]
  assign _T_7018 = valid_11_20 ? 5'h14 : _T_7017; // @[Mux.scala 31:69:@1898.4]
  assign _T_7019 = valid_11_19 ? 5'h13 : _T_7018; // @[Mux.scala 31:69:@1899.4]
  assign _T_7020 = valid_11_18 ? 5'h12 : _T_7019; // @[Mux.scala 31:69:@1900.4]
  assign _T_7021 = valid_11_17 ? 5'h11 : _T_7020; // @[Mux.scala 31:69:@1901.4]
  assign _T_7022 = valid_11_16 ? 5'h10 : _T_7021; // @[Mux.scala 31:69:@1902.4]
  assign _T_7023 = valid_11_15 ? 5'hf : _T_7022; // @[Mux.scala 31:69:@1903.4]
  assign _T_7024 = valid_11_14 ? 5'he : _T_7023; // @[Mux.scala 31:69:@1904.4]
  assign _T_7025 = valid_11_13 ? 5'hd : _T_7024; // @[Mux.scala 31:69:@1905.4]
  assign _T_7026 = valid_11_12 ? 5'hc : _T_7025; // @[Mux.scala 31:69:@1906.4]
  assign _T_7027 = valid_11_11 ? 5'hb : _T_7026; // @[Mux.scala 31:69:@1907.4]
  assign _T_7028 = valid_11_10 ? 5'ha : _T_7027; // @[Mux.scala 31:69:@1908.4]
  assign _T_7029 = valid_11_9 ? 5'h9 : _T_7028; // @[Mux.scala 31:69:@1909.4]
  assign _T_7030 = valid_11_8 ? 5'h8 : _T_7029; // @[Mux.scala 31:69:@1910.4]
  assign _T_7031 = valid_11_7 ? 5'h7 : _T_7030; // @[Mux.scala 31:69:@1911.4]
  assign _T_7032 = valid_11_6 ? 5'h6 : _T_7031; // @[Mux.scala 31:69:@1912.4]
  assign _T_7033 = valid_11_5 ? 5'h5 : _T_7032; // @[Mux.scala 31:69:@1913.4]
  assign _T_7034 = valid_11_4 ? 5'h4 : _T_7033; // @[Mux.scala 31:69:@1914.4]
  assign _T_7035 = valid_11_3 ? 5'h3 : _T_7034; // @[Mux.scala 31:69:@1915.4]
  assign _T_7036 = valid_11_2 ? 5'h2 : _T_7035; // @[Mux.scala 31:69:@1916.4]
  assign _T_7037 = valid_11_1 ? 5'h1 : _T_7036; // @[Mux.scala 31:69:@1917.4]
  assign select_11 = valid_11_0 ? 5'h0 : _T_7037; // @[Mux.scala 31:69:@1918.4]
  assign _GEN_353 = 5'h1 == select_11 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@1920.4]
  assign _GEN_354 = 5'h2 == select_11 ? io_inData_2 : _GEN_353; // @[Switch.scala 33:19:@1920.4]
  assign _GEN_355 = 5'h3 == select_11 ? io_inData_3 : _GEN_354; // @[Switch.scala 33:19:@1920.4]
  assign _GEN_356 = 5'h4 == select_11 ? io_inData_4 : _GEN_355; // @[Switch.scala 33:19:@1920.4]
  assign _GEN_357 = 5'h5 == select_11 ? io_inData_5 : _GEN_356; // @[Switch.scala 33:19:@1920.4]
  assign _GEN_358 = 5'h6 == select_11 ? io_inData_6 : _GEN_357; // @[Switch.scala 33:19:@1920.4]
  assign _GEN_359 = 5'h7 == select_11 ? io_inData_7 : _GEN_358; // @[Switch.scala 33:19:@1920.4]
  assign _GEN_360 = 5'h8 == select_11 ? io_inData_8 : _GEN_359; // @[Switch.scala 33:19:@1920.4]
  assign _GEN_361 = 5'h9 == select_11 ? io_inData_9 : _GEN_360; // @[Switch.scala 33:19:@1920.4]
  assign _GEN_362 = 5'ha == select_11 ? io_inData_10 : _GEN_361; // @[Switch.scala 33:19:@1920.4]
  assign _GEN_363 = 5'hb == select_11 ? io_inData_11 : _GEN_362; // @[Switch.scala 33:19:@1920.4]
  assign _GEN_364 = 5'hc == select_11 ? io_inData_12 : _GEN_363; // @[Switch.scala 33:19:@1920.4]
  assign _GEN_365 = 5'hd == select_11 ? io_inData_13 : _GEN_364; // @[Switch.scala 33:19:@1920.4]
  assign _GEN_366 = 5'he == select_11 ? io_inData_14 : _GEN_365; // @[Switch.scala 33:19:@1920.4]
  assign _GEN_367 = 5'hf == select_11 ? io_inData_15 : _GEN_366; // @[Switch.scala 33:19:@1920.4]
  assign _GEN_368 = 5'h10 == select_11 ? io_inData_16 : _GEN_367; // @[Switch.scala 33:19:@1920.4]
  assign _GEN_369 = 5'h11 == select_11 ? io_inData_17 : _GEN_368; // @[Switch.scala 33:19:@1920.4]
  assign _GEN_370 = 5'h12 == select_11 ? io_inData_18 : _GEN_369; // @[Switch.scala 33:19:@1920.4]
  assign _GEN_371 = 5'h13 == select_11 ? io_inData_19 : _GEN_370; // @[Switch.scala 33:19:@1920.4]
  assign _GEN_372 = 5'h14 == select_11 ? io_inData_20 : _GEN_371; // @[Switch.scala 33:19:@1920.4]
  assign _GEN_373 = 5'h15 == select_11 ? io_inData_21 : _GEN_372; // @[Switch.scala 33:19:@1920.4]
  assign _GEN_374 = 5'h16 == select_11 ? io_inData_22 : _GEN_373; // @[Switch.scala 33:19:@1920.4]
  assign _GEN_375 = 5'h17 == select_11 ? io_inData_23 : _GEN_374; // @[Switch.scala 33:19:@1920.4]
  assign _GEN_376 = 5'h18 == select_11 ? io_inData_24 : _GEN_375; // @[Switch.scala 33:19:@1920.4]
  assign _GEN_377 = 5'h19 == select_11 ? io_inData_25 : _GEN_376; // @[Switch.scala 33:19:@1920.4]
  assign _GEN_378 = 5'h1a == select_11 ? io_inData_26 : _GEN_377; // @[Switch.scala 33:19:@1920.4]
  assign _GEN_379 = 5'h1b == select_11 ? io_inData_27 : _GEN_378; // @[Switch.scala 33:19:@1920.4]
  assign _GEN_380 = 5'h1c == select_11 ? io_inData_28 : _GEN_379; // @[Switch.scala 33:19:@1920.4]
  assign _GEN_381 = 5'h1d == select_11 ? io_inData_29 : _GEN_380; // @[Switch.scala 33:19:@1920.4]
  assign _GEN_382 = 5'h1e == select_11 ? io_inData_30 : _GEN_381; // @[Switch.scala 33:19:@1920.4]
  assign _T_7046 = {valid_11_7,valid_11_6,valid_11_5,valid_11_4,valid_11_3,valid_11_2,valid_11_1,valid_11_0}; // @[Switch.scala 34:32:@1927.4]
  assign _T_7054 = {valid_11_15,valid_11_14,valid_11_13,valid_11_12,valid_11_11,valid_11_10,valid_11_9,valid_11_8,_T_7046}; // @[Switch.scala 34:32:@1935.4]
  assign _T_7061 = {valid_11_23,valid_11_22,valid_11_21,valid_11_20,valid_11_19,valid_11_18,valid_11_17,valid_11_16}; // @[Switch.scala 34:32:@1942.4]
  assign _T_7070 = {valid_11_31,valid_11_30,valid_11_29,valid_11_28,valid_11_27,valid_11_26,valid_11_25,valid_11_24,_T_7061,_T_7054}; // @[Switch.scala 34:32:@1951.4]
  assign _T_7074 = io_inAddr_0 == 5'hc; // @[Switch.scala 30:53:@1954.4]
  assign valid_12_0 = io_inValid_0 & _T_7074; // @[Switch.scala 30:36:@1955.4]
  assign _T_7077 = io_inAddr_1 == 5'hc; // @[Switch.scala 30:53:@1957.4]
  assign valid_12_1 = io_inValid_1 & _T_7077; // @[Switch.scala 30:36:@1958.4]
  assign _T_7080 = io_inAddr_2 == 5'hc; // @[Switch.scala 30:53:@1960.4]
  assign valid_12_2 = io_inValid_2 & _T_7080; // @[Switch.scala 30:36:@1961.4]
  assign _T_7083 = io_inAddr_3 == 5'hc; // @[Switch.scala 30:53:@1963.4]
  assign valid_12_3 = io_inValid_3 & _T_7083; // @[Switch.scala 30:36:@1964.4]
  assign _T_7086 = io_inAddr_4 == 5'hc; // @[Switch.scala 30:53:@1966.4]
  assign valid_12_4 = io_inValid_4 & _T_7086; // @[Switch.scala 30:36:@1967.4]
  assign _T_7089 = io_inAddr_5 == 5'hc; // @[Switch.scala 30:53:@1969.4]
  assign valid_12_5 = io_inValid_5 & _T_7089; // @[Switch.scala 30:36:@1970.4]
  assign _T_7092 = io_inAddr_6 == 5'hc; // @[Switch.scala 30:53:@1972.4]
  assign valid_12_6 = io_inValid_6 & _T_7092; // @[Switch.scala 30:36:@1973.4]
  assign _T_7095 = io_inAddr_7 == 5'hc; // @[Switch.scala 30:53:@1975.4]
  assign valid_12_7 = io_inValid_7 & _T_7095; // @[Switch.scala 30:36:@1976.4]
  assign _T_7098 = io_inAddr_8 == 5'hc; // @[Switch.scala 30:53:@1978.4]
  assign valid_12_8 = io_inValid_8 & _T_7098; // @[Switch.scala 30:36:@1979.4]
  assign _T_7101 = io_inAddr_9 == 5'hc; // @[Switch.scala 30:53:@1981.4]
  assign valid_12_9 = io_inValid_9 & _T_7101; // @[Switch.scala 30:36:@1982.4]
  assign _T_7104 = io_inAddr_10 == 5'hc; // @[Switch.scala 30:53:@1984.4]
  assign valid_12_10 = io_inValid_10 & _T_7104; // @[Switch.scala 30:36:@1985.4]
  assign _T_7107 = io_inAddr_11 == 5'hc; // @[Switch.scala 30:53:@1987.4]
  assign valid_12_11 = io_inValid_11 & _T_7107; // @[Switch.scala 30:36:@1988.4]
  assign _T_7110 = io_inAddr_12 == 5'hc; // @[Switch.scala 30:53:@1990.4]
  assign valid_12_12 = io_inValid_12 & _T_7110; // @[Switch.scala 30:36:@1991.4]
  assign _T_7113 = io_inAddr_13 == 5'hc; // @[Switch.scala 30:53:@1993.4]
  assign valid_12_13 = io_inValid_13 & _T_7113; // @[Switch.scala 30:36:@1994.4]
  assign _T_7116 = io_inAddr_14 == 5'hc; // @[Switch.scala 30:53:@1996.4]
  assign valid_12_14 = io_inValid_14 & _T_7116; // @[Switch.scala 30:36:@1997.4]
  assign _T_7119 = io_inAddr_15 == 5'hc; // @[Switch.scala 30:53:@1999.4]
  assign valid_12_15 = io_inValid_15 & _T_7119; // @[Switch.scala 30:36:@2000.4]
  assign _T_7122 = io_inAddr_16 == 5'hc; // @[Switch.scala 30:53:@2002.4]
  assign valid_12_16 = io_inValid_16 & _T_7122; // @[Switch.scala 30:36:@2003.4]
  assign _T_7125 = io_inAddr_17 == 5'hc; // @[Switch.scala 30:53:@2005.4]
  assign valid_12_17 = io_inValid_17 & _T_7125; // @[Switch.scala 30:36:@2006.4]
  assign _T_7128 = io_inAddr_18 == 5'hc; // @[Switch.scala 30:53:@2008.4]
  assign valid_12_18 = io_inValid_18 & _T_7128; // @[Switch.scala 30:36:@2009.4]
  assign _T_7131 = io_inAddr_19 == 5'hc; // @[Switch.scala 30:53:@2011.4]
  assign valid_12_19 = io_inValid_19 & _T_7131; // @[Switch.scala 30:36:@2012.4]
  assign _T_7134 = io_inAddr_20 == 5'hc; // @[Switch.scala 30:53:@2014.4]
  assign valid_12_20 = io_inValid_20 & _T_7134; // @[Switch.scala 30:36:@2015.4]
  assign _T_7137 = io_inAddr_21 == 5'hc; // @[Switch.scala 30:53:@2017.4]
  assign valid_12_21 = io_inValid_21 & _T_7137; // @[Switch.scala 30:36:@2018.4]
  assign _T_7140 = io_inAddr_22 == 5'hc; // @[Switch.scala 30:53:@2020.4]
  assign valid_12_22 = io_inValid_22 & _T_7140; // @[Switch.scala 30:36:@2021.4]
  assign _T_7143 = io_inAddr_23 == 5'hc; // @[Switch.scala 30:53:@2023.4]
  assign valid_12_23 = io_inValid_23 & _T_7143; // @[Switch.scala 30:36:@2024.4]
  assign _T_7146 = io_inAddr_24 == 5'hc; // @[Switch.scala 30:53:@2026.4]
  assign valid_12_24 = io_inValid_24 & _T_7146; // @[Switch.scala 30:36:@2027.4]
  assign _T_7149 = io_inAddr_25 == 5'hc; // @[Switch.scala 30:53:@2029.4]
  assign valid_12_25 = io_inValid_25 & _T_7149; // @[Switch.scala 30:36:@2030.4]
  assign _T_7152 = io_inAddr_26 == 5'hc; // @[Switch.scala 30:53:@2032.4]
  assign valid_12_26 = io_inValid_26 & _T_7152; // @[Switch.scala 30:36:@2033.4]
  assign _T_7155 = io_inAddr_27 == 5'hc; // @[Switch.scala 30:53:@2035.4]
  assign valid_12_27 = io_inValid_27 & _T_7155; // @[Switch.scala 30:36:@2036.4]
  assign _T_7158 = io_inAddr_28 == 5'hc; // @[Switch.scala 30:53:@2038.4]
  assign valid_12_28 = io_inValid_28 & _T_7158; // @[Switch.scala 30:36:@2039.4]
  assign _T_7161 = io_inAddr_29 == 5'hc; // @[Switch.scala 30:53:@2041.4]
  assign valid_12_29 = io_inValid_29 & _T_7161; // @[Switch.scala 30:36:@2042.4]
  assign _T_7164 = io_inAddr_30 == 5'hc; // @[Switch.scala 30:53:@2044.4]
  assign valid_12_30 = io_inValid_30 & _T_7164; // @[Switch.scala 30:36:@2045.4]
  assign _T_7167 = io_inAddr_31 == 5'hc; // @[Switch.scala 30:53:@2047.4]
  assign valid_12_31 = io_inValid_31 & _T_7167; // @[Switch.scala 30:36:@2048.4]
  assign _T_7201 = valid_12_30 ? 5'h1e : 5'h1f; // @[Mux.scala 31:69:@2050.4]
  assign _T_7202 = valid_12_29 ? 5'h1d : _T_7201; // @[Mux.scala 31:69:@2051.4]
  assign _T_7203 = valid_12_28 ? 5'h1c : _T_7202; // @[Mux.scala 31:69:@2052.4]
  assign _T_7204 = valid_12_27 ? 5'h1b : _T_7203; // @[Mux.scala 31:69:@2053.4]
  assign _T_7205 = valid_12_26 ? 5'h1a : _T_7204; // @[Mux.scala 31:69:@2054.4]
  assign _T_7206 = valid_12_25 ? 5'h19 : _T_7205; // @[Mux.scala 31:69:@2055.4]
  assign _T_7207 = valid_12_24 ? 5'h18 : _T_7206; // @[Mux.scala 31:69:@2056.4]
  assign _T_7208 = valid_12_23 ? 5'h17 : _T_7207; // @[Mux.scala 31:69:@2057.4]
  assign _T_7209 = valid_12_22 ? 5'h16 : _T_7208; // @[Mux.scala 31:69:@2058.4]
  assign _T_7210 = valid_12_21 ? 5'h15 : _T_7209; // @[Mux.scala 31:69:@2059.4]
  assign _T_7211 = valid_12_20 ? 5'h14 : _T_7210; // @[Mux.scala 31:69:@2060.4]
  assign _T_7212 = valid_12_19 ? 5'h13 : _T_7211; // @[Mux.scala 31:69:@2061.4]
  assign _T_7213 = valid_12_18 ? 5'h12 : _T_7212; // @[Mux.scala 31:69:@2062.4]
  assign _T_7214 = valid_12_17 ? 5'h11 : _T_7213; // @[Mux.scala 31:69:@2063.4]
  assign _T_7215 = valid_12_16 ? 5'h10 : _T_7214; // @[Mux.scala 31:69:@2064.4]
  assign _T_7216 = valid_12_15 ? 5'hf : _T_7215; // @[Mux.scala 31:69:@2065.4]
  assign _T_7217 = valid_12_14 ? 5'he : _T_7216; // @[Mux.scala 31:69:@2066.4]
  assign _T_7218 = valid_12_13 ? 5'hd : _T_7217; // @[Mux.scala 31:69:@2067.4]
  assign _T_7219 = valid_12_12 ? 5'hc : _T_7218; // @[Mux.scala 31:69:@2068.4]
  assign _T_7220 = valid_12_11 ? 5'hb : _T_7219; // @[Mux.scala 31:69:@2069.4]
  assign _T_7221 = valid_12_10 ? 5'ha : _T_7220; // @[Mux.scala 31:69:@2070.4]
  assign _T_7222 = valid_12_9 ? 5'h9 : _T_7221; // @[Mux.scala 31:69:@2071.4]
  assign _T_7223 = valid_12_8 ? 5'h8 : _T_7222; // @[Mux.scala 31:69:@2072.4]
  assign _T_7224 = valid_12_7 ? 5'h7 : _T_7223; // @[Mux.scala 31:69:@2073.4]
  assign _T_7225 = valid_12_6 ? 5'h6 : _T_7224; // @[Mux.scala 31:69:@2074.4]
  assign _T_7226 = valid_12_5 ? 5'h5 : _T_7225; // @[Mux.scala 31:69:@2075.4]
  assign _T_7227 = valid_12_4 ? 5'h4 : _T_7226; // @[Mux.scala 31:69:@2076.4]
  assign _T_7228 = valid_12_3 ? 5'h3 : _T_7227; // @[Mux.scala 31:69:@2077.4]
  assign _T_7229 = valid_12_2 ? 5'h2 : _T_7228; // @[Mux.scala 31:69:@2078.4]
  assign _T_7230 = valid_12_1 ? 5'h1 : _T_7229; // @[Mux.scala 31:69:@2079.4]
  assign select_12 = valid_12_0 ? 5'h0 : _T_7230; // @[Mux.scala 31:69:@2080.4]
  assign _GEN_385 = 5'h1 == select_12 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@2082.4]
  assign _GEN_386 = 5'h2 == select_12 ? io_inData_2 : _GEN_385; // @[Switch.scala 33:19:@2082.4]
  assign _GEN_387 = 5'h3 == select_12 ? io_inData_3 : _GEN_386; // @[Switch.scala 33:19:@2082.4]
  assign _GEN_388 = 5'h4 == select_12 ? io_inData_4 : _GEN_387; // @[Switch.scala 33:19:@2082.4]
  assign _GEN_389 = 5'h5 == select_12 ? io_inData_5 : _GEN_388; // @[Switch.scala 33:19:@2082.4]
  assign _GEN_390 = 5'h6 == select_12 ? io_inData_6 : _GEN_389; // @[Switch.scala 33:19:@2082.4]
  assign _GEN_391 = 5'h7 == select_12 ? io_inData_7 : _GEN_390; // @[Switch.scala 33:19:@2082.4]
  assign _GEN_392 = 5'h8 == select_12 ? io_inData_8 : _GEN_391; // @[Switch.scala 33:19:@2082.4]
  assign _GEN_393 = 5'h9 == select_12 ? io_inData_9 : _GEN_392; // @[Switch.scala 33:19:@2082.4]
  assign _GEN_394 = 5'ha == select_12 ? io_inData_10 : _GEN_393; // @[Switch.scala 33:19:@2082.4]
  assign _GEN_395 = 5'hb == select_12 ? io_inData_11 : _GEN_394; // @[Switch.scala 33:19:@2082.4]
  assign _GEN_396 = 5'hc == select_12 ? io_inData_12 : _GEN_395; // @[Switch.scala 33:19:@2082.4]
  assign _GEN_397 = 5'hd == select_12 ? io_inData_13 : _GEN_396; // @[Switch.scala 33:19:@2082.4]
  assign _GEN_398 = 5'he == select_12 ? io_inData_14 : _GEN_397; // @[Switch.scala 33:19:@2082.4]
  assign _GEN_399 = 5'hf == select_12 ? io_inData_15 : _GEN_398; // @[Switch.scala 33:19:@2082.4]
  assign _GEN_400 = 5'h10 == select_12 ? io_inData_16 : _GEN_399; // @[Switch.scala 33:19:@2082.4]
  assign _GEN_401 = 5'h11 == select_12 ? io_inData_17 : _GEN_400; // @[Switch.scala 33:19:@2082.4]
  assign _GEN_402 = 5'h12 == select_12 ? io_inData_18 : _GEN_401; // @[Switch.scala 33:19:@2082.4]
  assign _GEN_403 = 5'h13 == select_12 ? io_inData_19 : _GEN_402; // @[Switch.scala 33:19:@2082.4]
  assign _GEN_404 = 5'h14 == select_12 ? io_inData_20 : _GEN_403; // @[Switch.scala 33:19:@2082.4]
  assign _GEN_405 = 5'h15 == select_12 ? io_inData_21 : _GEN_404; // @[Switch.scala 33:19:@2082.4]
  assign _GEN_406 = 5'h16 == select_12 ? io_inData_22 : _GEN_405; // @[Switch.scala 33:19:@2082.4]
  assign _GEN_407 = 5'h17 == select_12 ? io_inData_23 : _GEN_406; // @[Switch.scala 33:19:@2082.4]
  assign _GEN_408 = 5'h18 == select_12 ? io_inData_24 : _GEN_407; // @[Switch.scala 33:19:@2082.4]
  assign _GEN_409 = 5'h19 == select_12 ? io_inData_25 : _GEN_408; // @[Switch.scala 33:19:@2082.4]
  assign _GEN_410 = 5'h1a == select_12 ? io_inData_26 : _GEN_409; // @[Switch.scala 33:19:@2082.4]
  assign _GEN_411 = 5'h1b == select_12 ? io_inData_27 : _GEN_410; // @[Switch.scala 33:19:@2082.4]
  assign _GEN_412 = 5'h1c == select_12 ? io_inData_28 : _GEN_411; // @[Switch.scala 33:19:@2082.4]
  assign _GEN_413 = 5'h1d == select_12 ? io_inData_29 : _GEN_412; // @[Switch.scala 33:19:@2082.4]
  assign _GEN_414 = 5'h1e == select_12 ? io_inData_30 : _GEN_413; // @[Switch.scala 33:19:@2082.4]
  assign _T_7239 = {valid_12_7,valid_12_6,valid_12_5,valid_12_4,valid_12_3,valid_12_2,valid_12_1,valid_12_0}; // @[Switch.scala 34:32:@2089.4]
  assign _T_7247 = {valid_12_15,valid_12_14,valid_12_13,valid_12_12,valid_12_11,valid_12_10,valid_12_9,valid_12_8,_T_7239}; // @[Switch.scala 34:32:@2097.4]
  assign _T_7254 = {valid_12_23,valid_12_22,valid_12_21,valid_12_20,valid_12_19,valid_12_18,valid_12_17,valid_12_16}; // @[Switch.scala 34:32:@2104.4]
  assign _T_7263 = {valid_12_31,valid_12_30,valid_12_29,valid_12_28,valid_12_27,valid_12_26,valid_12_25,valid_12_24,_T_7254,_T_7247}; // @[Switch.scala 34:32:@2113.4]
  assign _T_7267 = io_inAddr_0 == 5'hd; // @[Switch.scala 30:53:@2116.4]
  assign valid_13_0 = io_inValid_0 & _T_7267; // @[Switch.scala 30:36:@2117.4]
  assign _T_7270 = io_inAddr_1 == 5'hd; // @[Switch.scala 30:53:@2119.4]
  assign valid_13_1 = io_inValid_1 & _T_7270; // @[Switch.scala 30:36:@2120.4]
  assign _T_7273 = io_inAddr_2 == 5'hd; // @[Switch.scala 30:53:@2122.4]
  assign valid_13_2 = io_inValid_2 & _T_7273; // @[Switch.scala 30:36:@2123.4]
  assign _T_7276 = io_inAddr_3 == 5'hd; // @[Switch.scala 30:53:@2125.4]
  assign valid_13_3 = io_inValid_3 & _T_7276; // @[Switch.scala 30:36:@2126.4]
  assign _T_7279 = io_inAddr_4 == 5'hd; // @[Switch.scala 30:53:@2128.4]
  assign valid_13_4 = io_inValid_4 & _T_7279; // @[Switch.scala 30:36:@2129.4]
  assign _T_7282 = io_inAddr_5 == 5'hd; // @[Switch.scala 30:53:@2131.4]
  assign valid_13_5 = io_inValid_5 & _T_7282; // @[Switch.scala 30:36:@2132.4]
  assign _T_7285 = io_inAddr_6 == 5'hd; // @[Switch.scala 30:53:@2134.4]
  assign valid_13_6 = io_inValid_6 & _T_7285; // @[Switch.scala 30:36:@2135.4]
  assign _T_7288 = io_inAddr_7 == 5'hd; // @[Switch.scala 30:53:@2137.4]
  assign valid_13_7 = io_inValid_7 & _T_7288; // @[Switch.scala 30:36:@2138.4]
  assign _T_7291 = io_inAddr_8 == 5'hd; // @[Switch.scala 30:53:@2140.4]
  assign valid_13_8 = io_inValid_8 & _T_7291; // @[Switch.scala 30:36:@2141.4]
  assign _T_7294 = io_inAddr_9 == 5'hd; // @[Switch.scala 30:53:@2143.4]
  assign valid_13_9 = io_inValid_9 & _T_7294; // @[Switch.scala 30:36:@2144.4]
  assign _T_7297 = io_inAddr_10 == 5'hd; // @[Switch.scala 30:53:@2146.4]
  assign valid_13_10 = io_inValid_10 & _T_7297; // @[Switch.scala 30:36:@2147.4]
  assign _T_7300 = io_inAddr_11 == 5'hd; // @[Switch.scala 30:53:@2149.4]
  assign valid_13_11 = io_inValid_11 & _T_7300; // @[Switch.scala 30:36:@2150.4]
  assign _T_7303 = io_inAddr_12 == 5'hd; // @[Switch.scala 30:53:@2152.4]
  assign valid_13_12 = io_inValid_12 & _T_7303; // @[Switch.scala 30:36:@2153.4]
  assign _T_7306 = io_inAddr_13 == 5'hd; // @[Switch.scala 30:53:@2155.4]
  assign valid_13_13 = io_inValid_13 & _T_7306; // @[Switch.scala 30:36:@2156.4]
  assign _T_7309 = io_inAddr_14 == 5'hd; // @[Switch.scala 30:53:@2158.4]
  assign valid_13_14 = io_inValid_14 & _T_7309; // @[Switch.scala 30:36:@2159.4]
  assign _T_7312 = io_inAddr_15 == 5'hd; // @[Switch.scala 30:53:@2161.4]
  assign valid_13_15 = io_inValid_15 & _T_7312; // @[Switch.scala 30:36:@2162.4]
  assign _T_7315 = io_inAddr_16 == 5'hd; // @[Switch.scala 30:53:@2164.4]
  assign valid_13_16 = io_inValid_16 & _T_7315; // @[Switch.scala 30:36:@2165.4]
  assign _T_7318 = io_inAddr_17 == 5'hd; // @[Switch.scala 30:53:@2167.4]
  assign valid_13_17 = io_inValid_17 & _T_7318; // @[Switch.scala 30:36:@2168.4]
  assign _T_7321 = io_inAddr_18 == 5'hd; // @[Switch.scala 30:53:@2170.4]
  assign valid_13_18 = io_inValid_18 & _T_7321; // @[Switch.scala 30:36:@2171.4]
  assign _T_7324 = io_inAddr_19 == 5'hd; // @[Switch.scala 30:53:@2173.4]
  assign valid_13_19 = io_inValid_19 & _T_7324; // @[Switch.scala 30:36:@2174.4]
  assign _T_7327 = io_inAddr_20 == 5'hd; // @[Switch.scala 30:53:@2176.4]
  assign valid_13_20 = io_inValid_20 & _T_7327; // @[Switch.scala 30:36:@2177.4]
  assign _T_7330 = io_inAddr_21 == 5'hd; // @[Switch.scala 30:53:@2179.4]
  assign valid_13_21 = io_inValid_21 & _T_7330; // @[Switch.scala 30:36:@2180.4]
  assign _T_7333 = io_inAddr_22 == 5'hd; // @[Switch.scala 30:53:@2182.4]
  assign valid_13_22 = io_inValid_22 & _T_7333; // @[Switch.scala 30:36:@2183.4]
  assign _T_7336 = io_inAddr_23 == 5'hd; // @[Switch.scala 30:53:@2185.4]
  assign valid_13_23 = io_inValid_23 & _T_7336; // @[Switch.scala 30:36:@2186.4]
  assign _T_7339 = io_inAddr_24 == 5'hd; // @[Switch.scala 30:53:@2188.4]
  assign valid_13_24 = io_inValid_24 & _T_7339; // @[Switch.scala 30:36:@2189.4]
  assign _T_7342 = io_inAddr_25 == 5'hd; // @[Switch.scala 30:53:@2191.4]
  assign valid_13_25 = io_inValid_25 & _T_7342; // @[Switch.scala 30:36:@2192.4]
  assign _T_7345 = io_inAddr_26 == 5'hd; // @[Switch.scala 30:53:@2194.4]
  assign valid_13_26 = io_inValid_26 & _T_7345; // @[Switch.scala 30:36:@2195.4]
  assign _T_7348 = io_inAddr_27 == 5'hd; // @[Switch.scala 30:53:@2197.4]
  assign valid_13_27 = io_inValid_27 & _T_7348; // @[Switch.scala 30:36:@2198.4]
  assign _T_7351 = io_inAddr_28 == 5'hd; // @[Switch.scala 30:53:@2200.4]
  assign valid_13_28 = io_inValid_28 & _T_7351; // @[Switch.scala 30:36:@2201.4]
  assign _T_7354 = io_inAddr_29 == 5'hd; // @[Switch.scala 30:53:@2203.4]
  assign valid_13_29 = io_inValid_29 & _T_7354; // @[Switch.scala 30:36:@2204.4]
  assign _T_7357 = io_inAddr_30 == 5'hd; // @[Switch.scala 30:53:@2206.4]
  assign valid_13_30 = io_inValid_30 & _T_7357; // @[Switch.scala 30:36:@2207.4]
  assign _T_7360 = io_inAddr_31 == 5'hd; // @[Switch.scala 30:53:@2209.4]
  assign valid_13_31 = io_inValid_31 & _T_7360; // @[Switch.scala 30:36:@2210.4]
  assign _T_7394 = valid_13_30 ? 5'h1e : 5'h1f; // @[Mux.scala 31:69:@2212.4]
  assign _T_7395 = valid_13_29 ? 5'h1d : _T_7394; // @[Mux.scala 31:69:@2213.4]
  assign _T_7396 = valid_13_28 ? 5'h1c : _T_7395; // @[Mux.scala 31:69:@2214.4]
  assign _T_7397 = valid_13_27 ? 5'h1b : _T_7396; // @[Mux.scala 31:69:@2215.4]
  assign _T_7398 = valid_13_26 ? 5'h1a : _T_7397; // @[Mux.scala 31:69:@2216.4]
  assign _T_7399 = valid_13_25 ? 5'h19 : _T_7398; // @[Mux.scala 31:69:@2217.4]
  assign _T_7400 = valid_13_24 ? 5'h18 : _T_7399; // @[Mux.scala 31:69:@2218.4]
  assign _T_7401 = valid_13_23 ? 5'h17 : _T_7400; // @[Mux.scala 31:69:@2219.4]
  assign _T_7402 = valid_13_22 ? 5'h16 : _T_7401; // @[Mux.scala 31:69:@2220.4]
  assign _T_7403 = valid_13_21 ? 5'h15 : _T_7402; // @[Mux.scala 31:69:@2221.4]
  assign _T_7404 = valid_13_20 ? 5'h14 : _T_7403; // @[Mux.scala 31:69:@2222.4]
  assign _T_7405 = valid_13_19 ? 5'h13 : _T_7404; // @[Mux.scala 31:69:@2223.4]
  assign _T_7406 = valid_13_18 ? 5'h12 : _T_7405; // @[Mux.scala 31:69:@2224.4]
  assign _T_7407 = valid_13_17 ? 5'h11 : _T_7406; // @[Mux.scala 31:69:@2225.4]
  assign _T_7408 = valid_13_16 ? 5'h10 : _T_7407; // @[Mux.scala 31:69:@2226.4]
  assign _T_7409 = valid_13_15 ? 5'hf : _T_7408; // @[Mux.scala 31:69:@2227.4]
  assign _T_7410 = valid_13_14 ? 5'he : _T_7409; // @[Mux.scala 31:69:@2228.4]
  assign _T_7411 = valid_13_13 ? 5'hd : _T_7410; // @[Mux.scala 31:69:@2229.4]
  assign _T_7412 = valid_13_12 ? 5'hc : _T_7411; // @[Mux.scala 31:69:@2230.4]
  assign _T_7413 = valid_13_11 ? 5'hb : _T_7412; // @[Mux.scala 31:69:@2231.4]
  assign _T_7414 = valid_13_10 ? 5'ha : _T_7413; // @[Mux.scala 31:69:@2232.4]
  assign _T_7415 = valid_13_9 ? 5'h9 : _T_7414; // @[Mux.scala 31:69:@2233.4]
  assign _T_7416 = valid_13_8 ? 5'h8 : _T_7415; // @[Mux.scala 31:69:@2234.4]
  assign _T_7417 = valid_13_7 ? 5'h7 : _T_7416; // @[Mux.scala 31:69:@2235.4]
  assign _T_7418 = valid_13_6 ? 5'h6 : _T_7417; // @[Mux.scala 31:69:@2236.4]
  assign _T_7419 = valid_13_5 ? 5'h5 : _T_7418; // @[Mux.scala 31:69:@2237.4]
  assign _T_7420 = valid_13_4 ? 5'h4 : _T_7419; // @[Mux.scala 31:69:@2238.4]
  assign _T_7421 = valid_13_3 ? 5'h3 : _T_7420; // @[Mux.scala 31:69:@2239.4]
  assign _T_7422 = valid_13_2 ? 5'h2 : _T_7421; // @[Mux.scala 31:69:@2240.4]
  assign _T_7423 = valid_13_1 ? 5'h1 : _T_7422; // @[Mux.scala 31:69:@2241.4]
  assign select_13 = valid_13_0 ? 5'h0 : _T_7423; // @[Mux.scala 31:69:@2242.4]
  assign _GEN_417 = 5'h1 == select_13 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@2244.4]
  assign _GEN_418 = 5'h2 == select_13 ? io_inData_2 : _GEN_417; // @[Switch.scala 33:19:@2244.4]
  assign _GEN_419 = 5'h3 == select_13 ? io_inData_3 : _GEN_418; // @[Switch.scala 33:19:@2244.4]
  assign _GEN_420 = 5'h4 == select_13 ? io_inData_4 : _GEN_419; // @[Switch.scala 33:19:@2244.4]
  assign _GEN_421 = 5'h5 == select_13 ? io_inData_5 : _GEN_420; // @[Switch.scala 33:19:@2244.4]
  assign _GEN_422 = 5'h6 == select_13 ? io_inData_6 : _GEN_421; // @[Switch.scala 33:19:@2244.4]
  assign _GEN_423 = 5'h7 == select_13 ? io_inData_7 : _GEN_422; // @[Switch.scala 33:19:@2244.4]
  assign _GEN_424 = 5'h8 == select_13 ? io_inData_8 : _GEN_423; // @[Switch.scala 33:19:@2244.4]
  assign _GEN_425 = 5'h9 == select_13 ? io_inData_9 : _GEN_424; // @[Switch.scala 33:19:@2244.4]
  assign _GEN_426 = 5'ha == select_13 ? io_inData_10 : _GEN_425; // @[Switch.scala 33:19:@2244.4]
  assign _GEN_427 = 5'hb == select_13 ? io_inData_11 : _GEN_426; // @[Switch.scala 33:19:@2244.4]
  assign _GEN_428 = 5'hc == select_13 ? io_inData_12 : _GEN_427; // @[Switch.scala 33:19:@2244.4]
  assign _GEN_429 = 5'hd == select_13 ? io_inData_13 : _GEN_428; // @[Switch.scala 33:19:@2244.4]
  assign _GEN_430 = 5'he == select_13 ? io_inData_14 : _GEN_429; // @[Switch.scala 33:19:@2244.4]
  assign _GEN_431 = 5'hf == select_13 ? io_inData_15 : _GEN_430; // @[Switch.scala 33:19:@2244.4]
  assign _GEN_432 = 5'h10 == select_13 ? io_inData_16 : _GEN_431; // @[Switch.scala 33:19:@2244.4]
  assign _GEN_433 = 5'h11 == select_13 ? io_inData_17 : _GEN_432; // @[Switch.scala 33:19:@2244.4]
  assign _GEN_434 = 5'h12 == select_13 ? io_inData_18 : _GEN_433; // @[Switch.scala 33:19:@2244.4]
  assign _GEN_435 = 5'h13 == select_13 ? io_inData_19 : _GEN_434; // @[Switch.scala 33:19:@2244.4]
  assign _GEN_436 = 5'h14 == select_13 ? io_inData_20 : _GEN_435; // @[Switch.scala 33:19:@2244.4]
  assign _GEN_437 = 5'h15 == select_13 ? io_inData_21 : _GEN_436; // @[Switch.scala 33:19:@2244.4]
  assign _GEN_438 = 5'h16 == select_13 ? io_inData_22 : _GEN_437; // @[Switch.scala 33:19:@2244.4]
  assign _GEN_439 = 5'h17 == select_13 ? io_inData_23 : _GEN_438; // @[Switch.scala 33:19:@2244.4]
  assign _GEN_440 = 5'h18 == select_13 ? io_inData_24 : _GEN_439; // @[Switch.scala 33:19:@2244.4]
  assign _GEN_441 = 5'h19 == select_13 ? io_inData_25 : _GEN_440; // @[Switch.scala 33:19:@2244.4]
  assign _GEN_442 = 5'h1a == select_13 ? io_inData_26 : _GEN_441; // @[Switch.scala 33:19:@2244.4]
  assign _GEN_443 = 5'h1b == select_13 ? io_inData_27 : _GEN_442; // @[Switch.scala 33:19:@2244.4]
  assign _GEN_444 = 5'h1c == select_13 ? io_inData_28 : _GEN_443; // @[Switch.scala 33:19:@2244.4]
  assign _GEN_445 = 5'h1d == select_13 ? io_inData_29 : _GEN_444; // @[Switch.scala 33:19:@2244.4]
  assign _GEN_446 = 5'h1e == select_13 ? io_inData_30 : _GEN_445; // @[Switch.scala 33:19:@2244.4]
  assign _T_7432 = {valid_13_7,valid_13_6,valid_13_5,valid_13_4,valid_13_3,valid_13_2,valid_13_1,valid_13_0}; // @[Switch.scala 34:32:@2251.4]
  assign _T_7440 = {valid_13_15,valid_13_14,valid_13_13,valid_13_12,valid_13_11,valid_13_10,valid_13_9,valid_13_8,_T_7432}; // @[Switch.scala 34:32:@2259.4]
  assign _T_7447 = {valid_13_23,valid_13_22,valid_13_21,valid_13_20,valid_13_19,valid_13_18,valid_13_17,valid_13_16}; // @[Switch.scala 34:32:@2266.4]
  assign _T_7456 = {valid_13_31,valid_13_30,valid_13_29,valid_13_28,valid_13_27,valid_13_26,valid_13_25,valid_13_24,_T_7447,_T_7440}; // @[Switch.scala 34:32:@2275.4]
  assign _T_7460 = io_inAddr_0 == 5'he; // @[Switch.scala 30:53:@2278.4]
  assign valid_14_0 = io_inValid_0 & _T_7460; // @[Switch.scala 30:36:@2279.4]
  assign _T_7463 = io_inAddr_1 == 5'he; // @[Switch.scala 30:53:@2281.4]
  assign valid_14_1 = io_inValid_1 & _T_7463; // @[Switch.scala 30:36:@2282.4]
  assign _T_7466 = io_inAddr_2 == 5'he; // @[Switch.scala 30:53:@2284.4]
  assign valid_14_2 = io_inValid_2 & _T_7466; // @[Switch.scala 30:36:@2285.4]
  assign _T_7469 = io_inAddr_3 == 5'he; // @[Switch.scala 30:53:@2287.4]
  assign valid_14_3 = io_inValid_3 & _T_7469; // @[Switch.scala 30:36:@2288.4]
  assign _T_7472 = io_inAddr_4 == 5'he; // @[Switch.scala 30:53:@2290.4]
  assign valid_14_4 = io_inValid_4 & _T_7472; // @[Switch.scala 30:36:@2291.4]
  assign _T_7475 = io_inAddr_5 == 5'he; // @[Switch.scala 30:53:@2293.4]
  assign valid_14_5 = io_inValid_5 & _T_7475; // @[Switch.scala 30:36:@2294.4]
  assign _T_7478 = io_inAddr_6 == 5'he; // @[Switch.scala 30:53:@2296.4]
  assign valid_14_6 = io_inValid_6 & _T_7478; // @[Switch.scala 30:36:@2297.4]
  assign _T_7481 = io_inAddr_7 == 5'he; // @[Switch.scala 30:53:@2299.4]
  assign valid_14_7 = io_inValid_7 & _T_7481; // @[Switch.scala 30:36:@2300.4]
  assign _T_7484 = io_inAddr_8 == 5'he; // @[Switch.scala 30:53:@2302.4]
  assign valid_14_8 = io_inValid_8 & _T_7484; // @[Switch.scala 30:36:@2303.4]
  assign _T_7487 = io_inAddr_9 == 5'he; // @[Switch.scala 30:53:@2305.4]
  assign valid_14_9 = io_inValid_9 & _T_7487; // @[Switch.scala 30:36:@2306.4]
  assign _T_7490 = io_inAddr_10 == 5'he; // @[Switch.scala 30:53:@2308.4]
  assign valid_14_10 = io_inValid_10 & _T_7490; // @[Switch.scala 30:36:@2309.4]
  assign _T_7493 = io_inAddr_11 == 5'he; // @[Switch.scala 30:53:@2311.4]
  assign valid_14_11 = io_inValid_11 & _T_7493; // @[Switch.scala 30:36:@2312.4]
  assign _T_7496 = io_inAddr_12 == 5'he; // @[Switch.scala 30:53:@2314.4]
  assign valid_14_12 = io_inValid_12 & _T_7496; // @[Switch.scala 30:36:@2315.4]
  assign _T_7499 = io_inAddr_13 == 5'he; // @[Switch.scala 30:53:@2317.4]
  assign valid_14_13 = io_inValid_13 & _T_7499; // @[Switch.scala 30:36:@2318.4]
  assign _T_7502 = io_inAddr_14 == 5'he; // @[Switch.scala 30:53:@2320.4]
  assign valid_14_14 = io_inValid_14 & _T_7502; // @[Switch.scala 30:36:@2321.4]
  assign _T_7505 = io_inAddr_15 == 5'he; // @[Switch.scala 30:53:@2323.4]
  assign valid_14_15 = io_inValid_15 & _T_7505; // @[Switch.scala 30:36:@2324.4]
  assign _T_7508 = io_inAddr_16 == 5'he; // @[Switch.scala 30:53:@2326.4]
  assign valid_14_16 = io_inValid_16 & _T_7508; // @[Switch.scala 30:36:@2327.4]
  assign _T_7511 = io_inAddr_17 == 5'he; // @[Switch.scala 30:53:@2329.4]
  assign valid_14_17 = io_inValid_17 & _T_7511; // @[Switch.scala 30:36:@2330.4]
  assign _T_7514 = io_inAddr_18 == 5'he; // @[Switch.scala 30:53:@2332.4]
  assign valid_14_18 = io_inValid_18 & _T_7514; // @[Switch.scala 30:36:@2333.4]
  assign _T_7517 = io_inAddr_19 == 5'he; // @[Switch.scala 30:53:@2335.4]
  assign valid_14_19 = io_inValid_19 & _T_7517; // @[Switch.scala 30:36:@2336.4]
  assign _T_7520 = io_inAddr_20 == 5'he; // @[Switch.scala 30:53:@2338.4]
  assign valid_14_20 = io_inValid_20 & _T_7520; // @[Switch.scala 30:36:@2339.4]
  assign _T_7523 = io_inAddr_21 == 5'he; // @[Switch.scala 30:53:@2341.4]
  assign valid_14_21 = io_inValid_21 & _T_7523; // @[Switch.scala 30:36:@2342.4]
  assign _T_7526 = io_inAddr_22 == 5'he; // @[Switch.scala 30:53:@2344.4]
  assign valid_14_22 = io_inValid_22 & _T_7526; // @[Switch.scala 30:36:@2345.4]
  assign _T_7529 = io_inAddr_23 == 5'he; // @[Switch.scala 30:53:@2347.4]
  assign valid_14_23 = io_inValid_23 & _T_7529; // @[Switch.scala 30:36:@2348.4]
  assign _T_7532 = io_inAddr_24 == 5'he; // @[Switch.scala 30:53:@2350.4]
  assign valid_14_24 = io_inValid_24 & _T_7532; // @[Switch.scala 30:36:@2351.4]
  assign _T_7535 = io_inAddr_25 == 5'he; // @[Switch.scala 30:53:@2353.4]
  assign valid_14_25 = io_inValid_25 & _T_7535; // @[Switch.scala 30:36:@2354.4]
  assign _T_7538 = io_inAddr_26 == 5'he; // @[Switch.scala 30:53:@2356.4]
  assign valid_14_26 = io_inValid_26 & _T_7538; // @[Switch.scala 30:36:@2357.4]
  assign _T_7541 = io_inAddr_27 == 5'he; // @[Switch.scala 30:53:@2359.4]
  assign valid_14_27 = io_inValid_27 & _T_7541; // @[Switch.scala 30:36:@2360.4]
  assign _T_7544 = io_inAddr_28 == 5'he; // @[Switch.scala 30:53:@2362.4]
  assign valid_14_28 = io_inValid_28 & _T_7544; // @[Switch.scala 30:36:@2363.4]
  assign _T_7547 = io_inAddr_29 == 5'he; // @[Switch.scala 30:53:@2365.4]
  assign valid_14_29 = io_inValid_29 & _T_7547; // @[Switch.scala 30:36:@2366.4]
  assign _T_7550 = io_inAddr_30 == 5'he; // @[Switch.scala 30:53:@2368.4]
  assign valid_14_30 = io_inValid_30 & _T_7550; // @[Switch.scala 30:36:@2369.4]
  assign _T_7553 = io_inAddr_31 == 5'he; // @[Switch.scala 30:53:@2371.4]
  assign valid_14_31 = io_inValid_31 & _T_7553; // @[Switch.scala 30:36:@2372.4]
  assign _T_7587 = valid_14_30 ? 5'h1e : 5'h1f; // @[Mux.scala 31:69:@2374.4]
  assign _T_7588 = valid_14_29 ? 5'h1d : _T_7587; // @[Mux.scala 31:69:@2375.4]
  assign _T_7589 = valid_14_28 ? 5'h1c : _T_7588; // @[Mux.scala 31:69:@2376.4]
  assign _T_7590 = valid_14_27 ? 5'h1b : _T_7589; // @[Mux.scala 31:69:@2377.4]
  assign _T_7591 = valid_14_26 ? 5'h1a : _T_7590; // @[Mux.scala 31:69:@2378.4]
  assign _T_7592 = valid_14_25 ? 5'h19 : _T_7591; // @[Mux.scala 31:69:@2379.4]
  assign _T_7593 = valid_14_24 ? 5'h18 : _T_7592; // @[Mux.scala 31:69:@2380.4]
  assign _T_7594 = valid_14_23 ? 5'h17 : _T_7593; // @[Mux.scala 31:69:@2381.4]
  assign _T_7595 = valid_14_22 ? 5'h16 : _T_7594; // @[Mux.scala 31:69:@2382.4]
  assign _T_7596 = valid_14_21 ? 5'h15 : _T_7595; // @[Mux.scala 31:69:@2383.4]
  assign _T_7597 = valid_14_20 ? 5'h14 : _T_7596; // @[Mux.scala 31:69:@2384.4]
  assign _T_7598 = valid_14_19 ? 5'h13 : _T_7597; // @[Mux.scala 31:69:@2385.4]
  assign _T_7599 = valid_14_18 ? 5'h12 : _T_7598; // @[Mux.scala 31:69:@2386.4]
  assign _T_7600 = valid_14_17 ? 5'h11 : _T_7599; // @[Mux.scala 31:69:@2387.4]
  assign _T_7601 = valid_14_16 ? 5'h10 : _T_7600; // @[Mux.scala 31:69:@2388.4]
  assign _T_7602 = valid_14_15 ? 5'hf : _T_7601; // @[Mux.scala 31:69:@2389.4]
  assign _T_7603 = valid_14_14 ? 5'he : _T_7602; // @[Mux.scala 31:69:@2390.4]
  assign _T_7604 = valid_14_13 ? 5'hd : _T_7603; // @[Mux.scala 31:69:@2391.4]
  assign _T_7605 = valid_14_12 ? 5'hc : _T_7604; // @[Mux.scala 31:69:@2392.4]
  assign _T_7606 = valid_14_11 ? 5'hb : _T_7605; // @[Mux.scala 31:69:@2393.4]
  assign _T_7607 = valid_14_10 ? 5'ha : _T_7606; // @[Mux.scala 31:69:@2394.4]
  assign _T_7608 = valid_14_9 ? 5'h9 : _T_7607; // @[Mux.scala 31:69:@2395.4]
  assign _T_7609 = valid_14_8 ? 5'h8 : _T_7608; // @[Mux.scala 31:69:@2396.4]
  assign _T_7610 = valid_14_7 ? 5'h7 : _T_7609; // @[Mux.scala 31:69:@2397.4]
  assign _T_7611 = valid_14_6 ? 5'h6 : _T_7610; // @[Mux.scala 31:69:@2398.4]
  assign _T_7612 = valid_14_5 ? 5'h5 : _T_7611; // @[Mux.scala 31:69:@2399.4]
  assign _T_7613 = valid_14_4 ? 5'h4 : _T_7612; // @[Mux.scala 31:69:@2400.4]
  assign _T_7614 = valid_14_3 ? 5'h3 : _T_7613; // @[Mux.scala 31:69:@2401.4]
  assign _T_7615 = valid_14_2 ? 5'h2 : _T_7614; // @[Mux.scala 31:69:@2402.4]
  assign _T_7616 = valid_14_1 ? 5'h1 : _T_7615; // @[Mux.scala 31:69:@2403.4]
  assign select_14 = valid_14_0 ? 5'h0 : _T_7616; // @[Mux.scala 31:69:@2404.4]
  assign _GEN_449 = 5'h1 == select_14 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@2406.4]
  assign _GEN_450 = 5'h2 == select_14 ? io_inData_2 : _GEN_449; // @[Switch.scala 33:19:@2406.4]
  assign _GEN_451 = 5'h3 == select_14 ? io_inData_3 : _GEN_450; // @[Switch.scala 33:19:@2406.4]
  assign _GEN_452 = 5'h4 == select_14 ? io_inData_4 : _GEN_451; // @[Switch.scala 33:19:@2406.4]
  assign _GEN_453 = 5'h5 == select_14 ? io_inData_5 : _GEN_452; // @[Switch.scala 33:19:@2406.4]
  assign _GEN_454 = 5'h6 == select_14 ? io_inData_6 : _GEN_453; // @[Switch.scala 33:19:@2406.4]
  assign _GEN_455 = 5'h7 == select_14 ? io_inData_7 : _GEN_454; // @[Switch.scala 33:19:@2406.4]
  assign _GEN_456 = 5'h8 == select_14 ? io_inData_8 : _GEN_455; // @[Switch.scala 33:19:@2406.4]
  assign _GEN_457 = 5'h9 == select_14 ? io_inData_9 : _GEN_456; // @[Switch.scala 33:19:@2406.4]
  assign _GEN_458 = 5'ha == select_14 ? io_inData_10 : _GEN_457; // @[Switch.scala 33:19:@2406.4]
  assign _GEN_459 = 5'hb == select_14 ? io_inData_11 : _GEN_458; // @[Switch.scala 33:19:@2406.4]
  assign _GEN_460 = 5'hc == select_14 ? io_inData_12 : _GEN_459; // @[Switch.scala 33:19:@2406.4]
  assign _GEN_461 = 5'hd == select_14 ? io_inData_13 : _GEN_460; // @[Switch.scala 33:19:@2406.4]
  assign _GEN_462 = 5'he == select_14 ? io_inData_14 : _GEN_461; // @[Switch.scala 33:19:@2406.4]
  assign _GEN_463 = 5'hf == select_14 ? io_inData_15 : _GEN_462; // @[Switch.scala 33:19:@2406.4]
  assign _GEN_464 = 5'h10 == select_14 ? io_inData_16 : _GEN_463; // @[Switch.scala 33:19:@2406.4]
  assign _GEN_465 = 5'h11 == select_14 ? io_inData_17 : _GEN_464; // @[Switch.scala 33:19:@2406.4]
  assign _GEN_466 = 5'h12 == select_14 ? io_inData_18 : _GEN_465; // @[Switch.scala 33:19:@2406.4]
  assign _GEN_467 = 5'h13 == select_14 ? io_inData_19 : _GEN_466; // @[Switch.scala 33:19:@2406.4]
  assign _GEN_468 = 5'h14 == select_14 ? io_inData_20 : _GEN_467; // @[Switch.scala 33:19:@2406.4]
  assign _GEN_469 = 5'h15 == select_14 ? io_inData_21 : _GEN_468; // @[Switch.scala 33:19:@2406.4]
  assign _GEN_470 = 5'h16 == select_14 ? io_inData_22 : _GEN_469; // @[Switch.scala 33:19:@2406.4]
  assign _GEN_471 = 5'h17 == select_14 ? io_inData_23 : _GEN_470; // @[Switch.scala 33:19:@2406.4]
  assign _GEN_472 = 5'h18 == select_14 ? io_inData_24 : _GEN_471; // @[Switch.scala 33:19:@2406.4]
  assign _GEN_473 = 5'h19 == select_14 ? io_inData_25 : _GEN_472; // @[Switch.scala 33:19:@2406.4]
  assign _GEN_474 = 5'h1a == select_14 ? io_inData_26 : _GEN_473; // @[Switch.scala 33:19:@2406.4]
  assign _GEN_475 = 5'h1b == select_14 ? io_inData_27 : _GEN_474; // @[Switch.scala 33:19:@2406.4]
  assign _GEN_476 = 5'h1c == select_14 ? io_inData_28 : _GEN_475; // @[Switch.scala 33:19:@2406.4]
  assign _GEN_477 = 5'h1d == select_14 ? io_inData_29 : _GEN_476; // @[Switch.scala 33:19:@2406.4]
  assign _GEN_478 = 5'h1e == select_14 ? io_inData_30 : _GEN_477; // @[Switch.scala 33:19:@2406.4]
  assign _T_7625 = {valid_14_7,valid_14_6,valid_14_5,valid_14_4,valid_14_3,valid_14_2,valid_14_1,valid_14_0}; // @[Switch.scala 34:32:@2413.4]
  assign _T_7633 = {valid_14_15,valid_14_14,valid_14_13,valid_14_12,valid_14_11,valid_14_10,valid_14_9,valid_14_8,_T_7625}; // @[Switch.scala 34:32:@2421.4]
  assign _T_7640 = {valid_14_23,valid_14_22,valid_14_21,valid_14_20,valid_14_19,valid_14_18,valid_14_17,valid_14_16}; // @[Switch.scala 34:32:@2428.4]
  assign _T_7649 = {valid_14_31,valid_14_30,valid_14_29,valid_14_28,valid_14_27,valid_14_26,valid_14_25,valid_14_24,_T_7640,_T_7633}; // @[Switch.scala 34:32:@2437.4]
  assign _T_7653 = io_inAddr_0 == 5'hf; // @[Switch.scala 30:53:@2440.4]
  assign valid_15_0 = io_inValid_0 & _T_7653; // @[Switch.scala 30:36:@2441.4]
  assign _T_7656 = io_inAddr_1 == 5'hf; // @[Switch.scala 30:53:@2443.4]
  assign valid_15_1 = io_inValid_1 & _T_7656; // @[Switch.scala 30:36:@2444.4]
  assign _T_7659 = io_inAddr_2 == 5'hf; // @[Switch.scala 30:53:@2446.4]
  assign valid_15_2 = io_inValid_2 & _T_7659; // @[Switch.scala 30:36:@2447.4]
  assign _T_7662 = io_inAddr_3 == 5'hf; // @[Switch.scala 30:53:@2449.4]
  assign valid_15_3 = io_inValid_3 & _T_7662; // @[Switch.scala 30:36:@2450.4]
  assign _T_7665 = io_inAddr_4 == 5'hf; // @[Switch.scala 30:53:@2452.4]
  assign valid_15_4 = io_inValid_4 & _T_7665; // @[Switch.scala 30:36:@2453.4]
  assign _T_7668 = io_inAddr_5 == 5'hf; // @[Switch.scala 30:53:@2455.4]
  assign valid_15_5 = io_inValid_5 & _T_7668; // @[Switch.scala 30:36:@2456.4]
  assign _T_7671 = io_inAddr_6 == 5'hf; // @[Switch.scala 30:53:@2458.4]
  assign valid_15_6 = io_inValid_6 & _T_7671; // @[Switch.scala 30:36:@2459.4]
  assign _T_7674 = io_inAddr_7 == 5'hf; // @[Switch.scala 30:53:@2461.4]
  assign valid_15_7 = io_inValid_7 & _T_7674; // @[Switch.scala 30:36:@2462.4]
  assign _T_7677 = io_inAddr_8 == 5'hf; // @[Switch.scala 30:53:@2464.4]
  assign valid_15_8 = io_inValid_8 & _T_7677; // @[Switch.scala 30:36:@2465.4]
  assign _T_7680 = io_inAddr_9 == 5'hf; // @[Switch.scala 30:53:@2467.4]
  assign valid_15_9 = io_inValid_9 & _T_7680; // @[Switch.scala 30:36:@2468.4]
  assign _T_7683 = io_inAddr_10 == 5'hf; // @[Switch.scala 30:53:@2470.4]
  assign valid_15_10 = io_inValid_10 & _T_7683; // @[Switch.scala 30:36:@2471.4]
  assign _T_7686 = io_inAddr_11 == 5'hf; // @[Switch.scala 30:53:@2473.4]
  assign valid_15_11 = io_inValid_11 & _T_7686; // @[Switch.scala 30:36:@2474.4]
  assign _T_7689 = io_inAddr_12 == 5'hf; // @[Switch.scala 30:53:@2476.4]
  assign valid_15_12 = io_inValid_12 & _T_7689; // @[Switch.scala 30:36:@2477.4]
  assign _T_7692 = io_inAddr_13 == 5'hf; // @[Switch.scala 30:53:@2479.4]
  assign valid_15_13 = io_inValid_13 & _T_7692; // @[Switch.scala 30:36:@2480.4]
  assign _T_7695 = io_inAddr_14 == 5'hf; // @[Switch.scala 30:53:@2482.4]
  assign valid_15_14 = io_inValid_14 & _T_7695; // @[Switch.scala 30:36:@2483.4]
  assign _T_7698 = io_inAddr_15 == 5'hf; // @[Switch.scala 30:53:@2485.4]
  assign valid_15_15 = io_inValid_15 & _T_7698; // @[Switch.scala 30:36:@2486.4]
  assign _T_7701 = io_inAddr_16 == 5'hf; // @[Switch.scala 30:53:@2488.4]
  assign valid_15_16 = io_inValid_16 & _T_7701; // @[Switch.scala 30:36:@2489.4]
  assign _T_7704 = io_inAddr_17 == 5'hf; // @[Switch.scala 30:53:@2491.4]
  assign valid_15_17 = io_inValid_17 & _T_7704; // @[Switch.scala 30:36:@2492.4]
  assign _T_7707 = io_inAddr_18 == 5'hf; // @[Switch.scala 30:53:@2494.4]
  assign valid_15_18 = io_inValid_18 & _T_7707; // @[Switch.scala 30:36:@2495.4]
  assign _T_7710 = io_inAddr_19 == 5'hf; // @[Switch.scala 30:53:@2497.4]
  assign valid_15_19 = io_inValid_19 & _T_7710; // @[Switch.scala 30:36:@2498.4]
  assign _T_7713 = io_inAddr_20 == 5'hf; // @[Switch.scala 30:53:@2500.4]
  assign valid_15_20 = io_inValid_20 & _T_7713; // @[Switch.scala 30:36:@2501.4]
  assign _T_7716 = io_inAddr_21 == 5'hf; // @[Switch.scala 30:53:@2503.4]
  assign valid_15_21 = io_inValid_21 & _T_7716; // @[Switch.scala 30:36:@2504.4]
  assign _T_7719 = io_inAddr_22 == 5'hf; // @[Switch.scala 30:53:@2506.4]
  assign valid_15_22 = io_inValid_22 & _T_7719; // @[Switch.scala 30:36:@2507.4]
  assign _T_7722 = io_inAddr_23 == 5'hf; // @[Switch.scala 30:53:@2509.4]
  assign valid_15_23 = io_inValid_23 & _T_7722; // @[Switch.scala 30:36:@2510.4]
  assign _T_7725 = io_inAddr_24 == 5'hf; // @[Switch.scala 30:53:@2512.4]
  assign valid_15_24 = io_inValid_24 & _T_7725; // @[Switch.scala 30:36:@2513.4]
  assign _T_7728 = io_inAddr_25 == 5'hf; // @[Switch.scala 30:53:@2515.4]
  assign valid_15_25 = io_inValid_25 & _T_7728; // @[Switch.scala 30:36:@2516.4]
  assign _T_7731 = io_inAddr_26 == 5'hf; // @[Switch.scala 30:53:@2518.4]
  assign valid_15_26 = io_inValid_26 & _T_7731; // @[Switch.scala 30:36:@2519.4]
  assign _T_7734 = io_inAddr_27 == 5'hf; // @[Switch.scala 30:53:@2521.4]
  assign valid_15_27 = io_inValid_27 & _T_7734; // @[Switch.scala 30:36:@2522.4]
  assign _T_7737 = io_inAddr_28 == 5'hf; // @[Switch.scala 30:53:@2524.4]
  assign valid_15_28 = io_inValid_28 & _T_7737; // @[Switch.scala 30:36:@2525.4]
  assign _T_7740 = io_inAddr_29 == 5'hf; // @[Switch.scala 30:53:@2527.4]
  assign valid_15_29 = io_inValid_29 & _T_7740; // @[Switch.scala 30:36:@2528.4]
  assign _T_7743 = io_inAddr_30 == 5'hf; // @[Switch.scala 30:53:@2530.4]
  assign valid_15_30 = io_inValid_30 & _T_7743; // @[Switch.scala 30:36:@2531.4]
  assign _T_7746 = io_inAddr_31 == 5'hf; // @[Switch.scala 30:53:@2533.4]
  assign valid_15_31 = io_inValid_31 & _T_7746; // @[Switch.scala 30:36:@2534.4]
  assign _T_7780 = valid_15_30 ? 5'h1e : 5'h1f; // @[Mux.scala 31:69:@2536.4]
  assign _T_7781 = valid_15_29 ? 5'h1d : _T_7780; // @[Mux.scala 31:69:@2537.4]
  assign _T_7782 = valid_15_28 ? 5'h1c : _T_7781; // @[Mux.scala 31:69:@2538.4]
  assign _T_7783 = valid_15_27 ? 5'h1b : _T_7782; // @[Mux.scala 31:69:@2539.4]
  assign _T_7784 = valid_15_26 ? 5'h1a : _T_7783; // @[Mux.scala 31:69:@2540.4]
  assign _T_7785 = valid_15_25 ? 5'h19 : _T_7784; // @[Mux.scala 31:69:@2541.4]
  assign _T_7786 = valid_15_24 ? 5'h18 : _T_7785; // @[Mux.scala 31:69:@2542.4]
  assign _T_7787 = valid_15_23 ? 5'h17 : _T_7786; // @[Mux.scala 31:69:@2543.4]
  assign _T_7788 = valid_15_22 ? 5'h16 : _T_7787; // @[Mux.scala 31:69:@2544.4]
  assign _T_7789 = valid_15_21 ? 5'h15 : _T_7788; // @[Mux.scala 31:69:@2545.4]
  assign _T_7790 = valid_15_20 ? 5'h14 : _T_7789; // @[Mux.scala 31:69:@2546.4]
  assign _T_7791 = valid_15_19 ? 5'h13 : _T_7790; // @[Mux.scala 31:69:@2547.4]
  assign _T_7792 = valid_15_18 ? 5'h12 : _T_7791; // @[Mux.scala 31:69:@2548.4]
  assign _T_7793 = valid_15_17 ? 5'h11 : _T_7792; // @[Mux.scala 31:69:@2549.4]
  assign _T_7794 = valid_15_16 ? 5'h10 : _T_7793; // @[Mux.scala 31:69:@2550.4]
  assign _T_7795 = valid_15_15 ? 5'hf : _T_7794; // @[Mux.scala 31:69:@2551.4]
  assign _T_7796 = valid_15_14 ? 5'he : _T_7795; // @[Mux.scala 31:69:@2552.4]
  assign _T_7797 = valid_15_13 ? 5'hd : _T_7796; // @[Mux.scala 31:69:@2553.4]
  assign _T_7798 = valid_15_12 ? 5'hc : _T_7797; // @[Mux.scala 31:69:@2554.4]
  assign _T_7799 = valid_15_11 ? 5'hb : _T_7798; // @[Mux.scala 31:69:@2555.4]
  assign _T_7800 = valid_15_10 ? 5'ha : _T_7799; // @[Mux.scala 31:69:@2556.4]
  assign _T_7801 = valid_15_9 ? 5'h9 : _T_7800; // @[Mux.scala 31:69:@2557.4]
  assign _T_7802 = valid_15_8 ? 5'h8 : _T_7801; // @[Mux.scala 31:69:@2558.4]
  assign _T_7803 = valid_15_7 ? 5'h7 : _T_7802; // @[Mux.scala 31:69:@2559.4]
  assign _T_7804 = valid_15_6 ? 5'h6 : _T_7803; // @[Mux.scala 31:69:@2560.4]
  assign _T_7805 = valid_15_5 ? 5'h5 : _T_7804; // @[Mux.scala 31:69:@2561.4]
  assign _T_7806 = valid_15_4 ? 5'h4 : _T_7805; // @[Mux.scala 31:69:@2562.4]
  assign _T_7807 = valid_15_3 ? 5'h3 : _T_7806; // @[Mux.scala 31:69:@2563.4]
  assign _T_7808 = valid_15_2 ? 5'h2 : _T_7807; // @[Mux.scala 31:69:@2564.4]
  assign _T_7809 = valid_15_1 ? 5'h1 : _T_7808; // @[Mux.scala 31:69:@2565.4]
  assign select_15 = valid_15_0 ? 5'h0 : _T_7809; // @[Mux.scala 31:69:@2566.4]
  assign _GEN_481 = 5'h1 == select_15 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@2568.4]
  assign _GEN_482 = 5'h2 == select_15 ? io_inData_2 : _GEN_481; // @[Switch.scala 33:19:@2568.4]
  assign _GEN_483 = 5'h3 == select_15 ? io_inData_3 : _GEN_482; // @[Switch.scala 33:19:@2568.4]
  assign _GEN_484 = 5'h4 == select_15 ? io_inData_4 : _GEN_483; // @[Switch.scala 33:19:@2568.4]
  assign _GEN_485 = 5'h5 == select_15 ? io_inData_5 : _GEN_484; // @[Switch.scala 33:19:@2568.4]
  assign _GEN_486 = 5'h6 == select_15 ? io_inData_6 : _GEN_485; // @[Switch.scala 33:19:@2568.4]
  assign _GEN_487 = 5'h7 == select_15 ? io_inData_7 : _GEN_486; // @[Switch.scala 33:19:@2568.4]
  assign _GEN_488 = 5'h8 == select_15 ? io_inData_8 : _GEN_487; // @[Switch.scala 33:19:@2568.4]
  assign _GEN_489 = 5'h9 == select_15 ? io_inData_9 : _GEN_488; // @[Switch.scala 33:19:@2568.4]
  assign _GEN_490 = 5'ha == select_15 ? io_inData_10 : _GEN_489; // @[Switch.scala 33:19:@2568.4]
  assign _GEN_491 = 5'hb == select_15 ? io_inData_11 : _GEN_490; // @[Switch.scala 33:19:@2568.4]
  assign _GEN_492 = 5'hc == select_15 ? io_inData_12 : _GEN_491; // @[Switch.scala 33:19:@2568.4]
  assign _GEN_493 = 5'hd == select_15 ? io_inData_13 : _GEN_492; // @[Switch.scala 33:19:@2568.4]
  assign _GEN_494 = 5'he == select_15 ? io_inData_14 : _GEN_493; // @[Switch.scala 33:19:@2568.4]
  assign _GEN_495 = 5'hf == select_15 ? io_inData_15 : _GEN_494; // @[Switch.scala 33:19:@2568.4]
  assign _GEN_496 = 5'h10 == select_15 ? io_inData_16 : _GEN_495; // @[Switch.scala 33:19:@2568.4]
  assign _GEN_497 = 5'h11 == select_15 ? io_inData_17 : _GEN_496; // @[Switch.scala 33:19:@2568.4]
  assign _GEN_498 = 5'h12 == select_15 ? io_inData_18 : _GEN_497; // @[Switch.scala 33:19:@2568.4]
  assign _GEN_499 = 5'h13 == select_15 ? io_inData_19 : _GEN_498; // @[Switch.scala 33:19:@2568.4]
  assign _GEN_500 = 5'h14 == select_15 ? io_inData_20 : _GEN_499; // @[Switch.scala 33:19:@2568.4]
  assign _GEN_501 = 5'h15 == select_15 ? io_inData_21 : _GEN_500; // @[Switch.scala 33:19:@2568.4]
  assign _GEN_502 = 5'h16 == select_15 ? io_inData_22 : _GEN_501; // @[Switch.scala 33:19:@2568.4]
  assign _GEN_503 = 5'h17 == select_15 ? io_inData_23 : _GEN_502; // @[Switch.scala 33:19:@2568.4]
  assign _GEN_504 = 5'h18 == select_15 ? io_inData_24 : _GEN_503; // @[Switch.scala 33:19:@2568.4]
  assign _GEN_505 = 5'h19 == select_15 ? io_inData_25 : _GEN_504; // @[Switch.scala 33:19:@2568.4]
  assign _GEN_506 = 5'h1a == select_15 ? io_inData_26 : _GEN_505; // @[Switch.scala 33:19:@2568.4]
  assign _GEN_507 = 5'h1b == select_15 ? io_inData_27 : _GEN_506; // @[Switch.scala 33:19:@2568.4]
  assign _GEN_508 = 5'h1c == select_15 ? io_inData_28 : _GEN_507; // @[Switch.scala 33:19:@2568.4]
  assign _GEN_509 = 5'h1d == select_15 ? io_inData_29 : _GEN_508; // @[Switch.scala 33:19:@2568.4]
  assign _GEN_510 = 5'h1e == select_15 ? io_inData_30 : _GEN_509; // @[Switch.scala 33:19:@2568.4]
  assign _T_7818 = {valid_15_7,valid_15_6,valid_15_5,valid_15_4,valid_15_3,valid_15_2,valid_15_1,valid_15_0}; // @[Switch.scala 34:32:@2575.4]
  assign _T_7826 = {valid_15_15,valid_15_14,valid_15_13,valid_15_12,valid_15_11,valid_15_10,valid_15_9,valid_15_8,_T_7818}; // @[Switch.scala 34:32:@2583.4]
  assign _T_7833 = {valid_15_23,valid_15_22,valid_15_21,valid_15_20,valid_15_19,valid_15_18,valid_15_17,valid_15_16}; // @[Switch.scala 34:32:@2590.4]
  assign _T_7842 = {valid_15_31,valid_15_30,valid_15_29,valid_15_28,valid_15_27,valid_15_26,valid_15_25,valid_15_24,_T_7833,_T_7826}; // @[Switch.scala 34:32:@2599.4]
  assign _T_7846 = io_inAddr_0 == 5'h10; // @[Switch.scala 30:53:@2602.4]
  assign valid_16_0 = io_inValid_0 & _T_7846; // @[Switch.scala 30:36:@2603.4]
  assign _T_7849 = io_inAddr_1 == 5'h10; // @[Switch.scala 30:53:@2605.4]
  assign valid_16_1 = io_inValid_1 & _T_7849; // @[Switch.scala 30:36:@2606.4]
  assign _T_7852 = io_inAddr_2 == 5'h10; // @[Switch.scala 30:53:@2608.4]
  assign valid_16_2 = io_inValid_2 & _T_7852; // @[Switch.scala 30:36:@2609.4]
  assign _T_7855 = io_inAddr_3 == 5'h10; // @[Switch.scala 30:53:@2611.4]
  assign valid_16_3 = io_inValid_3 & _T_7855; // @[Switch.scala 30:36:@2612.4]
  assign _T_7858 = io_inAddr_4 == 5'h10; // @[Switch.scala 30:53:@2614.4]
  assign valid_16_4 = io_inValid_4 & _T_7858; // @[Switch.scala 30:36:@2615.4]
  assign _T_7861 = io_inAddr_5 == 5'h10; // @[Switch.scala 30:53:@2617.4]
  assign valid_16_5 = io_inValid_5 & _T_7861; // @[Switch.scala 30:36:@2618.4]
  assign _T_7864 = io_inAddr_6 == 5'h10; // @[Switch.scala 30:53:@2620.4]
  assign valid_16_6 = io_inValid_6 & _T_7864; // @[Switch.scala 30:36:@2621.4]
  assign _T_7867 = io_inAddr_7 == 5'h10; // @[Switch.scala 30:53:@2623.4]
  assign valid_16_7 = io_inValid_7 & _T_7867; // @[Switch.scala 30:36:@2624.4]
  assign _T_7870 = io_inAddr_8 == 5'h10; // @[Switch.scala 30:53:@2626.4]
  assign valid_16_8 = io_inValid_8 & _T_7870; // @[Switch.scala 30:36:@2627.4]
  assign _T_7873 = io_inAddr_9 == 5'h10; // @[Switch.scala 30:53:@2629.4]
  assign valid_16_9 = io_inValid_9 & _T_7873; // @[Switch.scala 30:36:@2630.4]
  assign _T_7876 = io_inAddr_10 == 5'h10; // @[Switch.scala 30:53:@2632.4]
  assign valid_16_10 = io_inValid_10 & _T_7876; // @[Switch.scala 30:36:@2633.4]
  assign _T_7879 = io_inAddr_11 == 5'h10; // @[Switch.scala 30:53:@2635.4]
  assign valid_16_11 = io_inValid_11 & _T_7879; // @[Switch.scala 30:36:@2636.4]
  assign _T_7882 = io_inAddr_12 == 5'h10; // @[Switch.scala 30:53:@2638.4]
  assign valid_16_12 = io_inValid_12 & _T_7882; // @[Switch.scala 30:36:@2639.4]
  assign _T_7885 = io_inAddr_13 == 5'h10; // @[Switch.scala 30:53:@2641.4]
  assign valid_16_13 = io_inValid_13 & _T_7885; // @[Switch.scala 30:36:@2642.4]
  assign _T_7888 = io_inAddr_14 == 5'h10; // @[Switch.scala 30:53:@2644.4]
  assign valid_16_14 = io_inValid_14 & _T_7888; // @[Switch.scala 30:36:@2645.4]
  assign _T_7891 = io_inAddr_15 == 5'h10; // @[Switch.scala 30:53:@2647.4]
  assign valid_16_15 = io_inValid_15 & _T_7891; // @[Switch.scala 30:36:@2648.4]
  assign _T_7894 = io_inAddr_16 == 5'h10; // @[Switch.scala 30:53:@2650.4]
  assign valid_16_16 = io_inValid_16 & _T_7894; // @[Switch.scala 30:36:@2651.4]
  assign _T_7897 = io_inAddr_17 == 5'h10; // @[Switch.scala 30:53:@2653.4]
  assign valid_16_17 = io_inValid_17 & _T_7897; // @[Switch.scala 30:36:@2654.4]
  assign _T_7900 = io_inAddr_18 == 5'h10; // @[Switch.scala 30:53:@2656.4]
  assign valid_16_18 = io_inValid_18 & _T_7900; // @[Switch.scala 30:36:@2657.4]
  assign _T_7903 = io_inAddr_19 == 5'h10; // @[Switch.scala 30:53:@2659.4]
  assign valid_16_19 = io_inValid_19 & _T_7903; // @[Switch.scala 30:36:@2660.4]
  assign _T_7906 = io_inAddr_20 == 5'h10; // @[Switch.scala 30:53:@2662.4]
  assign valid_16_20 = io_inValid_20 & _T_7906; // @[Switch.scala 30:36:@2663.4]
  assign _T_7909 = io_inAddr_21 == 5'h10; // @[Switch.scala 30:53:@2665.4]
  assign valid_16_21 = io_inValid_21 & _T_7909; // @[Switch.scala 30:36:@2666.4]
  assign _T_7912 = io_inAddr_22 == 5'h10; // @[Switch.scala 30:53:@2668.4]
  assign valid_16_22 = io_inValid_22 & _T_7912; // @[Switch.scala 30:36:@2669.4]
  assign _T_7915 = io_inAddr_23 == 5'h10; // @[Switch.scala 30:53:@2671.4]
  assign valid_16_23 = io_inValid_23 & _T_7915; // @[Switch.scala 30:36:@2672.4]
  assign _T_7918 = io_inAddr_24 == 5'h10; // @[Switch.scala 30:53:@2674.4]
  assign valid_16_24 = io_inValid_24 & _T_7918; // @[Switch.scala 30:36:@2675.4]
  assign _T_7921 = io_inAddr_25 == 5'h10; // @[Switch.scala 30:53:@2677.4]
  assign valid_16_25 = io_inValid_25 & _T_7921; // @[Switch.scala 30:36:@2678.4]
  assign _T_7924 = io_inAddr_26 == 5'h10; // @[Switch.scala 30:53:@2680.4]
  assign valid_16_26 = io_inValid_26 & _T_7924; // @[Switch.scala 30:36:@2681.4]
  assign _T_7927 = io_inAddr_27 == 5'h10; // @[Switch.scala 30:53:@2683.4]
  assign valid_16_27 = io_inValid_27 & _T_7927; // @[Switch.scala 30:36:@2684.4]
  assign _T_7930 = io_inAddr_28 == 5'h10; // @[Switch.scala 30:53:@2686.4]
  assign valid_16_28 = io_inValid_28 & _T_7930; // @[Switch.scala 30:36:@2687.4]
  assign _T_7933 = io_inAddr_29 == 5'h10; // @[Switch.scala 30:53:@2689.4]
  assign valid_16_29 = io_inValid_29 & _T_7933; // @[Switch.scala 30:36:@2690.4]
  assign _T_7936 = io_inAddr_30 == 5'h10; // @[Switch.scala 30:53:@2692.4]
  assign valid_16_30 = io_inValid_30 & _T_7936; // @[Switch.scala 30:36:@2693.4]
  assign _T_7939 = io_inAddr_31 == 5'h10; // @[Switch.scala 30:53:@2695.4]
  assign valid_16_31 = io_inValid_31 & _T_7939; // @[Switch.scala 30:36:@2696.4]
  assign _T_7973 = valid_16_30 ? 5'h1e : 5'h1f; // @[Mux.scala 31:69:@2698.4]
  assign _T_7974 = valid_16_29 ? 5'h1d : _T_7973; // @[Mux.scala 31:69:@2699.4]
  assign _T_7975 = valid_16_28 ? 5'h1c : _T_7974; // @[Mux.scala 31:69:@2700.4]
  assign _T_7976 = valid_16_27 ? 5'h1b : _T_7975; // @[Mux.scala 31:69:@2701.4]
  assign _T_7977 = valid_16_26 ? 5'h1a : _T_7976; // @[Mux.scala 31:69:@2702.4]
  assign _T_7978 = valid_16_25 ? 5'h19 : _T_7977; // @[Mux.scala 31:69:@2703.4]
  assign _T_7979 = valid_16_24 ? 5'h18 : _T_7978; // @[Mux.scala 31:69:@2704.4]
  assign _T_7980 = valid_16_23 ? 5'h17 : _T_7979; // @[Mux.scala 31:69:@2705.4]
  assign _T_7981 = valid_16_22 ? 5'h16 : _T_7980; // @[Mux.scala 31:69:@2706.4]
  assign _T_7982 = valid_16_21 ? 5'h15 : _T_7981; // @[Mux.scala 31:69:@2707.4]
  assign _T_7983 = valid_16_20 ? 5'h14 : _T_7982; // @[Mux.scala 31:69:@2708.4]
  assign _T_7984 = valid_16_19 ? 5'h13 : _T_7983; // @[Mux.scala 31:69:@2709.4]
  assign _T_7985 = valid_16_18 ? 5'h12 : _T_7984; // @[Mux.scala 31:69:@2710.4]
  assign _T_7986 = valid_16_17 ? 5'h11 : _T_7985; // @[Mux.scala 31:69:@2711.4]
  assign _T_7987 = valid_16_16 ? 5'h10 : _T_7986; // @[Mux.scala 31:69:@2712.4]
  assign _T_7988 = valid_16_15 ? 5'hf : _T_7987; // @[Mux.scala 31:69:@2713.4]
  assign _T_7989 = valid_16_14 ? 5'he : _T_7988; // @[Mux.scala 31:69:@2714.4]
  assign _T_7990 = valid_16_13 ? 5'hd : _T_7989; // @[Mux.scala 31:69:@2715.4]
  assign _T_7991 = valid_16_12 ? 5'hc : _T_7990; // @[Mux.scala 31:69:@2716.4]
  assign _T_7992 = valid_16_11 ? 5'hb : _T_7991; // @[Mux.scala 31:69:@2717.4]
  assign _T_7993 = valid_16_10 ? 5'ha : _T_7992; // @[Mux.scala 31:69:@2718.4]
  assign _T_7994 = valid_16_9 ? 5'h9 : _T_7993; // @[Mux.scala 31:69:@2719.4]
  assign _T_7995 = valid_16_8 ? 5'h8 : _T_7994; // @[Mux.scala 31:69:@2720.4]
  assign _T_7996 = valid_16_7 ? 5'h7 : _T_7995; // @[Mux.scala 31:69:@2721.4]
  assign _T_7997 = valid_16_6 ? 5'h6 : _T_7996; // @[Mux.scala 31:69:@2722.4]
  assign _T_7998 = valid_16_5 ? 5'h5 : _T_7997; // @[Mux.scala 31:69:@2723.4]
  assign _T_7999 = valid_16_4 ? 5'h4 : _T_7998; // @[Mux.scala 31:69:@2724.4]
  assign _T_8000 = valid_16_3 ? 5'h3 : _T_7999; // @[Mux.scala 31:69:@2725.4]
  assign _T_8001 = valid_16_2 ? 5'h2 : _T_8000; // @[Mux.scala 31:69:@2726.4]
  assign _T_8002 = valid_16_1 ? 5'h1 : _T_8001; // @[Mux.scala 31:69:@2727.4]
  assign select_16 = valid_16_0 ? 5'h0 : _T_8002; // @[Mux.scala 31:69:@2728.4]
  assign _GEN_513 = 5'h1 == select_16 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@2730.4]
  assign _GEN_514 = 5'h2 == select_16 ? io_inData_2 : _GEN_513; // @[Switch.scala 33:19:@2730.4]
  assign _GEN_515 = 5'h3 == select_16 ? io_inData_3 : _GEN_514; // @[Switch.scala 33:19:@2730.4]
  assign _GEN_516 = 5'h4 == select_16 ? io_inData_4 : _GEN_515; // @[Switch.scala 33:19:@2730.4]
  assign _GEN_517 = 5'h5 == select_16 ? io_inData_5 : _GEN_516; // @[Switch.scala 33:19:@2730.4]
  assign _GEN_518 = 5'h6 == select_16 ? io_inData_6 : _GEN_517; // @[Switch.scala 33:19:@2730.4]
  assign _GEN_519 = 5'h7 == select_16 ? io_inData_7 : _GEN_518; // @[Switch.scala 33:19:@2730.4]
  assign _GEN_520 = 5'h8 == select_16 ? io_inData_8 : _GEN_519; // @[Switch.scala 33:19:@2730.4]
  assign _GEN_521 = 5'h9 == select_16 ? io_inData_9 : _GEN_520; // @[Switch.scala 33:19:@2730.4]
  assign _GEN_522 = 5'ha == select_16 ? io_inData_10 : _GEN_521; // @[Switch.scala 33:19:@2730.4]
  assign _GEN_523 = 5'hb == select_16 ? io_inData_11 : _GEN_522; // @[Switch.scala 33:19:@2730.4]
  assign _GEN_524 = 5'hc == select_16 ? io_inData_12 : _GEN_523; // @[Switch.scala 33:19:@2730.4]
  assign _GEN_525 = 5'hd == select_16 ? io_inData_13 : _GEN_524; // @[Switch.scala 33:19:@2730.4]
  assign _GEN_526 = 5'he == select_16 ? io_inData_14 : _GEN_525; // @[Switch.scala 33:19:@2730.4]
  assign _GEN_527 = 5'hf == select_16 ? io_inData_15 : _GEN_526; // @[Switch.scala 33:19:@2730.4]
  assign _GEN_528 = 5'h10 == select_16 ? io_inData_16 : _GEN_527; // @[Switch.scala 33:19:@2730.4]
  assign _GEN_529 = 5'h11 == select_16 ? io_inData_17 : _GEN_528; // @[Switch.scala 33:19:@2730.4]
  assign _GEN_530 = 5'h12 == select_16 ? io_inData_18 : _GEN_529; // @[Switch.scala 33:19:@2730.4]
  assign _GEN_531 = 5'h13 == select_16 ? io_inData_19 : _GEN_530; // @[Switch.scala 33:19:@2730.4]
  assign _GEN_532 = 5'h14 == select_16 ? io_inData_20 : _GEN_531; // @[Switch.scala 33:19:@2730.4]
  assign _GEN_533 = 5'h15 == select_16 ? io_inData_21 : _GEN_532; // @[Switch.scala 33:19:@2730.4]
  assign _GEN_534 = 5'h16 == select_16 ? io_inData_22 : _GEN_533; // @[Switch.scala 33:19:@2730.4]
  assign _GEN_535 = 5'h17 == select_16 ? io_inData_23 : _GEN_534; // @[Switch.scala 33:19:@2730.4]
  assign _GEN_536 = 5'h18 == select_16 ? io_inData_24 : _GEN_535; // @[Switch.scala 33:19:@2730.4]
  assign _GEN_537 = 5'h19 == select_16 ? io_inData_25 : _GEN_536; // @[Switch.scala 33:19:@2730.4]
  assign _GEN_538 = 5'h1a == select_16 ? io_inData_26 : _GEN_537; // @[Switch.scala 33:19:@2730.4]
  assign _GEN_539 = 5'h1b == select_16 ? io_inData_27 : _GEN_538; // @[Switch.scala 33:19:@2730.4]
  assign _GEN_540 = 5'h1c == select_16 ? io_inData_28 : _GEN_539; // @[Switch.scala 33:19:@2730.4]
  assign _GEN_541 = 5'h1d == select_16 ? io_inData_29 : _GEN_540; // @[Switch.scala 33:19:@2730.4]
  assign _GEN_542 = 5'h1e == select_16 ? io_inData_30 : _GEN_541; // @[Switch.scala 33:19:@2730.4]
  assign _T_8011 = {valid_16_7,valid_16_6,valid_16_5,valid_16_4,valid_16_3,valid_16_2,valid_16_1,valid_16_0}; // @[Switch.scala 34:32:@2737.4]
  assign _T_8019 = {valid_16_15,valid_16_14,valid_16_13,valid_16_12,valid_16_11,valid_16_10,valid_16_9,valid_16_8,_T_8011}; // @[Switch.scala 34:32:@2745.4]
  assign _T_8026 = {valid_16_23,valid_16_22,valid_16_21,valid_16_20,valid_16_19,valid_16_18,valid_16_17,valid_16_16}; // @[Switch.scala 34:32:@2752.4]
  assign _T_8035 = {valid_16_31,valid_16_30,valid_16_29,valid_16_28,valid_16_27,valid_16_26,valid_16_25,valid_16_24,_T_8026,_T_8019}; // @[Switch.scala 34:32:@2761.4]
  assign _T_8039 = io_inAddr_0 == 5'h11; // @[Switch.scala 30:53:@2764.4]
  assign valid_17_0 = io_inValid_0 & _T_8039; // @[Switch.scala 30:36:@2765.4]
  assign _T_8042 = io_inAddr_1 == 5'h11; // @[Switch.scala 30:53:@2767.4]
  assign valid_17_1 = io_inValid_1 & _T_8042; // @[Switch.scala 30:36:@2768.4]
  assign _T_8045 = io_inAddr_2 == 5'h11; // @[Switch.scala 30:53:@2770.4]
  assign valid_17_2 = io_inValid_2 & _T_8045; // @[Switch.scala 30:36:@2771.4]
  assign _T_8048 = io_inAddr_3 == 5'h11; // @[Switch.scala 30:53:@2773.4]
  assign valid_17_3 = io_inValid_3 & _T_8048; // @[Switch.scala 30:36:@2774.4]
  assign _T_8051 = io_inAddr_4 == 5'h11; // @[Switch.scala 30:53:@2776.4]
  assign valid_17_4 = io_inValid_4 & _T_8051; // @[Switch.scala 30:36:@2777.4]
  assign _T_8054 = io_inAddr_5 == 5'h11; // @[Switch.scala 30:53:@2779.4]
  assign valid_17_5 = io_inValid_5 & _T_8054; // @[Switch.scala 30:36:@2780.4]
  assign _T_8057 = io_inAddr_6 == 5'h11; // @[Switch.scala 30:53:@2782.4]
  assign valid_17_6 = io_inValid_6 & _T_8057; // @[Switch.scala 30:36:@2783.4]
  assign _T_8060 = io_inAddr_7 == 5'h11; // @[Switch.scala 30:53:@2785.4]
  assign valid_17_7 = io_inValid_7 & _T_8060; // @[Switch.scala 30:36:@2786.4]
  assign _T_8063 = io_inAddr_8 == 5'h11; // @[Switch.scala 30:53:@2788.4]
  assign valid_17_8 = io_inValid_8 & _T_8063; // @[Switch.scala 30:36:@2789.4]
  assign _T_8066 = io_inAddr_9 == 5'h11; // @[Switch.scala 30:53:@2791.4]
  assign valid_17_9 = io_inValid_9 & _T_8066; // @[Switch.scala 30:36:@2792.4]
  assign _T_8069 = io_inAddr_10 == 5'h11; // @[Switch.scala 30:53:@2794.4]
  assign valid_17_10 = io_inValid_10 & _T_8069; // @[Switch.scala 30:36:@2795.4]
  assign _T_8072 = io_inAddr_11 == 5'h11; // @[Switch.scala 30:53:@2797.4]
  assign valid_17_11 = io_inValid_11 & _T_8072; // @[Switch.scala 30:36:@2798.4]
  assign _T_8075 = io_inAddr_12 == 5'h11; // @[Switch.scala 30:53:@2800.4]
  assign valid_17_12 = io_inValid_12 & _T_8075; // @[Switch.scala 30:36:@2801.4]
  assign _T_8078 = io_inAddr_13 == 5'h11; // @[Switch.scala 30:53:@2803.4]
  assign valid_17_13 = io_inValid_13 & _T_8078; // @[Switch.scala 30:36:@2804.4]
  assign _T_8081 = io_inAddr_14 == 5'h11; // @[Switch.scala 30:53:@2806.4]
  assign valid_17_14 = io_inValid_14 & _T_8081; // @[Switch.scala 30:36:@2807.4]
  assign _T_8084 = io_inAddr_15 == 5'h11; // @[Switch.scala 30:53:@2809.4]
  assign valid_17_15 = io_inValid_15 & _T_8084; // @[Switch.scala 30:36:@2810.4]
  assign _T_8087 = io_inAddr_16 == 5'h11; // @[Switch.scala 30:53:@2812.4]
  assign valid_17_16 = io_inValid_16 & _T_8087; // @[Switch.scala 30:36:@2813.4]
  assign _T_8090 = io_inAddr_17 == 5'h11; // @[Switch.scala 30:53:@2815.4]
  assign valid_17_17 = io_inValid_17 & _T_8090; // @[Switch.scala 30:36:@2816.4]
  assign _T_8093 = io_inAddr_18 == 5'h11; // @[Switch.scala 30:53:@2818.4]
  assign valid_17_18 = io_inValid_18 & _T_8093; // @[Switch.scala 30:36:@2819.4]
  assign _T_8096 = io_inAddr_19 == 5'h11; // @[Switch.scala 30:53:@2821.4]
  assign valid_17_19 = io_inValid_19 & _T_8096; // @[Switch.scala 30:36:@2822.4]
  assign _T_8099 = io_inAddr_20 == 5'h11; // @[Switch.scala 30:53:@2824.4]
  assign valid_17_20 = io_inValid_20 & _T_8099; // @[Switch.scala 30:36:@2825.4]
  assign _T_8102 = io_inAddr_21 == 5'h11; // @[Switch.scala 30:53:@2827.4]
  assign valid_17_21 = io_inValid_21 & _T_8102; // @[Switch.scala 30:36:@2828.4]
  assign _T_8105 = io_inAddr_22 == 5'h11; // @[Switch.scala 30:53:@2830.4]
  assign valid_17_22 = io_inValid_22 & _T_8105; // @[Switch.scala 30:36:@2831.4]
  assign _T_8108 = io_inAddr_23 == 5'h11; // @[Switch.scala 30:53:@2833.4]
  assign valid_17_23 = io_inValid_23 & _T_8108; // @[Switch.scala 30:36:@2834.4]
  assign _T_8111 = io_inAddr_24 == 5'h11; // @[Switch.scala 30:53:@2836.4]
  assign valid_17_24 = io_inValid_24 & _T_8111; // @[Switch.scala 30:36:@2837.4]
  assign _T_8114 = io_inAddr_25 == 5'h11; // @[Switch.scala 30:53:@2839.4]
  assign valid_17_25 = io_inValid_25 & _T_8114; // @[Switch.scala 30:36:@2840.4]
  assign _T_8117 = io_inAddr_26 == 5'h11; // @[Switch.scala 30:53:@2842.4]
  assign valid_17_26 = io_inValid_26 & _T_8117; // @[Switch.scala 30:36:@2843.4]
  assign _T_8120 = io_inAddr_27 == 5'h11; // @[Switch.scala 30:53:@2845.4]
  assign valid_17_27 = io_inValid_27 & _T_8120; // @[Switch.scala 30:36:@2846.4]
  assign _T_8123 = io_inAddr_28 == 5'h11; // @[Switch.scala 30:53:@2848.4]
  assign valid_17_28 = io_inValid_28 & _T_8123; // @[Switch.scala 30:36:@2849.4]
  assign _T_8126 = io_inAddr_29 == 5'h11; // @[Switch.scala 30:53:@2851.4]
  assign valid_17_29 = io_inValid_29 & _T_8126; // @[Switch.scala 30:36:@2852.4]
  assign _T_8129 = io_inAddr_30 == 5'h11; // @[Switch.scala 30:53:@2854.4]
  assign valid_17_30 = io_inValid_30 & _T_8129; // @[Switch.scala 30:36:@2855.4]
  assign _T_8132 = io_inAddr_31 == 5'h11; // @[Switch.scala 30:53:@2857.4]
  assign valid_17_31 = io_inValid_31 & _T_8132; // @[Switch.scala 30:36:@2858.4]
  assign _T_8166 = valid_17_30 ? 5'h1e : 5'h1f; // @[Mux.scala 31:69:@2860.4]
  assign _T_8167 = valid_17_29 ? 5'h1d : _T_8166; // @[Mux.scala 31:69:@2861.4]
  assign _T_8168 = valid_17_28 ? 5'h1c : _T_8167; // @[Mux.scala 31:69:@2862.4]
  assign _T_8169 = valid_17_27 ? 5'h1b : _T_8168; // @[Mux.scala 31:69:@2863.4]
  assign _T_8170 = valid_17_26 ? 5'h1a : _T_8169; // @[Mux.scala 31:69:@2864.4]
  assign _T_8171 = valid_17_25 ? 5'h19 : _T_8170; // @[Mux.scala 31:69:@2865.4]
  assign _T_8172 = valid_17_24 ? 5'h18 : _T_8171; // @[Mux.scala 31:69:@2866.4]
  assign _T_8173 = valid_17_23 ? 5'h17 : _T_8172; // @[Mux.scala 31:69:@2867.4]
  assign _T_8174 = valid_17_22 ? 5'h16 : _T_8173; // @[Mux.scala 31:69:@2868.4]
  assign _T_8175 = valid_17_21 ? 5'h15 : _T_8174; // @[Mux.scala 31:69:@2869.4]
  assign _T_8176 = valid_17_20 ? 5'h14 : _T_8175; // @[Mux.scala 31:69:@2870.4]
  assign _T_8177 = valid_17_19 ? 5'h13 : _T_8176; // @[Mux.scala 31:69:@2871.4]
  assign _T_8178 = valid_17_18 ? 5'h12 : _T_8177; // @[Mux.scala 31:69:@2872.4]
  assign _T_8179 = valid_17_17 ? 5'h11 : _T_8178; // @[Mux.scala 31:69:@2873.4]
  assign _T_8180 = valid_17_16 ? 5'h10 : _T_8179; // @[Mux.scala 31:69:@2874.4]
  assign _T_8181 = valid_17_15 ? 5'hf : _T_8180; // @[Mux.scala 31:69:@2875.4]
  assign _T_8182 = valid_17_14 ? 5'he : _T_8181; // @[Mux.scala 31:69:@2876.4]
  assign _T_8183 = valid_17_13 ? 5'hd : _T_8182; // @[Mux.scala 31:69:@2877.4]
  assign _T_8184 = valid_17_12 ? 5'hc : _T_8183; // @[Mux.scala 31:69:@2878.4]
  assign _T_8185 = valid_17_11 ? 5'hb : _T_8184; // @[Mux.scala 31:69:@2879.4]
  assign _T_8186 = valid_17_10 ? 5'ha : _T_8185; // @[Mux.scala 31:69:@2880.4]
  assign _T_8187 = valid_17_9 ? 5'h9 : _T_8186; // @[Mux.scala 31:69:@2881.4]
  assign _T_8188 = valid_17_8 ? 5'h8 : _T_8187; // @[Mux.scala 31:69:@2882.4]
  assign _T_8189 = valid_17_7 ? 5'h7 : _T_8188; // @[Mux.scala 31:69:@2883.4]
  assign _T_8190 = valid_17_6 ? 5'h6 : _T_8189; // @[Mux.scala 31:69:@2884.4]
  assign _T_8191 = valid_17_5 ? 5'h5 : _T_8190; // @[Mux.scala 31:69:@2885.4]
  assign _T_8192 = valid_17_4 ? 5'h4 : _T_8191; // @[Mux.scala 31:69:@2886.4]
  assign _T_8193 = valid_17_3 ? 5'h3 : _T_8192; // @[Mux.scala 31:69:@2887.4]
  assign _T_8194 = valid_17_2 ? 5'h2 : _T_8193; // @[Mux.scala 31:69:@2888.4]
  assign _T_8195 = valid_17_1 ? 5'h1 : _T_8194; // @[Mux.scala 31:69:@2889.4]
  assign select_17 = valid_17_0 ? 5'h0 : _T_8195; // @[Mux.scala 31:69:@2890.4]
  assign _GEN_545 = 5'h1 == select_17 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@2892.4]
  assign _GEN_546 = 5'h2 == select_17 ? io_inData_2 : _GEN_545; // @[Switch.scala 33:19:@2892.4]
  assign _GEN_547 = 5'h3 == select_17 ? io_inData_3 : _GEN_546; // @[Switch.scala 33:19:@2892.4]
  assign _GEN_548 = 5'h4 == select_17 ? io_inData_4 : _GEN_547; // @[Switch.scala 33:19:@2892.4]
  assign _GEN_549 = 5'h5 == select_17 ? io_inData_5 : _GEN_548; // @[Switch.scala 33:19:@2892.4]
  assign _GEN_550 = 5'h6 == select_17 ? io_inData_6 : _GEN_549; // @[Switch.scala 33:19:@2892.4]
  assign _GEN_551 = 5'h7 == select_17 ? io_inData_7 : _GEN_550; // @[Switch.scala 33:19:@2892.4]
  assign _GEN_552 = 5'h8 == select_17 ? io_inData_8 : _GEN_551; // @[Switch.scala 33:19:@2892.4]
  assign _GEN_553 = 5'h9 == select_17 ? io_inData_9 : _GEN_552; // @[Switch.scala 33:19:@2892.4]
  assign _GEN_554 = 5'ha == select_17 ? io_inData_10 : _GEN_553; // @[Switch.scala 33:19:@2892.4]
  assign _GEN_555 = 5'hb == select_17 ? io_inData_11 : _GEN_554; // @[Switch.scala 33:19:@2892.4]
  assign _GEN_556 = 5'hc == select_17 ? io_inData_12 : _GEN_555; // @[Switch.scala 33:19:@2892.4]
  assign _GEN_557 = 5'hd == select_17 ? io_inData_13 : _GEN_556; // @[Switch.scala 33:19:@2892.4]
  assign _GEN_558 = 5'he == select_17 ? io_inData_14 : _GEN_557; // @[Switch.scala 33:19:@2892.4]
  assign _GEN_559 = 5'hf == select_17 ? io_inData_15 : _GEN_558; // @[Switch.scala 33:19:@2892.4]
  assign _GEN_560 = 5'h10 == select_17 ? io_inData_16 : _GEN_559; // @[Switch.scala 33:19:@2892.4]
  assign _GEN_561 = 5'h11 == select_17 ? io_inData_17 : _GEN_560; // @[Switch.scala 33:19:@2892.4]
  assign _GEN_562 = 5'h12 == select_17 ? io_inData_18 : _GEN_561; // @[Switch.scala 33:19:@2892.4]
  assign _GEN_563 = 5'h13 == select_17 ? io_inData_19 : _GEN_562; // @[Switch.scala 33:19:@2892.4]
  assign _GEN_564 = 5'h14 == select_17 ? io_inData_20 : _GEN_563; // @[Switch.scala 33:19:@2892.4]
  assign _GEN_565 = 5'h15 == select_17 ? io_inData_21 : _GEN_564; // @[Switch.scala 33:19:@2892.4]
  assign _GEN_566 = 5'h16 == select_17 ? io_inData_22 : _GEN_565; // @[Switch.scala 33:19:@2892.4]
  assign _GEN_567 = 5'h17 == select_17 ? io_inData_23 : _GEN_566; // @[Switch.scala 33:19:@2892.4]
  assign _GEN_568 = 5'h18 == select_17 ? io_inData_24 : _GEN_567; // @[Switch.scala 33:19:@2892.4]
  assign _GEN_569 = 5'h19 == select_17 ? io_inData_25 : _GEN_568; // @[Switch.scala 33:19:@2892.4]
  assign _GEN_570 = 5'h1a == select_17 ? io_inData_26 : _GEN_569; // @[Switch.scala 33:19:@2892.4]
  assign _GEN_571 = 5'h1b == select_17 ? io_inData_27 : _GEN_570; // @[Switch.scala 33:19:@2892.4]
  assign _GEN_572 = 5'h1c == select_17 ? io_inData_28 : _GEN_571; // @[Switch.scala 33:19:@2892.4]
  assign _GEN_573 = 5'h1d == select_17 ? io_inData_29 : _GEN_572; // @[Switch.scala 33:19:@2892.4]
  assign _GEN_574 = 5'h1e == select_17 ? io_inData_30 : _GEN_573; // @[Switch.scala 33:19:@2892.4]
  assign _T_8204 = {valid_17_7,valid_17_6,valid_17_5,valid_17_4,valid_17_3,valid_17_2,valid_17_1,valid_17_0}; // @[Switch.scala 34:32:@2899.4]
  assign _T_8212 = {valid_17_15,valid_17_14,valid_17_13,valid_17_12,valid_17_11,valid_17_10,valid_17_9,valid_17_8,_T_8204}; // @[Switch.scala 34:32:@2907.4]
  assign _T_8219 = {valid_17_23,valid_17_22,valid_17_21,valid_17_20,valid_17_19,valid_17_18,valid_17_17,valid_17_16}; // @[Switch.scala 34:32:@2914.4]
  assign _T_8228 = {valid_17_31,valid_17_30,valid_17_29,valid_17_28,valid_17_27,valid_17_26,valid_17_25,valid_17_24,_T_8219,_T_8212}; // @[Switch.scala 34:32:@2923.4]
  assign _T_8232 = io_inAddr_0 == 5'h12; // @[Switch.scala 30:53:@2926.4]
  assign valid_18_0 = io_inValid_0 & _T_8232; // @[Switch.scala 30:36:@2927.4]
  assign _T_8235 = io_inAddr_1 == 5'h12; // @[Switch.scala 30:53:@2929.4]
  assign valid_18_1 = io_inValid_1 & _T_8235; // @[Switch.scala 30:36:@2930.4]
  assign _T_8238 = io_inAddr_2 == 5'h12; // @[Switch.scala 30:53:@2932.4]
  assign valid_18_2 = io_inValid_2 & _T_8238; // @[Switch.scala 30:36:@2933.4]
  assign _T_8241 = io_inAddr_3 == 5'h12; // @[Switch.scala 30:53:@2935.4]
  assign valid_18_3 = io_inValid_3 & _T_8241; // @[Switch.scala 30:36:@2936.4]
  assign _T_8244 = io_inAddr_4 == 5'h12; // @[Switch.scala 30:53:@2938.4]
  assign valid_18_4 = io_inValid_4 & _T_8244; // @[Switch.scala 30:36:@2939.4]
  assign _T_8247 = io_inAddr_5 == 5'h12; // @[Switch.scala 30:53:@2941.4]
  assign valid_18_5 = io_inValid_5 & _T_8247; // @[Switch.scala 30:36:@2942.4]
  assign _T_8250 = io_inAddr_6 == 5'h12; // @[Switch.scala 30:53:@2944.4]
  assign valid_18_6 = io_inValid_6 & _T_8250; // @[Switch.scala 30:36:@2945.4]
  assign _T_8253 = io_inAddr_7 == 5'h12; // @[Switch.scala 30:53:@2947.4]
  assign valid_18_7 = io_inValid_7 & _T_8253; // @[Switch.scala 30:36:@2948.4]
  assign _T_8256 = io_inAddr_8 == 5'h12; // @[Switch.scala 30:53:@2950.4]
  assign valid_18_8 = io_inValid_8 & _T_8256; // @[Switch.scala 30:36:@2951.4]
  assign _T_8259 = io_inAddr_9 == 5'h12; // @[Switch.scala 30:53:@2953.4]
  assign valid_18_9 = io_inValid_9 & _T_8259; // @[Switch.scala 30:36:@2954.4]
  assign _T_8262 = io_inAddr_10 == 5'h12; // @[Switch.scala 30:53:@2956.4]
  assign valid_18_10 = io_inValid_10 & _T_8262; // @[Switch.scala 30:36:@2957.4]
  assign _T_8265 = io_inAddr_11 == 5'h12; // @[Switch.scala 30:53:@2959.4]
  assign valid_18_11 = io_inValid_11 & _T_8265; // @[Switch.scala 30:36:@2960.4]
  assign _T_8268 = io_inAddr_12 == 5'h12; // @[Switch.scala 30:53:@2962.4]
  assign valid_18_12 = io_inValid_12 & _T_8268; // @[Switch.scala 30:36:@2963.4]
  assign _T_8271 = io_inAddr_13 == 5'h12; // @[Switch.scala 30:53:@2965.4]
  assign valid_18_13 = io_inValid_13 & _T_8271; // @[Switch.scala 30:36:@2966.4]
  assign _T_8274 = io_inAddr_14 == 5'h12; // @[Switch.scala 30:53:@2968.4]
  assign valid_18_14 = io_inValid_14 & _T_8274; // @[Switch.scala 30:36:@2969.4]
  assign _T_8277 = io_inAddr_15 == 5'h12; // @[Switch.scala 30:53:@2971.4]
  assign valid_18_15 = io_inValid_15 & _T_8277; // @[Switch.scala 30:36:@2972.4]
  assign _T_8280 = io_inAddr_16 == 5'h12; // @[Switch.scala 30:53:@2974.4]
  assign valid_18_16 = io_inValid_16 & _T_8280; // @[Switch.scala 30:36:@2975.4]
  assign _T_8283 = io_inAddr_17 == 5'h12; // @[Switch.scala 30:53:@2977.4]
  assign valid_18_17 = io_inValid_17 & _T_8283; // @[Switch.scala 30:36:@2978.4]
  assign _T_8286 = io_inAddr_18 == 5'h12; // @[Switch.scala 30:53:@2980.4]
  assign valid_18_18 = io_inValid_18 & _T_8286; // @[Switch.scala 30:36:@2981.4]
  assign _T_8289 = io_inAddr_19 == 5'h12; // @[Switch.scala 30:53:@2983.4]
  assign valid_18_19 = io_inValid_19 & _T_8289; // @[Switch.scala 30:36:@2984.4]
  assign _T_8292 = io_inAddr_20 == 5'h12; // @[Switch.scala 30:53:@2986.4]
  assign valid_18_20 = io_inValid_20 & _T_8292; // @[Switch.scala 30:36:@2987.4]
  assign _T_8295 = io_inAddr_21 == 5'h12; // @[Switch.scala 30:53:@2989.4]
  assign valid_18_21 = io_inValid_21 & _T_8295; // @[Switch.scala 30:36:@2990.4]
  assign _T_8298 = io_inAddr_22 == 5'h12; // @[Switch.scala 30:53:@2992.4]
  assign valid_18_22 = io_inValid_22 & _T_8298; // @[Switch.scala 30:36:@2993.4]
  assign _T_8301 = io_inAddr_23 == 5'h12; // @[Switch.scala 30:53:@2995.4]
  assign valid_18_23 = io_inValid_23 & _T_8301; // @[Switch.scala 30:36:@2996.4]
  assign _T_8304 = io_inAddr_24 == 5'h12; // @[Switch.scala 30:53:@2998.4]
  assign valid_18_24 = io_inValid_24 & _T_8304; // @[Switch.scala 30:36:@2999.4]
  assign _T_8307 = io_inAddr_25 == 5'h12; // @[Switch.scala 30:53:@3001.4]
  assign valid_18_25 = io_inValid_25 & _T_8307; // @[Switch.scala 30:36:@3002.4]
  assign _T_8310 = io_inAddr_26 == 5'h12; // @[Switch.scala 30:53:@3004.4]
  assign valid_18_26 = io_inValid_26 & _T_8310; // @[Switch.scala 30:36:@3005.4]
  assign _T_8313 = io_inAddr_27 == 5'h12; // @[Switch.scala 30:53:@3007.4]
  assign valid_18_27 = io_inValid_27 & _T_8313; // @[Switch.scala 30:36:@3008.4]
  assign _T_8316 = io_inAddr_28 == 5'h12; // @[Switch.scala 30:53:@3010.4]
  assign valid_18_28 = io_inValid_28 & _T_8316; // @[Switch.scala 30:36:@3011.4]
  assign _T_8319 = io_inAddr_29 == 5'h12; // @[Switch.scala 30:53:@3013.4]
  assign valid_18_29 = io_inValid_29 & _T_8319; // @[Switch.scala 30:36:@3014.4]
  assign _T_8322 = io_inAddr_30 == 5'h12; // @[Switch.scala 30:53:@3016.4]
  assign valid_18_30 = io_inValid_30 & _T_8322; // @[Switch.scala 30:36:@3017.4]
  assign _T_8325 = io_inAddr_31 == 5'h12; // @[Switch.scala 30:53:@3019.4]
  assign valid_18_31 = io_inValid_31 & _T_8325; // @[Switch.scala 30:36:@3020.4]
  assign _T_8359 = valid_18_30 ? 5'h1e : 5'h1f; // @[Mux.scala 31:69:@3022.4]
  assign _T_8360 = valid_18_29 ? 5'h1d : _T_8359; // @[Mux.scala 31:69:@3023.4]
  assign _T_8361 = valid_18_28 ? 5'h1c : _T_8360; // @[Mux.scala 31:69:@3024.4]
  assign _T_8362 = valid_18_27 ? 5'h1b : _T_8361; // @[Mux.scala 31:69:@3025.4]
  assign _T_8363 = valid_18_26 ? 5'h1a : _T_8362; // @[Mux.scala 31:69:@3026.4]
  assign _T_8364 = valid_18_25 ? 5'h19 : _T_8363; // @[Mux.scala 31:69:@3027.4]
  assign _T_8365 = valid_18_24 ? 5'h18 : _T_8364; // @[Mux.scala 31:69:@3028.4]
  assign _T_8366 = valid_18_23 ? 5'h17 : _T_8365; // @[Mux.scala 31:69:@3029.4]
  assign _T_8367 = valid_18_22 ? 5'h16 : _T_8366; // @[Mux.scala 31:69:@3030.4]
  assign _T_8368 = valid_18_21 ? 5'h15 : _T_8367; // @[Mux.scala 31:69:@3031.4]
  assign _T_8369 = valid_18_20 ? 5'h14 : _T_8368; // @[Mux.scala 31:69:@3032.4]
  assign _T_8370 = valid_18_19 ? 5'h13 : _T_8369; // @[Mux.scala 31:69:@3033.4]
  assign _T_8371 = valid_18_18 ? 5'h12 : _T_8370; // @[Mux.scala 31:69:@3034.4]
  assign _T_8372 = valid_18_17 ? 5'h11 : _T_8371; // @[Mux.scala 31:69:@3035.4]
  assign _T_8373 = valid_18_16 ? 5'h10 : _T_8372; // @[Mux.scala 31:69:@3036.4]
  assign _T_8374 = valid_18_15 ? 5'hf : _T_8373; // @[Mux.scala 31:69:@3037.4]
  assign _T_8375 = valid_18_14 ? 5'he : _T_8374; // @[Mux.scala 31:69:@3038.4]
  assign _T_8376 = valid_18_13 ? 5'hd : _T_8375; // @[Mux.scala 31:69:@3039.4]
  assign _T_8377 = valid_18_12 ? 5'hc : _T_8376; // @[Mux.scala 31:69:@3040.4]
  assign _T_8378 = valid_18_11 ? 5'hb : _T_8377; // @[Mux.scala 31:69:@3041.4]
  assign _T_8379 = valid_18_10 ? 5'ha : _T_8378; // @[Mux.scala 31:69:@3042.4]
  assign _T_8380 = valid_18_9 ? 5'h9 : _T_8379; // @[Mux.scala 31:69:@3043.4]
  assign _T_8381 = valid_18_8 ? 5'h8 : _T_8380; // @[Mux.scala 31:69:@3044.4]
  assign _T_8382 = valid_18_7 ? 5'h7 : _T_8381; // @[Mux.scala 31:69:@3045.4]
  assign _T_8383 = valid_18_6 ? 5'h6 : _T_8382; // @[Mux.scala 31:69:@3046.4]
  assign _T_8384 = valid_18_5 ? 5'h5 : _T_8383; // @[Mux.scala 31:69:@3047.4]
  assign _T_8385 = valid_18_4 ? 5'h4 : _T_8384; // @[Mux.scala 31:69:@3048.4]
  assign _T_8386 = valid_18_3 ? 5'h3 : _T_8385; // @[Mux.scala 31:69:@3049.4]
  assign _T_8387 = valid_18_2 ? 5'h2 : _T_8386; // @[Mux.scala 31:69:@3050.4]
  assign _T_8388 = valid_18_1 ? 5'h1 : _T_8387; // @[Mux.scala 31:69:@3051.4]
  assign select_18 = valid_18_0 ? 5'h0 : _T_8388; // @[Mux.scala 31:69:@3052.4]
  assign _GEN_577 = 5'h1 == select_18 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@3054.4]
  assign _GEN_578 = 5'h2 == select_18 ? io_inData_2 : _GEN_577; // @[Switch.scala 33:19:@3054.4]
  assign _GEN_579 = 5'h3 == select_18 ? io_inData_3 : _GEN_578; // @[Switch.scala 33:19:@3054.4]
  assign _GEN_580 = 5'h4 == select_18 ? io_inData_4 : _GEN_579; // @[Switch.scala 33:19:@3054.4]
  assign _GEN_581 = 5'h5 == select_18 ? io_inData_5 : _GEN_580; // @[Switch.scala 33:19:@3054.4]
  assign _GEN_582 = 5'h6 == select_18 ? io_inData_6 : _GEN_581; // @[Switch.scala 33:19:@3054.4]
  assign _GEN_583 = 5'h7 == select_18 ? io_inData_7 : _GEN_582; // @[Switch.scala 33:19:@3054.4]
  assign _GEN_584 = 5'h8 == select_18 ? io_inData_8 : _GEN_583; // @[Switch.scala 33:19:@3054.4]
  assign _GEN_585 = 5'h9 == select_18 ? io_inData_9 : _GEN_584; // @[Switch.scala 33:19:@3054.4]
  assign _GEN_586 = 5'ha == select_18 ? io_inData_10 : _GEN_585; // @[Switch.scala 33:19:@3054.4]
  assign _GEN_587 = 5'hb == select_18 ? io_inData_11 : _GEN_586; // @[Switch.scala 33:19:@3054.4]
  assign _GEN_588 = 5'hc == select_18 ? io_inData_12 : _GEN_587; // @[Switch.scala 33:19:@3054.4]
  assign _GEN_589 = 5'hd == select_18 ? io_inData_13 : _GEN_588; // @[Switch.scala 33:19:@3054.4]
  assign _GEN_590 = 5'he == select_18 ? io_inData_14 : _GEN_589; // @[Switch.scala 33:19:@3054.4]
  assign _GEN_591 = 5'hf == select_18 ? io_inData_15 : _GEN_590; // @[Switch.scala 33:19:@3054.4]
  assign _GEN_592 = 5'h10 == select_18 ? io_inData_16 : _GEN_591; // @[Switch.scala 33:19:@3054.4]
  assign _GEN_593 = 5'h11 == select_18 ? io_inData_17 : _GEN_592; // @[Switch.scala 33:19:@3054.4]
  assign _GEN_594 = 5'h12 == select_18 ? io_inData_18 : _GEN_593; // @[Switch.scala 33:19:@3054.4]
  assign _GEN_595 = 5'h13 == select_18 ? io_inData_19 : _GEN_594; // @[Switch.scala 33:19:@3054.4]
  assign _GEN_596 = 5'h14 == select_18 ? io_inData_20 : _GEN_595; // @[Switch.scala 33:19:@3054.4]
  assign _GEN_597 = 5'h15 == select_18 ? io_inData_21 : _GEN_596; // @[Switch.scala 33:19:@3054.4]
  assign _GEN_598 = 5'h16 == select_18 ? io_inData_22 : _GEN_597; // @[Switch.scala 33:19:@3054.4]
  assign _GEN_599 = 5'h17 == select_18 ? io_inData_23 : _GEN_598; // @[Switch.scala 33:19:@3054.4]
  assign _GEN_600 = 5'h18 == select_18 ? io_inData_24 : _GEN_599; // @[Switch.scala 33:19:@3054.4]
  assign _GEN_601 = 5'h19 == select_18 ? io_inData_25 : _GEN_600; // @[Switch.scala 33:19:@3054.4]
  assign _GEN_602 = 5'h1a == select_18 ? io_inData_26 : _GEN_601; // @[Switch.scala 33:19:@3054.4]
  assign _GEN_603 = 5'h1b == select_18 ? io_inData_27 : _GEN_602; // @[Switch.scala 33:19:@3054.4]
  assign _GEN_604 = 5'h1c == select_18 ? io_inData_28 : _GEN_603; // @[Switch.scala 33:19:@3054.4]
  assign _GEN_605 = 5'h1d == select_18 ? io_inData_29 : _GEN_604; // @[Switch.scala 33:19:@3054.4]
  assign _GEN_606 = 5'h1e == select_18 ? io_inData_30 : _GEN_605; // @[Switch.scala 33:19:@3054.4]
  assign _T_8397 = {valid_18_7,valid_18_6,valid_18_5,valid_18_4,valid_18_3,valid_18_2,valid_18_1,valid_18_0}; // @[Switch.scala 34:32:@3061.4]
  assign _T_8405 = {valid_18_15,valid_18_14,valid_18_13,valid_18_12,valid_18_11,valid_18_10,valid_18_9,valid_18_8,_T_8397}; // @[Switch.scala 34:32:@3069.4]
  assign _T_8412 = {valid_18_23,valid_18_22,valid_18_21,valid_18_20,valid_18_19,valid_18_18,valid_18_17,valid_18_16}; // @[Switch.scala 34:32:@3076.4]
  assign _T_8421 = {valid_18_31,valid_18_30,valid_18_29,valid_18_28,valid_18_27,valid_18_26,valid_18_25,valid_18_24,_T_8412,_T_8405}; // @[Switch.scala 34:32:@3085.4]
  assign _T_8425 = io_inAddr_0 == 5'h13; // @[Switch.scala 30:53:@3088.4]
  assign valid_19_0 = io_inValid_0 & _T_8425; // @[Switch.scala 30:36:@3089.4]
  assign _T_8428 = io_inAddr_1 == 5'h13; // @[Switch.scala 30:53:@3091.4]
  assign valid_19_1 = io_inValid_1 & _T_8428; // @[Switch.scala 30:36:@3092.4]
  assign _T_8431 = io_inAddr_2 == 5'h13; // @[Switch.scala 30:53:@3094.4]
  assign valid_19_2 = io_inValid_2 & _T_8431; // @[Switch.scala 30:36:@3095.4]
  assign _T_8434 = io_inAddr_3 == 5'h13; // @[Switch.scala 30:53:@3097.4]
  assign valid_19_3 = io_inValid_3 & _T_8434; // @[Switch.scala 30:36:@3098.4]
  assign _T_8437 = io_inAddr_4 == 5'h13; // @[Switch.scala 30:53:@3100.4]
  assign valid_19_4 = io_inValid_4 & _T_8437; // @[Switch.scala 30:36:@3101.4]
  assign _T_8440 = io_inAddr_5 == 5'h13; // @[Switch.scala 30:53:@3103.4]
  assign valid_19_5 = io_inValid_5 & _T_8440; // @[Switch.scala 30:36:@3104.4]
  assign _T_8443 = io_inAddr_6 == 5'h13; // @[Switch.scala 30:53:@3106.4]
  assign valid_19_6 = io_inValid_6 & _T_8443; // @[Switch.scala 30:36:@3107.4]
  assign _T_8446 = io_inAddr_7 == 5'h13; // @[Switch.scala 30:53:@3109.4]
  assign valid_19_7 = io_inValid_7 & _T_8446; // @[Switch.scala 30:36:@3110.4]
  assign _T_8449 = io_inAddr_8 == 5'h13; // @[Switch.scala 30:53:@3112.4]
  assign valid_19_8 = io_inValid_8 & _T_8449; // @[Switch.scala 30:36:@3113.4]
  assign _T_8452 = io_inAddr_9 == 5'h13; // @[Switch.scala 30:53:@3115.4]
  assign valid_19_9 = io_inValid_9 & _T_8452; // @[Switch.scala 30:36:@3116.4]
  assign _T_8455 = io_inAddr_10 == 5'h13; // @[Switch.scala 30:53:@3118.4]
  assign valid_19_10 = io_inValid_10 & _T_8455; // @[Switch.scala 30:36:@3119.4]
  assign _T_8458 = io_inAddr_11 == 5'h13; // @[Switch.scala 30:53:@3121.4]
  assign valid_19_11 = io_inValid_11 & _T_8458; // @[Switch.scala 30:36:@3122.4]
  assign _T_8461 = io_inAddr_12 == 5'h13; // @[Switch.scala 30:53:@3124.4]
  assign valid_19_12 = io_inValid_12 & _T_8461; // @[Switch.scala 30:36:@3125.4]
  assign _T_8464 = io_inAddr_13 == 5'h13; // @[Switch.scala 30:53:@3127.4]
  assign valid_19_13 = io_inValid_13 & _T_8464; // @[Switch.scala 30:36:@3128.4]
  assign _T_8467 = io_inAddr_14 == 5'h13; // @[Switch.scala 30:53:@3130.4]
  assign valid_19_14 = io_inValid_14 & _T_8467; // @[Switch.scala 30:36:@3131.4]
  assign _T_8470 = io_inAddr_15 == 5'h13; // @[Switch.scala 30:53:@3133.4]
  assign valid_19_15 = io_inValid_15 & _T_8470; // @[Switch.scala 30:36:@3134.4]
  assign _T_8473 = io_inAddr_16 == 5'h13; // @[Switch.scala 30:53:@3136.4]
  assign valid_19_16 = io_inValid_16 & _T_8473; // @[Switch.scala 30:36:@3137.4]
  assign _T_8476 = io_inAddr_17 == 5'h13; // @[Switch.scala 30:53:@3139.4]
  assign valid_19_17 = io_inValid_17 & _T_8476; // @[Switch.scala 30:36:@3140.4]
  assign _T_8479 = io_inAddr_18 == 5'h13; // @[Switch.scala 30:53:@3142.4]
  assign valid_19_18 = io_inValid_18 & _T_8479; // @[Switch.scala 30:36:@3143.4]
  assign _T_8482 = io_inAddr_19 == 5'h13; // @[Switch.scala 30:53:@3145.4]
  assign valid_19_19 = io_inValid_19 & _T_8482; // @[Switch.scala 30:36:@3146.4]
  assign _T_8485 = io_inAddr_20 == 5'h13; // @[Switch.scala 30:53:@3148.4]
  assign valid_19_20 = io_inValid_20 & _T_8485; // @[Switch.scala 30:36:@3149.4]
  assign _T_8488 = io_inAddr_21 == 5'h13; // @[Switch.scala 30:53:@3151.4]
  assign valid_19_21 = io_inValid_21 & _T_8488; // @[Switch.scala 30:36:@3152.4]
  assign _T_8491 = io_inAddr_22 == 5'h13; // @[Switch.scala 30:53:@3154.4]
  assign valid_19_22 = io_inValid_22 & _T_8491; // @[Switch.scala 30:36:@3155.4]
  assign _T_8494 = io_inAddr_23 == 5'h13; // @[Switch.scala 30:53:@3157.4]
  assign valid_19_23 = io_inValid_23 & _T_8494; // @[Switch.scala 30:36:@3158.4]
  assign _T_8497 = io_inAddr_24 == 5'h13; // @[Switch.scala 30:53:@3160.4]
  assign valid_19_24 = io_inValid_24 & _T_8497; // @[Switch.scala 30:36:@3161.4]
  assign _T_8500 = io_inAddr_25 == 5'h13; // @[Switch.scala 30:53:@3163.4]
  assign valid_19_25 = io_inValid_25 & _T_8500; // @[Switch.scala 30:36:@3164.4]
  assign _T_8503 = io_inAddr_26 == 5'h13; // @[Switch.scala 30:53:@3166.4]
  assign valid_19_26 = io_inValid_26 & _T_8503; // @[Switch.scala 30:36:@3167.4]
  assign _T_8506 = io_inAddr_27 == 5'h13; // @[Switch.scala 30:53:@3169.4]
  assign valid_19_27 = io_inValid_27 & _T_8506; // @[Switch.scala 30:36:@3170.4]
  assign _T_8509 = io_inAddr_28 == 5'h13; // @[Switch.scala 30:53:@3172.4]
  assign valid_19_28 = io_inValid_28 & _T_8509; // @[Switch.scala 30:36:@3173.4]
  assign _T_8512 = io_inAddr_29 == 5'h13; // @[Switch.scala 30:53:@3175.4]
  assign valid_19_29 = io_inValid_29 & _T_8512; // @[Switch.scala 30:36:@3176.4]
  assign _T_8515 = io_inAddr_30 == 5'h13; // @[Switch.scala 30:53:@3178.4]
  assign valid_19_30 = io_inValid_30 & _T_8515; // @[Switch.scala 30:36:@3179.4]
  assign _T_8518 = io_inAddr_31 == 5'h13; // @[Switch.scala 30:53:@3181.4]
  assign valid_19_31 = io_inValid_31 & _T_8518; // @[Switch.scala 30:36:@3182.4]
  assign _T_8552 = valid_19_30 ? 5'h1e : 5'h1f; // @[Mux.scala 31:69:@3184.4]
  assign _T_8553 = valid_19_29 ? 5'h1d : _T_8552; // @[Mux.scala 31:69:@3185.4]
  assign _T_8554 = valid_19_28 ? 5'h1c : _T_8553; // @[Mux.scala 31:69:@3186.4]
  assign _T_8555 = valid_19_27 ? 5'h1b : _T_8554; // @[Mux.scala 31:69:@3187.4]
  assign _T_8556 = valid_19_26 ? 5'h1a : _T_8555; // @[Mux.scala 31:69:@3188.4]
  assign _T_8557 = valid_19_25 ? 5'h19 : _T_8556; // @[Mux.scala 31:69:@3189.4]
  assign _T_8558 = valid_19_24 ? 5'h18 : _T_8557; // @[Mux.scala 31:69:@3190.4]
  assign _T_8559 = valid_19_23 ? 5'h17 : _T_8558; // @[Mux.scala 31:69:@3191.4]
  assign _T_8560 = valid_19_22 ? 5'h16 : _T_8559; // @[Mux.scala 31:69:@3192.4]
  assign _T_8561 = valid_19_21 ? 5'h15 : _T_8560; // @[Mux.scala 31:69:@3193.4]
  assign _T_8562 = valid_19_20 ? 5'h14 : _T_8561; // @[Mux.scala 31:69:@3194.4]
  assign _T_8563 = valid_19_19 ? 5'h13 : _T_8562; // @[Mux.scala 31:69:@3195.4]
  assign _T_8564 = valid_19_18 ? 5'h12 : _T_8563; // @[Mux.scala 31:69:@3196.4]
  assign _T_8565 = valid_19_17 ? 5'h11 : _T_8564; // @[Mux.scala 31:69:@3197.4]
  assign _T_8566 = valid_19_16 ? 5'h10 : _T_8565; // @[Mux.scala 31:69:@3198.4]
  assign _T_8567 = valid_19_15 ? 5'hf : _T_8566; // @[Mux.scala 31:69:@3199.4]
  assign _T_8568 = valid_19_14 ? 5'he : _T_8567; // @[Mux.scala 31:69:@3200.4]
  assign _T_8569 = valid_19_13 ? 5'hd : _T_8568; // @[Mux.scala 31:69:@3201.4]
  assign _T_8570 = valid_19_12 ? 5'hc : _T_8569; // @[Mux.scala 31:69:@3202.4]
  assign _T_8571 = valid_19_11 ? 5'hb : _T_8570; // @[Mux.scala 31:69:@3203.4]
  assign _T_8572 = valid_19_10 ? 5'ha : _T_8571; // @[Mux.scala 31:69:@3204.4]
  assign _T_8573 = valid_19_9 ? 5'h9 : _T_8572; // @[Mux.scala 31:69:@3205.4]
  assign _T_8574 = valid_19_8 ? 5'h8 : _T_8573; // @[Mux.scala 31:69:@3206.4]
  assign _T_8575 = valid_19_7 ? 5'h7 : _T_8574; // @[Mux.scala 31:69:@3207.4]
  assign _T_8576 = valid_19_6 ? 5'h6 : _T_8575; // @[Mux.scala 31:69:@3208.4]
  assign _T_8577 = valid_19_5 ? 5'h5 : _T_8576; // @[Mux.scala 31:69:@3209.4]
  assign _T_8578 = valid_19_4 ? 5'h4 : _T_8577; // @[Mux.scala 31:69:@3210.4]
  assign _T_8579 = valid_19_3 ? 5'h3 : _T_8578; // @[Mux.scala 31:69:@3211.4]
  assign _T_8580 = valid_19_2 ? 5'h2 : _T_8579; // @[Mux.scala 31:69:@3212.4]
  assign _T_8581 = valid_19_1 ? 5'h1 : _T_8580; // @[Mux.scala 31:69:@3213.4]
  assign select_19 = valid_19_0 ? 5'h0 : _T_8581; // @[Mux.scala 31:69:@3214.4]
  assign _GEN_609 = 5'h1 == select_19 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@3216.4]
  assign _GEN_610 = 5'h2 == select_19 ? io_inData_2 : _GEN_609; // @[Switch.scala 33:19:@3216.4]
  assign _GEN_611 = 5'h3 == select_19 ? io_inData_3 : _GEN_610; // @[Switch.scala 33:19:@3216.4]
  assign _GEN_612 = 5'h4 == select_19 ? io_inData_4 : _GEN_611; // @[Switch.scala 33:19:@3216.4]
  assign _GEN_613 = 5'h5 == select_19 ? io_inData_5 : _GEN_612; // @[Switch.scala 33:19:@3216.4]
  assign _GEN_614 = 5'h6 == select_19 ? io_inData_6 : _GEN_613; // @[Switch.scala 33:19:@3216.4]
  assign _GEN_615 = 5'h7 == select_19 ? io_inData_7 : _GEN_614; // @[Switch.scala 33:19:@3216.4]
  assign _GEN_616 = 5'h8 == select_19 ? io_inData_8 : _GEN_615; // @[Switch.scala 33:19:@3216.4]
  assign _GEN_617 = 5'h9 == select_19 ? io_inData_9 : _GEN_616; // @[Switch.scala 33:19:@3216.4]
  assign _GEN_618 = 5'ha == select_19 ? io_inData_10 : _GEN_617; // @[Switch.scala 33:19:@3216.4]
  assign _GEN_619 = 5'hb == select_19 ? io_inData_11 : _GEN_618; // @[Switch.scala 33:19:@3216.4]
  assign _GEN_620 = 5'hc == select_19 ? io_inData_12 : _GEN_619; // @[Switch.scala 33:19:@3216.4]
  assign _GEN_621 = 5'hd == select_19 ? io_inData_13 : _GEN_620; // @[Switch.scala 33:19:@3216.4]
  assign _GEN_622 = 5'he == select_19 ? io_inData_14 : _GEN_621; // @[Switch.scala 33:19:@3216.4]
  assign _GEN_623 = 5'hf == select_19 ? io_inData_15 : _GEN_622; // @[Switch.scala 33:19:@3216.4]
  assign _GEN_624 = 5'h10 == select_19 ? io_inData_16 : _GEN_623; // @[Switch.scala 33:19:@3216.4]
  assign _GEN_625 = 5'h11 == select_19 ? io_inData_17 : _GEN_624; // @[Switch.scala 33:19:@3216.4]
  assign _GEN_626 = 5'h12 == select_19 ? io_inData_18 : _GEN_625; // @[Switch.scala 33:19:@3216.4]
  assign _GEN_627 = 5'h13 == select_19 ? io_inData_19 : _GEN_626; // @[Switch.scala 33:19:@3216.4]
  assign _GEN_628 = 5'h14 == select_19 ? io_inData_20 : _GEN_627; // @[Switch.scala 33:19:@3216.4]
  assign _GEN_629 = 5'h15 == select_19 ? io_inData_21 : _GEN_628; // @[Switch.scala 33:19:@3216.4]
  assign _GEN_630 = 5'h16 == select_19 ? io_inData_22 : _GEN_629; // @[Switch.scala 33:19:@3216.4]
  assign _GEN_631 = 5'h17 == select_19 ? io_inData_23 : _GEN_630; // @[Switch.scala 33:19:@3216.4]
  assign _GEN_632 = 5'h18 == select_19 ? io_inData_24 : _GEN_631; // @[Switch.scala 33:19:@3216.4]
  assign _GEN_633 = 5'h19 == select_19 ? io_inData_25 : _GEN_632; // @[Switch.scala 33:19:@3216.4]
  assign _GEN_634 = 5'h1a == select_19 ? io_inData_26 : _GEN_633; // @[Switch.scala 33:19:@3216.4]
  assign _GEN_635 = 5'h1b == select_19 ? io_inData_27 : _GEN_634; // @[Switch.scala 33:19:@3216.4]
  assign _GEN_636 = 5'h1c == select_19 ? io_inData_28 : _GEN_635; // @[Switch.scala 33:19:@3216.4]
  assign _GEN_637 = 5'h1d == select_19 ? io_inData_29 : _GEN_636; // @[Switch.scala 33:19:@3216.4]
  assign _GEN_638 = 5'h1e == select_19 ? io_inData_30 : _GEN_637; // @[Switch.scala 33:19:@3216.4]
  assign _T_8590 = {valid_19_7,valid_19_6,valid_19_5,valid_19_4,valid_19_3,valid_19_2,valid_19_1,valid_19_0}; // @[Switch.scala 34:32:@3223.4]
  assign _T_8598 = {valid_19_15,valid_19_14,valid_19_13,valid_19_12,valid_19_11,valid_19_10,valid_19_9,valid_19_8,_T_8590}; // @[Switch.scala 34:32:@3231.4]
  assign _T_8605 = {valid_19_23,valid_19_22,valid_19_21,valid_19_20,valid_19_19,valid_19_18,valid_19_17,valid_19_16}; // @[Switch.scala 34:32:@3238.4]
  assign _T_8614 = {valid_19_31,valid_19_30,valid_19_29,valid_19_28,valid_19_27,valid_19_26,valid_19_25,valid_19_24,_T_8605,_T_8598}; // @[Switch.scala 34:32:@3247.4]
  assign _T_8618 = io_inAddr_0 == 5'h14; // @[Switch.scala 30:53:@3250.4]
  assign valid_20_0 = io_inValid_0 & _T_8618; // @[Switch.scala 30:36:@3251.4]
  assign _T_8621 = io_inAddr_1 == 5'h14; // @[Switch.scala 30:53:@3253.4]
  assign valid_20_1 = io_inValid_1 & _T_8621; // @[Switch.scala 30:36:@3254.4]
  assign _T_8624 = io_inAddr_2 == 5'h14; // @[Switch.scala 30:53:@3256.4]
  assign valid_20_2 = io_inValid_2 & _T_8624; // @[Switch.scala 30:36:@3257.4]
  assign _T_8627 = io_inAddr_3 == 5'h14; // @[Switch.scala 30:53:@3259.4]
  assign valid_20_3 = io_inValid_3 & _T_8627; // @[Switch.scala 30:36:@3260.4]
  assign _T_8630 = io_inAddr_4 == 5'h14; // @[Switch.scala 30:53:@3262.4]
  assign valid_20_4 = io_inValid_4 & _T_8630; // @[Switch.scala 30:36:@3263.4]
  assign _T_8633 = io_inAddr_5 == 5'h14; // @[Switch.scala 30:53:@3265.4]
  assign valid_20_5 = io_inValid_5 & _T_8633; // @[Switch.scala 30:36:@3266.4]
  assign _T_8636 = io_inAddr_6 == 5'h14; // @[Switch.scala 30:53:@3268.4]
  assign valid_20_6 = io_inValid_6 & _T_8636; // @[Switch.scala 30:36:@3269.4]
  assign _T_8639 = io_inAddr_7 == 5'h14; // @[Switch.scala 30:53:@3271.4]
  assign valid_20_7 = io_inValid_7 & _T_8639; // @[Switch.scala 30:36:@3272.4]
  assign _T_8642 = io_inAddr_8 == 5'h14; // @[Switch.scala 30:53:@3274.4]
  assign valid_20_8 = io_inValid_8 & _T_8642; // @[Switch.scala 30:36:@3275.4]
  assign _T_8645 = io_inAddr_9 == 5'h14; // @[Switch.scala 30:53:@3277.4]
  assign valid_20_9 = io_inValid_9 & _T_8645; // @[Switch.scala 30:36:@3278.4]
  assign _T_8648 = io_inAddr_10 == 5'h14; // @[Switch.scala 30:53:@3280.4]
  assign valid_20_10 = io_inValid_10 & _T_8648; // @[Switch.scala 30:36:@3281.4]
  assign _T_8651 = io_inAddr_11 == 5'h14; // @[Switch.scala 30:53:@3283.4]
  assign valid_20_11 = io_inValid_11 & _T_8651; // @[Switch.scala 30:36:@3284.4]
  assign _T_8654 = io_inAddr_12 == 5'h14; // @[Switch.scala 30:53:@3286.4]
  assign valid_20_12 = io_inValid_12 & _T_8654; // @[Switch.scala 30:36:@3287.4]
  assign _T_8657 = io_inAddr_13 == 5'h14; // @[Switch.scala 30:53:@3289.4]
  assign valid_20_13 = io_inValid_13 & _T_8657; // @[Switch.scala 30:36:@3290.4]
  assign _T_8660 = io_inAddr_14 == 5'h14; // @[Switch.scala 30:53:@3292.4]
  assign valid_20_14 = io_inValid_14 & _T_8660; // @[Switch.scala 30:36:@3293.4]
  assign _T_8663 = io_inAddr_15 == 5'h14; // @[Switch.scala 30:53:@3295.4]
  assign valid_20_15 = io_inValid_15 & _T_8663; // @[Switch.scala 30:36:@3296.4]
  assign _T_8666 = io_inAddr_16 == 5'h14; // @[Switch.scala 30:53:@3298.4]
  assign valid_20_16 = io_inValid_16 & _T_8666; // @[Switch.scala 30:36:@3299.4]
  assign _T_8669 = io_inAddr_17 == 5'h14; // @[Switch.scala 30:53:@3301.4]
  assign valid_20_17 = io_inValid_17 & _T_8669; // @[Switch.scala 30:36:@3302.4]
  assign _T_8672 = io_inAddr_18 == 5'h14; // @[Switch.scala 30:53:@3304.4]
  assign valid_20_18 = io_inValid_18 & _T_8672; // @[Switch.scala 30:36:@3305.4]
  assign _T_8675 = io_inAddr_19 == 5'h14; // @[Switch.scala 30:53:@3307.4]
  assign valid_20_19 = io_inValid_19 & _T_8675; // @[Switch.scala 30:36:@3308.4]
  assign _T_8678 = io_inAddr_20 == 5'h14; // @[Switch.scala 30:53:@3310.4]
  assign valid_20_20 = io_inValid_20 & _T_8678; // @[Switch.scala 30:36:@3311.4]
  assign _T_8681 = io_inAddr_21 == 5'h14; // @[Switch.scala 30:53:@3313.4]
  assign valid_20_21 = io_inValid_21 & _T_8681; // @[Switch.scala 30:36:@3314.4]
  assign _T_8684 = io_inAddr_22 == 5'h14; // @[Switch.scala 30:53:@3316.4]
  assign valid_20_22 = io_inValid_22 & _T_8684; // @[Switch.scala 30:36:@3317.4]
  assign _T_8687 = io_inAddr_23 == 5'h14; // @[Switch.scala 30:53:@3319.4]
  assign valid_20_23 = io_inValid_23 & _T_8687; // @[Switch.scala 30:36:@3320.4]
  assign _T_8690 = io_inAddr_24 == 5'h14; // @[Switch.scala 30:53:@3322.4]
  assign valid_20_24 = io_inValid_24 & _T_8690; // @[Switch.scala 30:36:@3323.4]
  assign _T_8693 = io_inAddr_25 == 5'h14; // @[Switch.scala 30:53:@3325.4]
  assign valid_20_25 = io_inValid_25 & _T_8693; // @[Switch.scala 30:36:@3326.4]
  assign _T_8696 = io_inAddr_26 == 5'h14; // @[Switch.scala 30:53:@3328.4]
  assign valid_20_26 = io_inValid_26 & _T_8696; // @[Switch.scala 30:36:@3329.4]
  assign _T_8699 = io_inAddr_27 == 5'h14; // @[Switch.scala 30:53:@3331.4]
  assign valid_20_27 = io_inValid_27 & _T_8699; // @[Switch.scala 30:36:@3332.4]
  assign _T_8702 = io_inAddr_28 == 5'h14; // @[Switch.scala 30:53:@3334.4]
  assign valid_20_28 = io_inValid_28 & _T_8702; // @[Switch.scala 30:36:@3335.4]
  assign _T_8705 = io_inAddr_29 == 5'h14; // @[Switch.scala 30:53:@3337.4]
  assign valid_20_29 = io_inValid_29 & _T_8705; // @[Switch.scala 30:36:@3338.4]
  assign _T_8708 = io_inAddr_30 == 5'h14; // @[Switch.scala 30:53:@3340.4]
  assign valid_20_30 = io_inValid_30 & _T_8708; // @[Switch.scala 30:36:@3341.4]
  assign _T_8711 = io_inAddr_31 == 5'h14; // @[Switch.scala 30:53:@3343.4]
  assign valid_20_31 = io_inValid_31 & _T_8711; // @[Switch.scala 30:36:@3344.4]
  assign _T_8745 = valid_20_30 ? 5'h1e : 5'h1f; // @[Mux.scala 31:69:@3346.4]
  assign _T_8746 = valid_20_29 ? 5'h1d : _T_8745; // @[Mux.scala 31:69:@3347.4]
  assign _T_8747 = valid_20_28 ? 5'h1c : _T_8746; // @[Mux.scala 31:69:@3348.4]
  assign _T_8748 = valid_20_27 ? 5'h1b : _T_8747; // @[Mux.scala 31:69:@3349.4]
  assign _T_8749 = valid_20_26 ? 5'h1a : _T_8748; // @[Mux.scala 31:69:@3350.4]
  assign _T_8750 = valid_20_25 ? 5'h19 : _T_8749; // @[Mux.scala 31:69:@3351.4]
  assign _T_8751 = valid_20_24 ? 5'h18 : _T_8750; // @[Mux.scala 31:69:@3352.4]
  assign _T_8752 = valid_20_23 ? 5'h17 : _T_8751; // @[Mux.scala 31:69:@3353.4]
  assign _T_8753 = valid_20_22 ? 5'h16 : _T_8752; // @[Mux.scala 31:69:@3354.4]
  assign _T_8754 = valid_20_21 ? 5'h15 : _T_8753; // @[Mux.scala 31:69:@3355.4]
  assign _T_8755 = valid_20_20 ? 5'h14 : _T_8754; // @[Mux.scala 31:69:@3356.4]
  assign _T_8756 = valid_20_19 ? 5'h13 : _T_8755; // @[Mux.scala 31:69:@3357.4]
  assign _T_8757 = valid_20_18 ? 5'h12 : _T_8756; // @[Mux.scala 31:69:@3358.4]
  assign _T_8758 = valid_20_17 ? 5'h11 : _T_8757; // @[Mux.scala 31:69:@3359.4]
  assign _T_8759 = valid_20_16 ? 5'h10 : _T_8758; // @[Mux.scala 31:69:@3360.4]
  assign _T_8760 = valid_20_15 ? 5'hf : _T_8759; // @[Mux.scala 31:69:@3361.4]
  assign _T_8761 = valid_20_14 ? 5'he : _T_8760; // @[Mux.scala 31:69:@3362.4]
  assign _T_8762 = valid_20_13 ? 5'hd : _T_8761; // @[Mux.scala 31:69:@3363.4]
  assign _T_8763 = valid_20_12 ? 5'hc : _T_8762; // @[Mux.scala 31:69:@3364.4]
  assign _T_8764 = valid_20_11 ? 5'hb : _T_8763; // @[Mux.scala 31:69:@3365.4]
  assign _T_8765 = valid_20_10 ? 5'ha : _T_8764; // @[Mux.scala 31:69:@3366.4]
  assign _T_8766 = valid_20_9 ? 5'h9 : _T_8765; // @[Mux.scala 31:69:@3367.4]
  assign _T_8767 = valid_20_8 ? 5'h8 : _T_8766; // @[Mux.scala 31:69:@3368.4]
  assign _T_8768 = valid_20_7 ? 5'h7 : _T_8767; // @[Mux.scala 31:69:@3369.4]
  assign _T_8769 = valid_20_6 ? 5'h6 : _T_8768; // @[Mux.scala 31:69:@3370.4]
  assign _T_8770 = valid_20_5 ? 5'h5 : _T_8769; // @[Mux.scala 31:69:@3371.4]
  assign _T_8771 = valid_20_4 ? 5'h4 : _T_8770; // @[Mux.scala 31:69:@3372.4]
  assign _T_8772 = valid_20_3 ? 5'h3 : _T_8771; // @[Mux.scala 31:69:@3373.4]
  assign _T_8773 = valid_20_2 ? 5'h2 : _T_8772; // @[Mux.scala 31:69:@3374.4]
  assign _T_8774 = valid_20_1 ? 5'h1 : _T_8773; // @[Mux.scala 31:69:@3375.4]
  assign select_20 = valid_20_0 ? 5'h0 : _T_8774; // @[Mux.scala 31:69:@3376.4]
  assign _GEN_641 = 5'h1 == select_20 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@3378.4]
  assign _GEN_642 = 5'h2 == select_20 ? io_inData_2 : _GEN_641; // @[Switch.scala 33:19:@3378.4]
  assign _GEN_643 = 5'h3 == select_20 ? io_inData_3 : _GEN_642; // @[Switch.scala 33:19:@3378.4]
  assign _GEN_644 = 5'h4 == select_20 ? io_inData_4 : _GEN_643; // @[Switch.scala 33:19:@3378.4]
  assign _GEN_645 = 5'h5 == select_20 ? io_inData_5 : _GEN_644; // @[Switch.scala 33:19:@3378.4]
  assign _GEN_646 = 5'h6 == select_20 ? io_inData_6 : _GEN_645; // @[Switch.scala 33:19:@3378.4]
  assign _GEN_647 = 5'h7 == select_20 ? io_inData_7 : _GEN_646; // @[Switch.scala 33:19:@3378.4]
  assign _GEN_648 = 5'h8 == select_20 ? io_inData_8 : _GEN_647; // @[Switch.scala 33:19:@3378.4]
  assign _GEN_649 = 5'h9 == select_20 ? io_inData_9 : _GEN_648; // @[Switch.scala 33:19:@3378.4]
  assign _GEN_650 = 5'ha == select_20 ? io_inData_10 : _GEN_649; // @[Switch.scala 33:19:@3378.4]
  assign _GEN_651 = 5'hb == select_20 ? io_inData_11 : _GEN_650; // @[Switch.scala 33:19:@3378.4]
  assign _GEN_652 = 5'hc == select_20 ? io_inData_12 : _GEN_651; // @[Switch.scala 33:19:@3378.4]
  assign _GEN_653 = 5'hd == select_20 ? io_inData_13 : _GEN_652; // @[Switch.scala 33:19:@3378.4]
  assign _GEN_654 = 5'he == select_20 ? io_inData_14 : _GEN_653; // @[Switch.scala 33:19:@3378.4]
  assign _GEN_655 = 5'hf == select_20 ? io_inData_15 : _GEN_654; // @[Switch.scala 33:19:@3378.4]
  assign _GEN_656 = 5'h10 == select_20 ? io_inData_16 : _GEN_655; // @[Switch.scala 33:19:@3378.4]
  assign _GEN_657 = 5'h11 == select_20 ? io_inData_17 : _GEN_656; // @[Switch.scala 33:19:@3378.4]
  assign _GEN_658 = 5'h12 == select_20 ? io_inData_18 : _GEN_657; // @[Switch.scala 33:19:@3378.4]
  assign _GEN_659 = 5'h13 == select_20 ? io_inData_19 : _GEN_658; // @[Switch.scala 33:19:@3378.4]
  assign _GEN_660 = 5'h14 == select_20 ? io_inData_20 : _GEN_659; // @[Switch.scala 33:19:@3378.4]
  assign _GEN_661 = 5'h15 == select_20 ? io_inData_21 : _GEN_660; // @[Switch.scala 33:19:@3378.4]
  assign _GEN_662 = 5'h16 == select_20 ? io_inData_22 : _GEN_661; // @[Switch.scala 33:19:@3378.4]
  assign _GEN_663 = 5'h17 == select_20 ? io_inData_23 : _GEN_662; // @[Switch.scala 33:19:@3378.4]
  assign _GEN_664 = 5'h18 == select_20 ? io_inData_24 : _GEN_663; // @[Switch.scala 33:19:@3378.4]
  assign _GEN_665 = 5'h19 == select_20 ? io_inData_25 : _GEN_664; // @[Switch.scala 33:19:@3378.4]
  assign _GEN_666 = 5'h1a == select_20 ? io_inData_26 : _GEN_665; // @[Switch.scala 33:19:@3378.4]
  assign _GEN_667 = 5'h1b == select_20 ? io_inData_27 : _GEN_666; // @[Switch.scala 33:19:@3378.4]
  assign _GEN_668 = 5'h1c == select_20 ? io_inData_28 : _GEN_667; // @[Switch.scala 33:19:@3378.4]
  assign _GEN_669 = 5'h1d == select_20 ? io_inData_29 : _GEN_668; // @[Switch.scala 33:19:@3378.4]
  assign _GEN_670 = 5'h1e == select_20 ? io_inData_30 : _GEN_669; // @[Switch.scala 33:19:@3378.4]
  assign _T_8783 = {valid_20_7,valid_20_6,valid_20_5,valid_20_4,valid_20_3,valid_20_2,valid_20_1,valid_20_0}; // @[Switch.scala 34:32:@3385.4]
  assign _T_8791 = {valid_20_15,valid_20_14,valid_20_13,valid_20_12,valid_20_11,valid_20_10,valid_20_9,valid_20_8,_T_8783}; // @[Switch.scala 34:32:@3393.4]
  assign _T_8798 = {valid_20_23,valid_20_22,valid_20_21,valid_20_20,valid_20_19,valid_20_18,valid_20_17,valid_20_16}; // @[Switch.scala 34:32:@3400.4]
  assign _T_8807 = {valid_20_31,valid_20_30,valid_20_29,valid_20_28,valid_20_27,valid_20_26,valid_20_25,valid_20_24,_T_8798,_T_8791}; // @[Switch.scala 34:32:@3409.4]
  assign _T_8811 = io_inAddr_0 == 5'h15; // @[Switch.scala 30:53:@3412.4]
  assign valid_21_0 = io_inValid_0 & _T_8811; // @[Switch.scala 30:36:@3413.4]
  assign _T_8814 = io_inAddr_1 == 5'h15; // @[Switch.scala 30:53:@3415.4]
  assign valid_21_1 = io_inValid_1 & _T_8814; // @[Switch.scala 30:36:@3416.4]
  assign _T_8817 = io_inAddr_2 == 5'h15; // @[Switch.scala 30:53:@3418.4]
  assign valid_21_2 = io_inValid_2 & _T_8817; // @[Switch.scala 30:36:@3419.4]
  assign _T_8820 = io_inAddr_3 == 5'h15; // @[Switch.scala 30:53:@3421.4]
  assign valid_21_3 = io_inValid_3 & _T_8820; // @[Switch.scala 30:36:@3422.4]
  assign _T_8823 = io_inAddr_4 == 5'h15; // @[Switch.scala 30:53:@3424.4]
  assign valid_21_4 = io_inValid_4 & _T_8823; // @[Switch.scala 30:36:@3425.4]
  assign _T_8826 = io_inAddr_5 == 5'h15; // @[Switch.scala 30:53:@3427.4]
  assign valid_21_5 = io_inValid_5 & _T_8826; // @[Switch.scala 30:36:@3428.4]
  assign _T_8829 = io_inAddr_6 == 5'h15; // @[Switch.scala 30:53:@3430.4]
  assign valid_21_6 = io_inValid_6 & _T_8829; // @[Switch.scala 30:36:@3431.4]
  assign _T_8832 = io_inAddr_7 == 5'h15; // @[Switch.scala 30:53:@3433.4]
  assign valid_21_7 = io_inValid_7 & _T_8832; // @[Switch.scala 30:36:@3434.4]
  assign _T_8835 = io_inAddr_8 == 5'h15; // @[Switch.scala 30:53:@3436.4]
  assign valid_21_8 = io_inValid_8 & _T_8835; // @[Switch.scala 30:36:@3437.4]
  assign _T_8838 = io_inAddr_9 == 5'h15; // @[Switch.scala 30:53:@3439.4]
  assign valid_21_9 = io_inValid_9 & _T_8838; // @[Switch.scala 30:36:@3440.4]
  assign _T_8841 = io_inAddr_10 == 5'h15; // @[Switch.scala 30:53:@3442.4]
  assign valid_21_10 = io_inValid_10 & _T_8841; // @[Switch.scala 30:36:@3443.4]
  assign _T_8844 = io_inAddr_11 == 5'h15; // @[Switch.scala 30:53:@3445.4]
  assign valid_21_11 = io_inValid_11 & _T_8844; // @[Switch.scala 30:36:@3446.4]
  assign _T_8847 = io_inAddr_12 == 5'h15; // @[Switch.scala 30:53:@3448.4]
  assign valid_21_12 = io_inValid_12 & _T_8847; // @[Switch.scala 30:36:@3449.4]
  assign _T_8850 = io_inAddr_13 == 5'h15; // @[Switch.scala 30:53:@3451.4]
  assign valid_21_13 = io_inValid_13 & _T_8850; // @[Switch.scala 30:36:@3452.4]
  assign _T_8853 = io_inAddr_14 == 5'h15; // @[Switch.scala 30:53:@3454.4]
  assign valid_21_14 = io_inValid_14 & _T_8853; // @[Switch.scala 30:36:@3455.4]
  assign _T_8856 = io_inAddr_15 == 5'h15; // @[Switch.scala 30:53:@3457.4]
  assign valid_21_15 = io_inValid_15 & _T_8856; // @[Switch.scala 30:36:@3458.4]
  assign _T_8859 = io_inAddr_16 == 5'h15; // @[Switch.scala 30:53:@3460.4]
  assign valid_21_16 = io_inValid_16 & _T_8859; // @[Switch.scala 30:36:@3461.4]
  assign _T_8862 = io_inAddr_17 == 5'h15; // @[Switch.scala 30:53:@3463.4]
  assign valid_21_17 = io_inValid_17 & _T_8862; // @[Switch.scala 30:36:@3464.4]
  assign _T_8865 = io_inAddr_18 == 5'h15; // @[Switch.scala 30:53:@3466.4]
  assign valid_21_18 = io_inValid_18 & _T_8865; // @[Switch.scala 30:36:@3467.4]
  assign _T_8868 = io_inAddr_19 == 5'h15; // @[Switch.scala 30:53:@3469.4]
  assign valid_21_19 = io_inValid_19 & _T_8868; // @[Switch.scala 30:36:@3470.4]
  assign _T_8871 = io_inAddr_20 == 5'h15; // @[Switch.scala 30:53:@3472.4]
  assign valid_21_20 = io_inValid_20 & _T_8871; // @[Switch.scala 30:36:@3473.4]
  assign _T_8874 = io_inAddr_21 == 5'h15; // @[Switch.scala 30:53:@3475.4]
  assign valid_21_21 = io_inValid_21 & _T_8874; // @[Switch.scala 30:36:@3476.4]
  assign _T_8877 = io_inAddr_22 == 5'h15; // @[Switch.scala 30:53:@3478.4]
  assign valid_21_22 = io_inValid_22 & _T_8877; // @[Switch.scala 30:36:@3479.4]
  assign _T_8880 = io_inAddr_23 == 5'h15; // @[Switch.scala 30:53:@3481.4]
  assign valid_21_23 = io_inValid_23 & _T_8880; // @[Switch.scala 30:36:@3482.4]
  assign _T_8883 = io_inAddr_24 == 5'h15; // @[Switch.scala 30:53:@3484.4]
  assign valid_21_24 = io_inValid_24 & _T_8883; // @[Switch.scala 30:36:@3485.4]
  assign _T_8886 = io_inAddr_25 == 5'h15; // @[Switch.scala 30:53:@3487.4]
  assign valid_21_25 = io_inValid_25 & _T_8886; // @[Switch.scala 30:36:@3488.4]
  assign _T_8889 = io_inAddr_26 == 5'h15; // @[Switch.scala 30:53:@3490.4]
  assign valid_21_26 = io_inValid_26 & _T_8889; // @[Switch.scala 30:36:@3491.4]
  assign _T_8892 = io_inAddr_27 == 5'h15; // @[Switch.scala 30:53:@3493.4]
  assign valid_21_27 = io_inValid_27 & _T_8892; // @[Switch.scala 30:36:@3494.4]
  assign _T_8895 = io_inAddr_28 == 5'h15; // @[Switch.scala 30:53:@3496.4]
  assign valid_21_28 = io_inValid_28 & _T_8895; // @[Switch.scala 30:36:@3497.4]
  assign _T_8898 = io_inAddr_29 == 5'h15; // @[Switch.scala 30:53:@3499.4]
  assign valid_21_29 = io_inValid_29 & _T_8898; // @[Switch.scala 30:36:@3500.4]
  assign _T_8901 = io_inAddr_30 == 5'h15; // @[Switch.scala 30:53:@3502.4]
  assign valid_21_30 = io_inValid_30 & _T_8901; // @[Switch.scala 30:36:@3503.4]
  assign _T_8904 = io_inAddr_31 == 5'h15; // @[Switch.scala 30:53:@3505.4]
  assign valid_21_31 = io_inValid_31 & _T_8904; // @[Switch.scala 30:36:@3506.4]
  assign _T_8938 = valid_21_30 ? 5'h1e : 5'h1f; // @[Mux.scala 31:69:@3508.4]
  assign _T_8939 = valid_21_29 ? 5'h1d : _T_8938; // @[Mux.scala 31:69:@3509.4]
  assign _T_8940 = valid_21_28 ? 5'h1c : _T_8939; // @[Mux.scala 31:69:@3510.4]
  assign _T_8941 = valid_21_27 ? 5'h1b : _T_8940; // @[Mux.scala 31:69:@3511.4]
  assign _T_8942 = valid_21_26 ? 5'h1a : _T_8941; // @[Mux.scala 31:69:@3512.4]
  assign _T_8943 = valid_21_25 ? 5'h19 : _T_8942; // @[Mux.scala 31:69:@3513.4]
  assign _T_8944 = valid_21_24 ? 5'h18 : _T_8943; // @[Mux.scala 31:69:@3514.4]
  assign _T_8945 = valid_21_23 ? 5'h17 : _T_8944; // @[Mux.scala 31:69:@3515.4]
  assign _T_8946 = valid_21_22 ? 5'h16 : _T_8945; // @[Mux.scala 31:69:@3516.4]
  assign _T_8947 = valid_21_21 ? 5'h15 : _T_8946; // @[Mux.scala 31:69:@3517.4]
  assign _T_8948 = valid_21_20 ? 5'h14 : _T_8947; // @[Mux.scala 31:69:@3518.4]
  assign _T_8949 = valid_21_19 ? 5'h13 : _T_8948; // @[Mux.scala 31:69:@3519.4]
  assign _T_8950 = valid_21_18 ? 5'h12 : _T_8949; // @[Mux.scala 31:69:@3520.4]
  assign _T_8951 = valid_21_17 ? 5'h11 : _T_8950; // @[Mux.scala 31:69:@3521.4]
  assign _T_8952 = valid_21_16 ? 5'h10 : _T_8951; // @[Mux.scala 31:69:@3522.4]
  assign _T_8953 = valid_21_15 ? 5'hf : _T_8952; // @[Mux.scala 31:69:@3523.4]
  assign _T_8954 = valid_21_14 ? 5'he : _T_8953; // @[Mux.scala 31:69:@3524.4]
  assign _T_8955 = valid_21_13 ? 5'hd : _T_8954; // @[Mux.scala 31:69:@3525.4]
  assign _T_8956 = valid_21_12 ? 5'hc : _T_8955; // @[Mux.scala 31:69:@3526.4]
  assign _T_8957 = valid_21_11 ? 5'hb : _T_8956; // @[Mux.scala 31:69:@3527.4]
  assign _T_8958 = valid_21_10 ? 5'ha : _T_8957; // @[Mux.scala 31:69:@3528.4]
  assign _T_8959 = valid_21_9 ? 5'h9 : _T_8958; // @[Mux.scala 31:69:@3529.4]
  assign _T_8960 = valid_21_8 ? 5'h8 : _T_8959; // @[Mux.scala 31:69:@3530.4]
  assign _T_8961 = valid_21_7 ? 5'h7 : _T_8960; // @[Mux.scala 31:69:@3531.4]
  assign _T_8962 = valid_21_6 ? 5'h6 : _T_8961; // @[Mux.scala 31:69:@3532.4]
  assign _T_8963 = valid_21_5 ? 5'h5 : _T_8962; // @[Mux.scala 31:69:@3533.4]
  assign _T_8964 = valid_21_4 ? 5'h4 : _T_8963; // @[Mux.scala 31:69:@3534.4]
  assign _T_8965 = valid_21_3 ? 5'h3 : _T_8964; // @[Mux.scala 31:69:@3535.4]
  assign _T_8966 = valid_21_2 ? 5'h2 : _T_8965; // @[Mux.scala 31:69:@3536.4]
  assign _T_8967 = valid_21_1 ? 5'h1 : _T_8966; // @[Mux.scala 31:69:@3537.4]
  assign select_21 = valid_21_0 ? 5'h0 : _T_8967; // @[Mux.scala 31:69:@3538.4]
  assign _GEN_673 = 5'h1 == select_21 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@3540.4]
  assign _GEN_674 = 5'h2 == select_21 ? io_inData_2 : _GEN_673; // @[Switch.scala 33:19:@3540.4]
  assign _GEN_675 = 5'h3 == select_21 ? io_inData_3 : _GEN_674; // @[Switch.scala 33:19:@3540.4]
  assign _GEN_676 = 5'h4 == select_21 ? io_inData_4 : _GEN_675; // @[Switch.scala 33:19:@3540.4]
  assign _GEN_677 = 5'h5 == select_21 ? io_inData_5 : _GEN_676; // @[Switch.scala 33:19:@3540.4]
  assign _GEN_678 = 5'h6 == select_21 ? io_inData_6 : _GEN_677; // @[Switch.scala 33:19:@3540.4]
  assign _GEN_679 = 5'h7 == select_21 ? io_inData_7 : _GEN_678; // @[Switch.scala 33:19:@3540.4]
  assign _GEN_680 = 5'h8 == select_21 ? io_inData_8 : _GEN_679; // @[Switch.scala 33:19:@3540.4]
  assign _GEN_681 = 5'h9 == select_21 ? io_inData_9 : _GEN_680; // @[Switch.scala 33:19:@3540.4]
  assign _GEN_682 = 5'ha == select_21 ? io_inData_10 : _GEN_681; // @[Switch.scala 33:19:@3540.4]
  assign _GEN_683 = 5'hb == select_21 ? io_inData_11 : _GEN_682; // @[Switch.scala 33:19:@3540.4]
  assign _GEN_684 = 5'hc == select_21 ? io_inData_12 : _GEN_683; // @[Switch.scala 33:19:@3540.4]
  assign _GEN_685 = 5'hd == select_21 ? io_inData_13 : _GEN_684; // @[Switch.scala 33:19:@3540.4]
  assign _GEN_686 = 5'he == select_21 ? io_inData_14 : _GEN_685; // @[Switch.scala 33:19:@3540.4]
  assign _GEN_687 = 5'hf == select_21 ? io_inData_15 : _GEN_686; // @[Switch.scala 33:19:@3540.4]
  assign _GEN_688 = 5'h10 == select_21 ? io_inData_16 : _GEN_687; // @[Switch.scala 33:19:@3540.4]
  assign _GEN_689 = 5'h11 == select_21 ? io_inData_17 : _GEN_688; // @[Switch.scala 33:19:@3540.4]
  assign _GEN_690 = 5'h12 == select_21 ? io_inData_18 : _GEN_689; // @[Switch.scala 33:19:@3540.4]
  assign _GEN_691 = 5'h13 == select_21 ? io_inData_19 : _GEN_690; // @[Switch.scala 33:19:@3540.4]
  assign _GEN_692 = 5'h14 == select_21 ? io_inData_20 : _GEN_691; // @[Switch.scala 33:19:@3540.4]
  assign _GEN_693 = 5'h15 == select_21 ? io_inData_21 : _GEN_692; // @[Switch.scala 33:19:@3540.4]
  assign _GEN_694 = 5'h16 == select_21 ? io_inData_22 : _GEN_693; // @[Switch.scala 33:19:@3540.4]
  assign _GEN_695 = 5'h17 == select_21 ? io_inData_23 : _GEN_694; // @[Switch.scala 33:19:@3540.4]
  assign _GEN_696 = 5'h18 == select_21 ? io_inData_24 : _GEN_695; // @[Switch.scala 33:19:@3540.4]
  assign _GEN_697 = 5'h19 == select_21 ? io_inData_25 : _GEN_696; // @[Switch.scala 33:19:@3540.4]
  assign _GEN_698 = 5'h1a == select_21 ? io_inData_26 : _GEN_697; // @[Switch.scala 33:19:@3540.4]
  assign _GEN_699 = 5'h1b == select_21 ? io_inData_27 : _GEN_698; // @[Switch.scala 33:19:@3540.4]
  assign _GEN_700 = 5'h1c == select_21 ? io_inData_28 : _GEN_699; // @[Switch.scala 33:19:@3540.4]
  assign _GEN_701 = 5'h1d == select_21 ? io_inData_29 : _GEN_700; // @[Switch.scala 33:19:@3540.4]
  assign _GEN_702 = 5'h1e == select_21 ? io_inData_30 : _GEN_701; // @[Switch.scala 33:19:@3540.4]
  assign _T_8976 = {valid_21_7,valid_21_6,valid_21_5,valid_21_4,valid_21_3,valid_21_2,valid_21_1,valid_21_0}; // @[Switch.scala 34:32:@3547.4]
  assign _T_8984 = {valid_21_15,valid_21_14,valid_21_13,valid_21_12,valid_21_11,valid_21_10,valid_21_9,valid_21_8,_T_8976}; // @[Switch.scala 34:32:@3555.4]
  assign _T_8991 = {valid_21_23,valid_21_22,valid_21_21,valid_21_20,valid_21_19,valid_21_18,valid_21_17,valid_21_16}; // @[Switch.scala 34:32:@3562.4]
  assign _T_9000 = {valid_21_31,valid_21_30,valid_21_29,valid_21_28,valid_21_27,valid_21_26,valid_21_25,valid_21_24,_T_8991,_T_8984}; // @[Switch.scala 34:32:@3571.4]
  assign _T_9004 = io_inAddr_0 == 5'h16; // @[Switch.scala 30:53:@3574.4]
  assign valid_22_0 = io_inValid_0 & _T_9004; // @[Switch.scala 30:36:@3575.4]
  assign _T_9007 = io_inAddr_1 == 5'h16; // @[Switch.scala 30:53:@3577.4]
  assign valid_22_1 = io_inValid_1 & _T_9007; // @[Switch.scala 30:36:@3578.4]
  assign _T_9010 = io_inAddr_2 == 5'h16; // @[Switch.scala 30:53:@3580.4]
  assign valid_22_2 = io_inValid_2 & _T_9010; // @[Switch.scala 30:36:@3581.4]
  assign _T_9013 = io_inAddr_3 == 5'h16; // @[Switch.scala 30:53:@3583.4]
  assign valid_22_3 = io_inValid_3 & _T_9013; // @[Switch.scala 30:36:@3584.4]
  assign _T_9016 = io_inAddr_4 == 5'h16; // @[Switch.scala 30:53:@3586.4]
  assign valid_22_4 = io_inValid_4 & _T_9016; // @[Switch.scala 30:36:@3587.4]
  assign _T_9019 = io_inAddr_5 == 5'h16; // @[Switch.scala 30:53:@3589.4]
  assign valid_22_5 = io_inValid_5 & _T_9019; // @[Switch.scala 30:36:@3590.4]
  assign _T_9022 = io_inAddr_6 == 5'h16; // @[Switch.scala 30:53:@3592.4]
  assign valid_22_6 = io_inValid_6 & _T_9022; // @[Switch.scala 30:36:@3593.4]
  assign _T_9025 = io_inAddr_7 == 5'h16; // @[Switch.scala 30:53:@3595.4]
  assign valid_22_7 = io_inValid_7 & _T_9025; // @[Switch.scala 30:36:@3596.4]
  assign _T_9028 = io_inAddr_8 == 5'h16; // @[Switch.scala 30:53:@3598.4]
  assign valid_22_8 = io_inValid_8 & _T_9028; // @[Switch.scala 30:36:@3599.4]
  assign _T_9031 = io_inAddr_9 == 5'h16; // @[Switch.scala 30:53:@3601.4]
  assign valid_22_9 = io_inValid_9 & _T_9031; // @[Switch.scala 30:36:@3602.4]
  assign _T_9034 = io_inAddr_10 == 5'h16; // @[Switch.scala 30:53:@3604.4]
  assign valid_22_10 = io_inValid_10 & _T_9034; // @[Switch.scala 30:36:@3605.4]
  assign _T_9037 = io_inAddr_11 == 5'h16; // @[Switch.scala 30:53:@3607.4]
  assign valid_22_11 = io_inValid_11 & _T_9037; // @[Switch.scala 30:36:@3608.4]
  assign _T_9040 = io_inAddr_12 == 5'h16; // @[Switch.scala 30:53:@3610.4]
  assign valid_22_12 = io_inValid_12 & _T_9040; // @[Switch.scala 30:36:@3611.4]
  assign _T_9043 = io_inAddr_13 == 5'h16; // @[Switch.scala 30:53:@3613.4]
  assign valid_22_13 = io_inValid_13 & _T_9043; // @[Switch.scala 30:36:@3614.4]
  assign _T_9046 = io_inAddr_14 == 5'h16; // @[Switch.scala 30:53:@3616.4]
  assign valid_22_14 = io_inValid_14 & _T_9046; // @[Switch.scala 30:36:@3617.4]
  assign _T_9049 = io_inAddr_15 == 5'h16; // @[Switch.scala 30:53:@3619.4]
  assign valid_22_15 = io_inValid_15 & _T_9049; // @[Switch.scala 30:36:@3620.4]
  assign _T_9052 = io_inAddr_16 == 5'h16; // @[Switch.scala 30:53:@3622.4]
  assign valid_22_16 = io_inValid_16 & _T_9052; // @[Switch.scala 30:36:@3623.4]
  assign _T_9055 = io_inAddr_17 == 5'h16; // @[Switch.scala 30:53:@3625.4]
  assign valid_22_17 = io_inValid_17 & _T_9055; // @[Switch.scala 30:36:@3626.4]
  assign _T_9058 = io_inAddr_18 == 5'h16; // @[Switch.scala 30:53:@3628.4]
  assign valid_22_18 = io_inValid_18 & _T_9058; // @[Switch.scala 30:36:@3629.4]
  assign _T_9061 = io_inAddr_19 == 5'h16; // @[Switch.scala 30:53:@3631.4]
  assign valid_22_19 = io_inValid_19 & _T_9061; // @[Switch.scala 30:36:@3632.4]
  assign _T_9064 = io_inAddr_20 == 5'h16; // @[Switch.scala 30:53:@3634.4]
  assign valid_22_20 = io_inValid_20 & _T_9064; // @[Switch.scala 30:36:@3635.4]
  assign _T_9067 = io_inAddr_21 == 5'h16; // @[Switch.scala 30:53:@3637.4]
  assign valid_22_21 = io_inValid_21 & _T_9067; // @[Switch.scala 30:36:@3638.4]
  assign _T_9070 = io_inAddr_22 == 5'h16; // @[Switch.scala 30:53:@3640.4]
  assign valid_22_22 = io_inValid_22 & _T_9070; // @[Switch.scala 30:36:@3641.4]
  assign _T_9073 = io_inAddr_23 == 5'h16; // @[Switch.scala 30:53:@3643.4]
  assign valid_22_23 = io_inValid_23 & _T_9073; // @[Switch.scala 30:36:@3644.4]
  assign _T_9076 = io_inAddr_24 == 5'h16; // @[Switch.scala 30:53:@3646.4]
  assign valid_22_24 = io_inValid_24 & _T_9076; // @[Switch.scala 30:36:@3647.4]
  assign _T_9079 = io_inAddr_25 == 5'h16; // @[Switch.scala 30:53:@3649.4]
  assign valid_22_25 = io_inValid_25 & _T_9079; // @[Switch.scala 30:36:@3650.4]
  assign _T_9082 = io_inAddr_26 == 5'h16; // @[Switch.scala 30:53:@3652.4]
  assign valid_22_26 = io_inValid_26 & _T_9082; // @[Switch.scala 30:36:@3653.4]
  assign _T_9085 = io_inAddr_27 == 5'h16; // @[Switch.scala 30:53:@3655.4]
  assign valid_22_27 = io_inValid_27 & _T_9085; // @[Switch.scala 30:36:@3656.4]
  assign _T_9088 = io_inAddr_28 == 5'h16; // @[Switch.scala 30:53:@3658.4]
  assign valid_22_28 = io_inValid_28 & _T_9088; // @[Switch.scala 30:36:@3659.4]
  assign _T_9091 = io_inAddr_29 == 5'h16; // @[Switch.scala 30:53:@3661.4]
  assign valid_22_29 = io_inValid_29 & _T_9091; // @[Switch.scala 30:36:@3662.4]
  assign _T_9094 = io_inAddr_30 == 5'h16; // @[Switch.scala 30:53:@3664.4]
  assign valid_22_30 = io_inValid_30 & _T_9094; // @[Switch.scala 30:36:@3665.4]
  assign _T_9097 = io_inAddr_31 == 5'h16; // @[Switch.scala 30:53:@3667.4]
  assign valid_22_31 = io_inValid_31 & _T_9097; // @[Switch.scala 30:36:@3668.4]
  assign _T_9131 = valid_22_30 ? 5'h1e : 5'h1f; // @[Mux.scala 31:69:@3670.4]
  assign _T_9132 = valid_22_29 ? 5'h1d : _T_9131; // @[Mux.scala 31:69:@3671.4]
  assign _T_9133 = valid_22_28 ? 5'h1c : _T_9132; // @[Mux.scala 31:69:@3672.4]
  assign _T_9134 = valid_22_27 ? 5'h1b : _T_9133; // @[Mux.scala 31:69:@3673.4]
  assign _T_9135 = valid_22_26 ? 5'h1a : _T_9134; // @[Mux.scala 31:69:@3674.4]
  assign _T_9136 = valid_22_25 ? 5'h19 : _T_9135; // @[Mux.scala 31:69:@3675.4]
  assign _T_9137 = valid_22_24 ? 5'h18 : _T_9136; // @[Mux.scala 31:69:@3676.4]
  assign _T_9138 = valid_22_23 ? 5'h17 : _T_9137; // @[Mux.scala 31:69:@3677.4]
  assign _T_9139 = valid_22_22 ? 5'h16 : _T_9138; // @[Mux.scala 31:69:@3678.4]
  assign _T_9140 = valid_22_21 ? 5'h15 : _T_9139; // @[Mux.scala 31:69:@3679.4]
  assign _T_9141 = valid_22_20 ? 5'h14 : _T_9140; // @[Mux.scala 31:69:@3680.4]
  assign _T_9142 = valid_22_19 ? 5'h13 : _T_9141; // @[Mux.scala 31:69:@3681.4]
  assign _T_9143 = valid_22_18 ? 5'h12 : _T_9142; // @[Mux.scala 31:69:@3682.4]
  assign _T_9144 = valid_22_17 ? 5'h11 : _T_9143; // @[Mux.scala 31:69:@3683.4]
  assign _T_9145 = valid_22_16 ? 5'h10 : _T_9144; // @[Mux.scala 31:69:@3684.4]
  assign _T_9146 = valid_22_15 ? 5'hf : _T_9145; // @[Mux.scala 31:69:@3685.4]
  assign _T_9147 = valid_22_14 ? 5'he : _T_9146; // @[Mux.scala 31:69:@3686.4]
  assign _T_9148 = valid_22_13 ? 5'hd : _T_9147; // @[Mux.scala 31:69:@3687.4]
  assign _T_9149 = valid_22_12 ? 5'hc : _T_9148; // @[Mux.scala 31:69:@3688.4]
  assign _T_9150 = valid_22_11 ? 5'hb : _T_9149; // @[Mux.scala 31:69:@3689.4]
  assign _T_9151 = valid_22_10 ? 5'ha : _T_9150; // @[Mux.scala 31:69:@3690.4]
  assign _T_9152 = valid_22_9 ? 5'h9 : _T_9151; // @[Mux.scala 31:69:@3691.4]
  assign _T_9153 = valid_22_8 ? 5'h8 : _T_9152; // @[Mux.scala 31:69:@3692.4]
  assign _T_9154 = valid_22_7 ? 5'h7 : _T_9153; // @[Mux.scala 31:69:@3693.4]
  assign _T_9155 = valid_22_6 ? 5'h6 : _T_9154; // @[Mux.scala 31:69:@3694.4]
  assign _T_9156 = valid_22_5 ? 5'h5 : _T_9155; // @[Mux.scala 31:69:@3695.4]
  assign _T_9157 = valid_22_4 ? 5'h4 : _T_9156; // @[Mux.scala 31:69:@3696.4]
  assign _T_9158 = valid_22_3 ? 5'h3 : _T_9157; // @[Mux.scala 31:69:@3697.4]
  assign _T_9159 = valid_22_2 ? 5'h2 : _T_9158; // @[Mux.scala 31:69:@3698.4]
  assign _T_9160 = valid_22_1 ? 5'h1 : _T_9159; // @[Mux.scala 31:69:@3699.4]
  assign select_22 = valid_22_0 ? 5'h0 : _T_9160; // @[Mux.scala 31:69:@3700.4]
  assign _GEN_705 = 5'h1 == select_22 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@3702.4]
  assign _GEN_706 = 5'h2 == select_22 ? io_inData_2 : _GEN_705; // @[Switch.scala 33:19:@3702.4]
  assign _GEN_707 = 5'h3 == select_22 ? io_inData_3 : _GEN_706; // @[Switch.scala 33:19:@3702.4]
  assign _GEN_708 = 5'h4 == select_22 ? io_inData_4 : _GEN_707; // @[Switch.scala 33:19:@3702.4]
  assign _GEN_709 = 5'h5 == select_22 ? io_inData_5 : _GEN_708; // @[Switch.scala 33:19:@3702.4]
  assign _GEN_710 = 5'h6 == select_22 ? io_inData_6 : _GEN_709; // @[Switch.scala 33:19:@3702.4]
  assign _GEN_711 = 5'h7 == select_22 ? io_inData_7 : _GEN_710; // @[Switch.scala 33:19:@3702.4]
  assign _GEN_712 = 5'h8 == select_22 ? io_inData_8 : _GEN_711; // @[Switch.scala 33:19:@3702.4]
  assign _GEN_713 = 5'h9 == select_22 ? io_inData_9 : _GEN_712; // @[Switch.scala 33:19:@3702.4]
  assign _GEN_714 = 5'ha == select_22 ? io_inData_10 : _GEN_713; // @[Switch.scala 33:19:@3702.4]
  assign _GEN_715 = 5'hb == select_22 ? io_inData_11 : _GEN_714; // @[Switch.scala 33:19:@3702.4]
  assign _GEN_716 = 5'hc == select_22 ? io_inData_12 : _GEN_715; // @[Switch.scala 33:19:@3702.4]
  assign _GEN_717 = 5'hd == select_22 ? io_inData_13 : _GEN_716; // @[Switch.scala 33:19:@3702.4]
  assign _GEN_718 = 5'he == select_22 ? io_inData_14 : _GEN_717; // @[Switch.scala 33:19:@3702.4]
  assign _GEN_719 = 5'hf == select_22 ? io_inData_15 : _GEN_718; // @[Switch.scala 33:19:@3702.4]
  assign _GEN_720 = 5'h10 == select_22 ? io_inData_16 : _GEN_719; // @[Switch.scala 33:19:@3702.4]
  assign _GEN_721 = 5'h11 == select_22 ? io_inData_17 : _GEN_720; // @[Switch.scala 33:19:@3702.4]
  assign _GEN_722 = 5'h12 == select_22 ? io_inData_18 : _GEN_721; // @[Switch.scala 33:19:@3702.4]
  assign _GEN_723 = 5'h13 == select_22 ? io_inData_19 : _GEN_722; // @[Switch.scala 33:19:@3702.4]
  assign _GEN_724 = 5'h14 == select_22 ? io_inData_20 : _GEN_723; // @[Switch.scala 33:19:@3702.4]
  assign _GEN_725 = 5'h15 == select_22 ? io_inData_21 : _GEN_724; // @[Switch.scala 33:19:@3702.4]
  assign _GEN_726 = 5'h16 == select_22 ? io_inData_22 : _GEN_725; // @[Switch.scala 33:19:@3702.4]
  assign _GEN_727 = 5'h17 == select_22 ? io_inData_23 : _GEN_726; // @[Switch.scala 33:19:@3702.4]
  assign _GEN_728 = 5'h18 == select_22 ? io_inData_24 : _GEN_727; // @[Switch.scala 33:19:@3702.4]
  assign _GEN_729 = 5'h19 == select_22 ? io_inData_25 : _GEN_728; // @[Switch.scala 33:19:@3702.4]
  assign _GEN_730 = 5'h1a == select_22 ? io_inData_26 : _GEN_729; // @[Switch.scala 33:19:@3702.4]
  assign _GEN_731 = 5'h1b == select_22 ? io_inData_27 : _GEN_730; // @[Switch.scala 33:19:@3702.4]
  assign _GEN_732 = 5'h1c == select_22 ? io_inData_28 : _GEN_731; // @[Switch.scala 33:19:@3702.4]
  assign _GEN_733 = 5'h1d == select_22 ? io_inData_29 : _GEN_732; // @[Switch.scala 33:19:@3702.4]
  assign _GEN_734 = 5'h1e == select_22 ? io_inData_30 : _GEN_733; // @[Switch.scala 33:19:@3702.4]
  assign _T_9169 = {valid_22_7,valid_22_6,valid_22_5,valid_22_4,valid_22_3,valid_22_2,valid_22_1,valid_22_0}; // @[Switch.scala 34:32:@3709.4]
  assign _T_9177 = {valid_22_15,valid_22_14,valid_22_13,valid_22_12,valid_22_11,valid_22_10,valid_22_9,valid_22_8,_T_9169}; // @[Switch.scala 34:32:@3717.4]
  assign _T_9184 = {valid_22_23,valid_22_22,valid_22_21,valid_22_20,valid_22_19,valid_22_18,valid_22_17,valid_22_16}; // @[Switch.scala 34:32:@3724.4]
  assign _T_9193 = {valid_22_31,valid_22_30,valid_22_29,valid_22_28,valid_22_27,valid_22_26,valid_22_25,valid_22_24,_T_9184,_T_9177}; // @[Switch.scala 34:32:@3733.4]
  assign _T_9197 = io_inAddr_0 == 5'h17; // @[Switch.scala 30:53:@3736.4]
  assign valid_23_0 = io_inValid_0 & _T_9197; // @[Switch.scala 30:36:@3737.4]
  assign _T_9200 = io_inAddr_1 == 5'h17; // @[Switch.scala 30:53:@3739.4]
  assign valid_23_1 = io_inValid_1 & _T_9200; // @[Switch.scala 30:36:@3740.4]
  assign _T_9203 = io_inAddr_2 == 5'h17; // @[Switch.scala 30:53:@3742.4]
  assign valid_23_2 = io_inValid_2 & _T_9203; // @[Switch.scala 30:36:@3743.4]
  assign _T_9206 = io_inAddr_3 == 5'h17; // @[Switch.scala 30:53:@3745.4]
  assign valid_23_3 = io_inValid_3 & _T_9206; // @[Switch.scala 30:36:@3746.4]
  assign _T_9209 = io_inAddr_4 == 5'h17; // @[Switch.scala 30:53:@3748.4]
  assign valid_23_4 = io_inValid_4 & _T_9209; // @[Switch.scala 30:36:@3749.4]
  assign _T_9212 = io_inAddr_5 == 5'h17; // @[Switch.scala 30:53:@3751.4]
  assign valid_23_5 = io_inValid_5 & _T_9212; // @[Switch.scala 30:36:@3752.4]
  assign _T_9215 = io_inAddr_6 == 5'h17; // @[Switch.scala 30:53:@3754.4]
  assign valid_23_6 = io_inValid_6 & _T_9215; // @[Switch.scala 30:36:@3755.4]
  assign _T_9218 = io_inAddr_7 == 5'h17; // @[Switch.scala 30:53:@3757.4]
  assign valid_23_7 = io_inValid_7 & _T_9218; // @[Switch.scala 30:36:@3758.4]
  assign _T_9221 = io_inAddr_8 == 5'h17; // @[Switch.scala 30:53:@3760.4]
  assign valid_23_8 = io_inValid_8 & _T_9221; // @[Switch.scala 30:36:@3761.4]
  assign _T_9224 = io_inAddr_9 == 5'h17; // @[Switch.scala 30:53:@3763.4]
  assign valid_23_9 = io_inValid_9 & _T_9224; // @[Switch.scala 30:36:@3764.4]
  assign _T_9227 = io_inAddr_10 == 5'h17; // @[Switch.scala 30:53:@3766.4]
  assign valid_23_10 = io_inValid_10 & _T_9227; // @[Switch.scala 30:36:@3767.4]
  assign _T_9230 = io_inAddr_11 == 5'h17; // @[Switch.scala 30:53:@3769.4]
  assign valid_23_11 = io_inValid_11 & _T_9230; // @[Switch.scala 30:36:@3770.4]
  assign _T_9233 = io_inAddr_12 == 5'h17; // @[Switch.scala 30:53:@3772.4]
  assign valid_23_12 = io_inValid_12 & _T_9233; // @[Switch.scala 30:36:@3773.4]
  assign _T_9236 = io_inAddr_13 == 5'h17; // @[Switch.scala 30:53:@3775.4]
  assign valid_23_13 = io_inValid_13 & _T_9236; // @[Switch.scala 30:36:@3776.4]
  assign _T_9239 = io_inAddr_14 == 5'h17; // @[Switch.scala 30:53:@3778.4]
  assign valid_23_14 = io_inValid_14 & _T_9239; // @[Switch.scala 30:36:@3779.4]
  assign _T_9242 = io_inAddr_15 == 5'h17; // @[Switch.scala 30:53:@3781.4]
  assign valid_23_15 = io_inValid_15 & _T_9242; // @[Switch.scala 30:36:@3782.4]
  assign _T_9245 = io_inAddr_16 == 5'h17; // @[Switch.scala 30:53:@3784.4]
  assign valid_23_16 = io_inValid_16 & _T_9245; // @[Switch.scala 30:36:@3785.4]
  assign _T_9248 = io_inAddr_17 == 5'h17; // @[Switch.scala 30:53:@3787.4]
  assign valid_23_17 = io_inValid_17 & _T_9248; // @[Switch.scala 30:36:@3788.4]
  assign _T_9251 = io_inAddr_18 == 5'h17; // @[Switch.scala 30:53:@3790.4]
  assign valid_23_18 = io_inValid_18 & _T_9251; // @[Switch.scala 30:36:@3791.4]
  assign _T_9254 = io_inAddr_19 == 5'h17; // @[Switch.scala 30:53:@3793.4]
  assign valid_23_19 = io_inValid_19 & _T_9254; // @[Switch.scala 30:36:@3794.4]
  assign _T_9257 = io_inAddr_20 == 5'h17; // @[Switch.scala 30:53:@3796.4]
  assign valid_23_20 = io_inValid_20 & _T_9257; // @[Switch.scala 30:36:@3797.4]
  assign _T_9260 = io_inAddr_21 == 5'h17; // @[Switch.scala 30:53:@3799.4]
  assign valid_23_21 = io_inValid_21 & _T_9260; // @[Switch.scala 30:36:@3800.4]
  assign _T_9263 = io_inAddr_22 == 5'h17; // @[Switch.scala 30:53:@3802.4]
  assign valid_23_22 = io_inValid_22 & _T_9263; // @[Switch.scala 30:36:@3803.4]
  assign _T_9266 = io_inAddr_23 == 5'h17; // @[Switch.scala 30:53:@3805.4]
  assign valid_23_23 = io_inValid_23 & _T_9266; // @[Switch.scala 30:36:@3806.4]
  assign _T_9269 = io_inAddr_24 == 5'h17; // @[Switch.scala 30:53:@3808.4]
  assign valid_23_24 = io_inValid_24 & _T_9269; // @[Switch.scala 30:36:@3809.4]
  assign _T_9272 = io_inAddr_25 == 5'h17; // @[Switch.scala 30:53:@3811.4]
  assign valid_23_25 = io_inValid_25 & _T_9272; // @[Switch.scala 30:36:@3812.4]
  assign _T_9275 = io_inAddr_26 == 5'h17; // @[Switch.scala 30:53:@3814.4]
  assign valid_23_26 = io_inValid_26 & _T_9275; // @[Switch.scala 30:36:@3815.4]
  assign _T_9278 = io_inAddr_27 == 5'h17; // @[Switch.scala 30:53:@3817.4]
  assign valid_23_27 = io_inValid_27 & _T_9278; // @[Switch.scala 30:36:@3818.4]
  assign _T_9281 = io_inAddr_28 == 5'h17; // @[Switch.scala 30:53:@3820.4]
  assign valid_23_28 = io_inValid_28 & _T_9281; // @[Switch.scala 30:36:@3821.4]
  assign _T_9284 = io_inAddr_29 == 5'h17; // @[Switch.scala 30:53:@3823.4]
  assign valid_23_29 = io_inValid_29 & _T_9284; // @[Switch.scala 30:36:@3824.4]
  assign _T_9287 = io_inAddr_30 == 5'h17; // @[Switch.scala 30:53:@3826.4]
  assign valid_23_30 = io_inValid_30 & _T_9287; // @[Switch.scala 30:36:@3827.4]
  assign _T_9290 = io_inAddr_31 == 5'h17; // @[Switch.scala 30:53:@3829.4]
  assign valid_23_31 = io_inValid_31 & _T_9290; // @[Switch.scala 30:36:@3830.4]
  assign _T_9324 = valid_23_30 ? 5'h1e : 5'h1f; // @[Mux.scala 31:69:@3832.4]
  assign _T_9325 = valid_23_29 ? 5'h1d : _T_9324; // @[Mux.scala 31:69:@3833.4]
  assign _T_9326 = valid_23_28 ? 5'h1c : _T_9325; // @[Mux.scala 31:69:@3834.4]
  assign _T_9327 = valid_23_27 ? 5'h1b : _T_9326; // @[Mux.scala 31:69:@3835.4]
  assign _T_9328 = valid_23_26 ? 5'h1a : _T_9327; // @[Mux.scala 31:69:@3836.4]
  assign _T_9329 = valid_23_25 ? 5'h19 : _T_9328; // @[Mux.scala 31:69:@3837.4]
  assign _T_9330 = valid_23_24 ? 5'h18 : _T_9329; // @[Mux.scala 31:69:@3838.4]
  assign _T_9331 = valid_23_23 ? 5'h17 : _T_9330; // @[Mux.scala 31:69:@3839.4]
  assign _T_9332 = valid_23_22 ? 5'h16 : _T_9331; // @[Mux.scala 31:69:@3840.4]
  assign _T_9333 = valid_23_21 ? 5'h15 : _T_9332; // @[Mux.scala 31:69:@3841.4]
  assign _T_9334 = valid_23_20 ? 5'h14 : _T_9333; // @[Mux.scala 31:69:@3842.4]
  assign _T_9335 = valid_23_19 ? 5'h13 : _T_9334; // @[Mux.scala 31:69:@3843.4]
  assign _T_9336 = valid_23_18 ? 5'h12 : _T_9335; // @[Mux.scala 31:69:@3844.4]
  assign _T_9337 = valid_23_17 ? 5'h11 : _T_9336; // @[Mux.scala 31:69:@3845.4]
  assign _T_9338 = valid_23_16 ? 5'h10 : _T_9337; // @[Mux.scala 31:69:@3846.4]
  assign _T_9339 = valid_23_15 ? 5'hf : _T_9338; // @[Mux.scala 31:69:@3847.4]
  assign _T_9340 = valid_23_14 ? 5'he : _T_9339; // @[Mux.scala 31:69:@3848.4]
  assign _T_9341 = valid_23_13 ? 5'hd : _T_9340; // @[Mux.scala 31:69:@3849.4]
  assign _T_9342 = valid_23_12 ? 5'hc : _T_9341; // @[Mux.scala 31:69:@3850.4]
  assign _T_9343 = valid_23_11 ? 5'hb : _T_9342; // @[Mux.scala 31:69:@3851.4]
  assign _T_9344 = valid_23_10 ? 5'ha : _T_9343; // @[Mux.scala 31:69:@3852.4]
  assign _T_9345 = valid_23_9 ? 5'h9 : _T_9344; // @[Mux.scala 31:69:@3853.4]
  assign _T_9346 = valid_23_8 ? 5'h8 : _T_9345; // @[Mux.scala 31:69:@3854.4]
  assign _T_9347 = valid_23_7 ? 5'h7 : _T_9346; // @[Mux.scala 31:69:@3855.4]
  assign _T_9348 = valid_23_6 ? 5'h6 : _T_9347; // @[Mux.scala 31:69:@3856.4]
  assign _T_9349 = valid_23_5 ? 5'h5 : _T_9348; // @[Mux.scala 31:69:@3857.4]
  assign _T_9350 = valid_23_4 ? 5'h4 : _T_9349; // @[Mux.scala 31:69:@3858.4]
  assign _T_9351 = valid_23_3 ? 5'h3 : _T_9350; // @[Mux.scala 31:69:@3859.4]
  assign _T_9352 = valid_23_2 ? 5'h2 : _T_9351; // @[Mux.scala 31:69:@3860.4]
  assign _T_9353 = valid_23_1 ? 5'h1 : _T_9352; // @[Mux.scala 31:69:@3861.4]
  assign select_23 = valid_23_0 ? 5'h0 : _T_9353; // @[Mux.scala 31:69:@3862.4]
  assign _GEN_737 = 5'h1 == select_23 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@3864.4]
  assign _GEN_738 = 5'h2 == select_23 ? io_inData_2 : _GEN_737; // @[Switch.scala 33:19:@3864.4]
  assign _GEN_739 = 5'h3 == select_23 ? io_inData_3 : _GEN_738; // @[Switch.scala 33:19:@3864.4]
  assign _GEN_740 = 5'h4 == select_23 ? io_inData_4 : _GEN_739; // @[Switch.scala 33:19:@3864.4]
  assign _GEN_741 = 5'h5 == select_23 ? io_inData_5 : _GEN_740; // @[Switch.scala 33:19:@3864.4]
  assign _GEN_742 = 5'h6 == select_23 ? io_inData_6 : _GEN_741; // @[Switch.scala 33:19:@3864.4]
  assign _GEN_743 = 5'h7 == select_23 ? io_inData_7 : _GEN_742; // @[Switch.scala 33:19:@3864.4]
  assign _GEN_744 = 5'h8 == select_23 ? io_inData_8 : _GEN_743; // @[Switch.scala 33:19:@3864.4]
  assign _GEN_745 = 5'h9 == select_23 ? io_inData_9 : _GEN_744; // @[Switch.scala 33:19:@3864.4]
  assign _GEN_746 = 5'ha == select_23 ? io_inData_10 : _GEN_745; // @[Switch.scala 33:19:@3864.4]
  assign _GEN_747 = 5'hb == select_23 ? io_inData_11 : _GEN_746; // @[Switch.scala 33:19:@3864.4]
  assign _GEN_748 = 5'hc == select_23 ? io_inData_12 : _GEN_747; // @[Switch.scala 33:19:@3864.4]
  assign _GEN_749 = 5'hd == select_23 ? io_inData_13 : _GEN_748; // @[Switch.scala 33:19:@3864.4]
  assign _GEN_750 = 5'he == select_23 ? io_inData_14 : _GEN_749; // @[Switch.scala 33:19:@3864.4]
  assign _GEN_751 = 5'hf == select_23 ? io_inData_15 : _GEN_750; // @[Switch.scala 33:19:@3864.4]
  assign _GEN_752 = 5'h10 == select_23 ? io_inData_16 : _GEN_751; // @[Switch.scala 33:19:@3864.4]
  assign _GEN_753 = 5'h11 == select_23 ? io_inData_17 : _GEN_752; // @[Switch.scala 33:19:@3864.4]
  assign _GEN_754 = 5'h12 == select_23 ? io_inData_18 : _GEN_753; // @[Switch.scala 33:19:@3864.4]
  assign _GEN_755 = 5'h13 == select_23 ? io_inData_19 : _GEN_754; // @[Switch.scala 33:19:@3864.4]
  assign _GEN_756 = 5'h14 == select_23 ? io_inData_20 : _GEN_755; // @[Switch.scala 33:19:@3864.4]
  assign _GEN_757 = 5'h15 == select_23 ? io_inData_21 : _GEN_756; // @[Switch.scala 33:19:@3864.4]
  assign _GEN_758 = 5'h16 == select_23 ? io_inData_22 : _GEN_757; // @[Switch.scala 33:19:@3864.4]
  assign _GEN_759 = 5'h17 == select_23 ? io_inData_23 : _GEN_758; // @[Switch.scala 33:19:@3864.4]
  assign _GEN_760 = 5'h18 == select_23 ? io_inData_24 : _GEN_759; // @[Switch.scala 33:19:@3864.4]
  assign _GEN_761 = 5'h19 == select_23 ? io_inData_25 : _GEN_760; // @[Switch.scala 33:19:@3864.4]
  assign _GEN_762 = 5'h1a == select_23 ? io_inData_26 : _GEN_761; // @[Switch.scala 33:19:@3864.4]
  assign _GEN_763 = 5'h1b == select_23 ? io_inData_27 : _GEN_762; // @[Switch.scala 33:19:@3864.4]
  assign _GEN_764 = 5'h1c == select_23 ? io_inData_28 : _GEN_763; // @[Switch.scala 33:19:@3864.4]
  assign _GEN_765 = 5'h1d == select_23 ? io_inData_29 : _GEN_764; // @[Switch.scala 33:19:@3864.4]
  assign _GEN_766 = 5'h1e == select_23 ? io_inData_30 : _GEN_765; // @[Switch.scala 33:19:@3864.4]
  assign _T_9362 = {valid_23_7,valid_23_6,valid_23_5,valid_23_4,valid_23_3,valid_23_2,valid_23_1,valid_23_0}; // @[Switch.scala 34:32:@3871.4]
  assign _T_9370 = {valid_23_15,valid_23_14,valid_23_13,valid_23_12,valid_23_11,valid_23_10,valid_23_9,valid_23_8,_T_9362}; // @[Switch.scala 34:32:@3879.4]
  assign _T_9377 = {valid_23_23,valid_23_22,valid_23_21,valid_23_20,valid_23_19,valid_23_18,valid_23_17,valid_23_16}; // @[Switch.scala 34:32:@3886.4]
  assign _T_9386 = {valid_23_31,valid_23_30,valid_23_29,valid_23_28,valid_23_27,valid_23_26,valid_23_25,valid_23_24,_T_9377,_T_9370}; // @[Switch.scala 34:32:@3895.4]
  assign _T_9390 = io_inAddr_0 == 5'h18; // @[Switch.scala 30:53:@3898.4]
  assign valid_24_0 = io_inValid_0 & _T_9390; // @[Switch.scala 30:36:@3899.4]
  assign _T_9393 = io_inAddr_1 == 5'h18; // @[Switch.scala 30:53:@3901.4]
  assign valid_24_1 = io_inValid_1 & _T_9393; // @[Switch.scala 30:36:@3902.4]
  assign _T_9396 = io_inAddr_2 == 5'h18; // @[Switch.scala 30:53:@3904.4]
  assign valid_24_2 = io_inValid_2 & _T_9396; // @[Switch.scala 30:36:@3905.4]
  assign _T_9399 = io_inAddr_3 == 5'h18; // @[Switch.scala 30:53:@3907.4]
  assign valid_24_3 = io_inValid_3 & _T_9399; // @[Switch.scala 30:36:@3908.4]
  assign _T_9402 = io_inAddr_4 == 5'h18; // @[Switch.scala 30:53:@3910.4]
  assign valid_24_4 = io_inValid_4 & _T_9402; // @[Switch.scala 30:36:@3911.4]
  assign _T_9405 = io_inAddr_5 == 5'h18; // @[Switch.scala 30:53:@3913.4]
  assign valid_24_5 = io_inValid_5 & _T_9405; // @[Switch.scala 30:36:@3914.4]
  assign _T_9408 = io_inAddr_6 == 5'h18; // @[Switch.scala 30:53:@3916.4]
  assign valid_24_6 = io_inValid_6 & _T_9408; // @[Switch.scala 30:36:@3917.4]
  assign _T_9411 = io_inAddr_7 == 5'h18; // @[Switch.scala 30:53:@3919.4]
  assign valid_24_7 = io_inValid_7 & _T_9411; // @[Switch.scala 30:36:@3920.4]
  assign _T_9414 = io_inAddr_8 == 5'h18; // @[Switch.scala 30:53:@3922.4]
  assign valid_24_8 = io_inValid_8 & _T_9414; // @[Switch.scala 30:36:@3923.4]
  assign _T_9417 = io_inAddr_9 == 5'h18; // @[Switch.scala 30:53:@3925.4]
  assign valid_24_9 = io_inValid_9 & _T_9417; // @[Switch.scala 30:36:@3926.4]
  assign _T_9420 = io_inAddr_10 == 5'h18; // @[Switch.scala 30:53:@3928.4]
  assign valid_24_10 = io_inValid_10 & _T_9420; // @[Switch.scala 30:36:@3929.4]
  assign _T_9423 = io_inAddr_11 == 5'h18; // @[Switch.scala 30:53:@3931.4]
  assign valid_24_11 = io_inValid_11 & _T_9423; // @[Switch.scala 30:36:@3932.4]
  assign _T_9426 = io_inAddr_12 == 5'h18; // @[Switch.scala 30:53:@3934.4]
  assign valid_24_12 = io_inValid_12 & _T_9426; // @[Switch.scala 30:36:@3935.4]
  assign _T_9429 = io_inAddr_13 == 5'h18; // @[Switch.scala 30:53:@3937.4]
  assign valid_24_13 = io_inValid_13 & _T_9429; // @[Switch.scala 30:36:@3938.4]
  assign _T_9432 = io_inAddr_14 == 5'h18; // @[Switch.scala 30:53:@3940.4]
  assign valid_24_14 = io_inValid_14 & _T_9432; // @[Switch.scala 30:36:@3941.4]
  assign _T_9435 = io_inAddr_15 == 5'h18; // @[Switch.scala 30:53:@3943.4]
  assign valid_24_15 = io_inValid_15 & _T_9435; // @[Switch.scala 30:36:@3944.4]
  assign _T_9438 = io_inAddr_16 == 5'h18; // @[Switch.scala 30:53:@3946.4]
  assign valid_24_16 = io_inValid_16 & _T_9438; // @[Switch.scala 30:36:@3947.4]
  assign _T_9441 = io_inAddr_17 == 5'h18; // @[Switch.scala 30:53:@3949.4]
  assign valid_24_17 = io_inValid_17 & _T_9441; // @[Switch.scala 30:36:@3950.4]
  assign _T_9444 = io_inAddr_18 == 5'h18; // @[Switch.scala 30:53:@3952.4]
  assign valid_24_18 = io_inValid_18 & _T_9444; // @[Switch.scala 30:36:@3953.4]
  assign _T_9447 = io_inAddr_19 == 5'h18; // @[Switch.scala 30:53:@3955.4]
  assign valid_24_19 = io_inValid_19 & _T_9447; // @[Switch.scala 30:36:@3956.4]
  assign _T_9450 = io_inAddr_20 == 5'h18; // @[Switch.scala 30:53:@3958.4]
  assign valid_24_20 = io_inValid_20 & _T_9450; // @[Switch.scala 30:36:@3959.4]
  assign _T_9453 = io_inAddr_21 == 5'h18; // @[Switch.scala 30:53:@3961.4]
  assign valid_24_21 = io_inValid_21 & _T_9453; // @[Switch.scala 30:36:@3962.4]
  assign _T_9456 = io_inAddr_22 == 5'h18; // @[Switch.scala 30:53:@3964.4]
  assign valid_24_22 = io_inValid_22 & _T_9456; // @[Switch.scala 30:36:@3965.4]
  assign _T_9459 = io_inAddr_23 == 5'h18; // @[Switch.scala 30:53:@3967.4]
  assign valid_24_23 = io_inValid_23 & _T_9459; // @[Switch.scala 30:36:@3968.4]
  assign _T_9462 = io_inAddr_24 == 5'h18; // @[Switch.scala 30:53:@3970.4]
  assign valid_24_24 = io_inValid_24 & _T_9462; // @[Switch.scala 30:36:@3971.4]
  assign _T_9465 = io_inAddr_25 == 5'h18; // @[Switch.scala 30:53:@3973.4]
  assign valid_24_25 = io_inValid_25 & _T_9465; // @[Switch.scala 30:36:@3974.4]
  assign _T_9468 = io_inAddr_26 == 5'h18; // @[Switch.scala 30:53:@3976.4]
  assign valid_24_26 = io_inValid_26 & _T_9468; // @[Switch.scala 30:36:@3977.4]
  assign _T_9471 = io_inAddr_27 == 5'h18; // @[Switch.scala 30:53:@3979.4]
  assign valid_24_27 = io_inValid_27 & _T_9471; // @[Switch.scala 30:36:@3980.4]
  assign _T_9474 = io_inAddr_28 == 5'h18; // @[Switch.scala 30:53:@3982.4]
  assign valid_24_28 = io_inValid_28 & _T_9474; // @[Switch.scala 30:36:@3983.4]
  assign _T_9477 = io_inAddr_29 == 5'h18; // @[Switch.scala 30:53:@3985.4]
  assign valid_24_29 = io_inValid_29 & _T_9477; // @[Switch.scala 30:36:@3986.4]
  assign _T_9480 = io_inAddr_30 == 5'h18; // @[Switch.scala 30:53:@3988.4]
  assign valid_24_30 = io_inValid_30 & _T_9480; // @[Switch.scala 30:36:@3989.4]
  assign _T_9483 = io_inAddr_31 == 5'h18; // @[Switch.scala 30:53:@3991.4]
  assign valid_24_31 = io_inValid_31 & _T_9483; // @[Switch.scala 30:36:@3992.4]
  assign _T_9517 = valid_24_30 ? 5'h1e : 5'h1f; // @[Mux.scala 31:69:@3994.4]
  assign _T_9518 = valid_24_29 ? 5'h1d : _T_9517; // @[Mux.scala 31:69:@3995.4]
  assign _T_9519 = valid_24_28 ? 5'h1c : _T_9518; // @[Mux.scala 31:69:@3996.4]
  assign _T_9520 = valid_24_27 ? 5'h1b : _T_9519; // @[Mux.scala 31:69:@3997.4]
  assign _T_9521 = valid_24_26 ? 5'h1a : _T_9520; // @[Mux.scala 31:69:@3998.4]
  assign _T_9522 = valid_24_25 ? 5'h19 : _T_9521; // @[Mux.scala 31:69:@3999.4]
  assign _T_9523 = valid_24_24 ? 5'h18 : _T_9522; // @[Mux.scala 31:69:@4000.4]
  assign _T_9524 = valid_24_23 ? 5'h17 : _T_9523; // @[Mux.scala 31:69:@4001.4]
  assign _T_9525 = valid_24_22 ? 5'h16 : _T_9524; // @[Mux.scala 31:69:@4002.4]
  assign _T_9526 = valid_24_21 ? 5'h15 : _T_9525; // @[Mux.scala 31:69:@4003.4]
  assign _T_9527 = valid_24_20 ? 5'h14 : _T_9526; // @[Mux.scala 31:69:@4004.4]
  assign _T_9528 = valid_24_19 ? 5'h13 : _T_9527; // @[Mux.scala 31:69:@4005.4]
  assign _T_9529 = valid_24_18 ? 5'h12 : _T_9528; // @[Mux.scala 31:69:@4006.4]
  assign _T_9530 = valid_24_17 ? 5'h11 : _T_9529; // @[Mux.scala 31:69:@4007.4]
  assign _T_9531 = valid_24_16 ? 5'h10 : _T_9530; // @[Mux.scala 31:69:@4008.4]
  assign _T_9532 = valid_24_15 ? 5'hf : _T_9531; // @[Mux.scala 31:69:@4009.4]
  assign _T_9533 = valid_24_14 ? 5'he : _T_9532; // @[Mux.scala 31:69:@4010.4]
  assign _T_9534 = valid_24_13 ? 5'hd : _T_9533; // @[Mux.scala 31:69:@4011.4]
  assign _T_9535 = valid_24_12 ? 5'hc : _T_9534; // @[Mux.scala 31:69:@4012.4]
  assign _T_9536 = valid_24_11 ? 5'hb : _T_9535; // @[Mux.scala 31:69:@4013.4]
  assign _T_9537 = valid_24_10 ? 5'ha : _T_9536; // @[Mux.scala 31:69:@4014.4]
  assign _T_9538 = valid_24_9 ? 5'h9 : _T_9537; // @[Mux.scala 31:69:@4015.4]
  assign _T_9539 = valid_24_8 ? 5'h8 : _T_9538; // @[Mux.scala 31:69:@4016.4]
  assign _T_9540 = valid_24_7 ? 5'h7 : _T_9539; // @[Mux.scala 31:69:@4017.4]
  assign _T_9541 = valid_24_6 ? 5'h6 : _T_9540; // @[Mux.scala 31:69:@4018.4]
  assign _T_9542 = valid_24_5 ? 5'h5 : _T_9541; // @[Mux.scala 31:69:@4019.4]
  assign _T_9543 = valid_24_4 ? 5'h4 : _T_9542; // @[Mux.scala 31:69:@4020.4]
  assign _T_9544 = valid_24_3 ? 5'h3 : _T_9543; // @[Mux.scala 31:69:@4021.4]
  assign _T_9545 = valid_24_2 ? 5'h2 : _T_9544; // @[Mux.scala 31:69:@4022.4]
  assign _T_9546 = valid_24_1 ? 5'h1 : _T_9545; // @[Mux.scala 31:69:@4023.4]
  assign select_24 = valid_24_0 ? 5'h0 : _T_9546; // @[Mux.scala 31:69:@4024.4]
  assign _GEN_769 = 5'h1 == select_24 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@4026.4]
  assign _GEN_770 = 5'h2 == select_24 ? io_inData_2 : _GEN_769; // @[Switch.scala 33:19:@4026.4]
  assign _GEN_771 = 5'h3 == select_24 ? io_inData_3 : _GEN_770; // @[Switch.scala 33:19:@4026.4]
  assign _GEN_772 = 5'h4 == select_24 ? io_inData_4 : _GEN_771; // @[Switch.scala 33:19:@4026.4]
  assign _GEN_773 = 5'h5 == select_24 ? io_inData_5 : _GEN_772; // @[Switch.scala 33:19:@4026.4]
  assign _GEN_774 = 5'h6 == select_24 ? io_inData_6 : _GEN_773; // @[Switch.scala 33:19:@4026.4]
  assign _GEN_775 = 5'h7 == select_24 ? io_inData_7 : _GEN_774; // @[Switch.scala 33:19:@4026.4]
  assign _GEN_776 = 5'h8 == select_24 ? io_inData_8 : _GEN_775; // @[Switch.scala 33:19:@4026.4]
  assign _GEN_777 = 5'h9 == select_24 ? io_inData_9 : _GEN_776; // @[Switch.scala 33:19:@4026.4]
  assign _GEN_778 = 5'ha == select_24 ? io_inData_10 : _GEN_777; // @[Switch.scala 33:19:@4026.4]
  assign _GEN_779 = 5'hb == select_24 ? io_inData_11 : _GEN_778; // @[Switch.scala 33:19:@4026.4]
  assign _GEN_780 = 5'hc == select_24 ? io_inData_12 : _GEN_779; // @[Switch.scala 33:19:@4026.4]
  assign _GEN_781 = 5'hd == select_24 ? io_inData_13 : _GEN_780; // @[Switch.scala 33:19:@4026.4]
  assign _GEN_782 = 5'he == select_24 ? io_inData_14 : _GEN_781; // @[Switch.scala 33:19:@4026.4]
  assign _GEN_783 = 5'hf == select_24 ? io_inData_15 : _GEN_782; // @[Switch.scala 33:19:@4026.4]
  assign _GEN_784 = 5'h10 == select_24 ? io_inData_16 : _GEN_783; // @[Switch.scala 33:19:@4026.4]
  assign _GEN_785 = 5'h11 == select_24 ? io_inData_17 : _GEN_784; // @[Switch.scala 33:19:@4026.4]
  assign _GEN_786 = 5'h12 == select_24 ? io_inData_18 : _GEN_785; // @[Switch.scala 33:19:@4026.4]
  assign _GEN_787 = 5'h13 == select_24 ? io_inData_19 : _GEN_786; // @[Switch.scala 33:19:@4026.4]
  assign _GEN_788 = 5'h14 == select_24 ? io_inData_20 : _GEN_787; // @[Switch.scala 33:19:@4026.4]
  assign _GEN_789 = 5'h15 == select_24 ? io_inData_21 : _GEN_788; // @[Switch.scala 33:19:@4026.4]
  assign _GEN_790 = 5'h16 == select_24 ? io_inData_22 : _GEN_789; // @[Switch.scala 33:19:@4026.4]
  assign _GEN_791 = 5'h17 == select_24 ? io_inData_23 : _GEN_790; // @[Switch.scala 33:19:@4026.4]
  assign _GEN_792 = 5'h18 == select_24 ? io_inData_24 : _GEN_791; // @[Switch.scala 33:19:@4026.4]
  assign _GEN_793 = 5'h19 == select_24 ? io_inData_25 : _GEN_792; // @[Switch.scala 33:19:@4026.4]
  assign _GEN_794 = 5'h1a == select_24 ? io_inData_26 : _GEN_793; // @[Switch.scala 33:19:@4026.4]
  assign _GEN_795 = 5'h1b == select_24 ? io_inData_27 : _GEN_794; // @[Switch.scala 33:19:@4026.4]
  assign _GEN_796 = 5'h1c == select_24 ? io_inData_28 : _GEN_795; // @[Switch.scala 33:19:@4026.4]
  assign _GEN_797 = 5'h1d == select_24 ? io_inData_29 : _GEN_796; // @[Switch.scala 33:19:@4026.4]
  assign _GEN_798 = 5'h1e == select_24 ? io_inData_30 : _GEN_797; // @[Switch.scala 33:19:@4026.4]
  assign _T_9555 = {valid_24_7,valid_24_6,valid_24_5,valid_24_4,valid_24_3,valid_24_2,valid_24_1,valid_24_0}; // @[Switch.scala 34:32:@4033.4]
  assign _T_9563 = {valid_24_15,valid_24_14,valid_24_13,valid_24_12,valid_24_11,valid_24_10,valid_24_9,valid_24_8,_T_9555}; // @[Switch.scala 34:32:@4041.4]
  assign _T_9570 = {valid_24_23,valid_24_22,valid_24_21,valid_24_20,valid_24_19,valid_24_18,valid_24_17,valid_24_16}; // @[Switch.scala 34:32:@4048.4]
  assign _T_9579 = {valid_24_31,valid_24_30,valid_24_29,valid_24_28,valid_24_27,valid_24_26,valid_24_25,valid_24_24,_T_9570,_T_9563}; // @[Switch.scala 34:32:@4057.4]
  assign _T_9583 = io_inAddr_0 == 5'h19; // @[Switch.scala 30:53:@4060.4]
  assign valid_25_0 = io_inValid_0 & _T_9583; // @[Switch.scala 30:36:@4061.4]
  assign _T_9586 = io_inAddr_1 == 5'h19; // @[Switch.scala 30:53:@4063.4]
  assign valid_25_1 = io_inValid_1 & _T_9586; // @[Switch.scala 30:36:@4064.4]
  assign _T_9589 = io_inAddr_2 == 5'h19; // @[Switch.scala 30:53:@4066.4]
  assign valid_25_2 = io_inValid_2 & _T_9589; // @[Switch.scala 30:36:@4067.4]
  assign _T_9592 = io_inAddr_3 == 5'h19; // @[Switch.scala 30:53:@4069.4]
  assign valid_25_3 = io_inValid_3 & _T_9592; // @[Switch.scala 30:36:@4070.4]
  assign _T_9595 = io_inAddr_4 == 5'h19; // @[Switch.scala 30:53:@4072.4]
  assign valid_25_4 = io_inValid_4 & _T_9595; // @[Switch.scala 30:36:@4073.4]
  assign _T_9598 = io_inAddr_5 == 5'h19; // @[Switch.scala 30:53:@4075.4]
  assign valid_25_5 = io_inValid_5 & _T_9598; // @[Switch.scala 30:36:@4076.4]
  assign _T_9601 = io_inAddr_6 == 5'h19; // @[Switch.scala 30:53:@4078.4]
  assign valid_25_6 = io_inValid_6 & _T_9601; // @[Switch.scala 30:36:@4079.4]
  assign _T_9604 = io_inAddr_7 == 5'h19; // @[Switch.scala 30:53:@4081.4]
  assign valid_25_7 = io_inValid_7 & _T_9604; // @[Switch.scala 30:36:@4082.4]
  assign _T_9607 = io_inAddr_8 == 5'h19; // @[Switch.scala 30:53:@4084.4]
  assign valid_25_8 = io_inValid_8 & _T_9607; // @[Switch.scala 30:36:@4085.4]
  assign _T_9610 = io_inAddr_9 == 5'h19; // @[Switch.scala 30:53:@4087.4]
  assign valid_25_9 = io_inValid_9 & _T_9610; // @[Switch.scala 30:36:@4088.4]
  assign _T_9613 = io_inAddr_10 == 5'h19; // @[Switch.scala 30:53:@4090.4]
  assign valid_25_10 = io_inValid_10 & _T_9613; // @[Switch.scala 30:36:@4091.4]
  assign _T_9616 = io_inAddr_11 == 5'h19; // @[Switch.scala 30:53:@4093.4]
  assign valid_25_11 = io_inValid_11 & _T_9616; // @[Switch.scala 30:36:@4094.4]
  assign _T_9619 = io_inAddr_12 == 5'h19; // @[Switch.scala 30:53:@4096.4]
  assign valid_25_12 = io_inValid_12 & _T_9619; // @[Switch.scala 30:36:@4097.4]
  assign _T_9622 = io_inAddr_13 == 5'h19; // @[Switch.scala 30:53:@4099.4]
  assign valid_25_13 = io_inValid_13 & _T_9622; // @[Switch.scala 30:36:@4100.4]
  assign _T_9625 = io_inAddr_14 == 5'h19; // @[Switch.scala 30:53:@4102.4]
  assign valid_25_14 = io_inValid_14 & _T_9625; // @[Switch.scala 30:36:@4103.4]
  assign _T_9628 = io_inAddr_15 == 5'h19; // @[Switch.scala 30:53:@4105.4]
  assign valid_25_15 = io_inValid_15 & _T_9628; // @[Switch.scala 30:36:@4106.4]
  assign _T_9631 = io_inAddr_16 == 5'h19; // @[Switch.scala 30:53:@4108.4]
  assign valid_25_16 = io_inValid_16 & _T_9631; // @[Switch.scala 30:36:@4109.4]
  assign _T_9634 = io_inAddr_17 == 5'h19; // @[Switch.scala 30:53:@4111.4]
  assign valid_25_17 = io_inValid_17 & _T_9634; // @[Switch.scala 30:36:@4112.4]
  assign _T_9637 = io_inAddr_18 == 5'h19; // @[Switch.scala 30:53:@4114.4]
  assign valid_25_18 = io_inValid_18 & _T_9637; // @[Switch.scala 30:36:@4115.4]
  assign _T_9640 = io_inAddr_19 == 5'h19; // @[Switch.scala 30:53:@4117.4]
  assign valid_25_19 = io_inValid_19 & _T_9640; // @[Switch.scala 30:36:@4118.4]
  assign _T_9643 = io_inAddr_20 == 5'h19; // @[Switch.scala 30:53:@4120.4]
  assign valid_25_20 = io_inValid_20 & _T_9643; // @[Switch.scala 30:36:@4121.4]
  assign _T_9646 = io_inAddr_21 == 5'h19; // @[Switch.scala 30:53:@4123.4]
  assign valid_25_21 = io_inValid_21 & _T_9646; // @[Switch.scala 30:36:@4124.4]
  assign _T_9649 = io_inAddr_22 == 5'h19; // @[Switch.scala 30:53:@4126.4]
  assign valid_25_22 = io_inValid_22 & _T_9649; // @[Switch.scala 30:36:@4127.4]
  assign _T_9652 = io_inAddr_23 == 5'h19; // @[Switch.scala 30:53:@4129.4]
  assign valid_25_23 = io_inValid_23 & _T_9652; // @[Switch.scala 30:36:@4130.4]
  assign _T_9655 = io_inAddr_24 == 5'h19; // @[Switch.scala 30:53:@4132.4]
  assign valid_25_24 = io_inValid_24 & _T_9655; // @[Switch.scala 30:36:@4133.4]
  assign _T_9658 = io_inAddr_25 == 5'h19; // @[Switch.scala 30:53:@4135.4]
  assign valid_25_25 = io_inValid_25 & _T_9658; // @[Switch.scala 30:36:@4136.4]
  assign _T_9661 = io_inAddr_26 == 5'h19; // @[Switch.scala 30:53:@4138.4]
  assign valid_25_26 = io_inValid_26 & _T_9661; // @[Switch.scala 30:36:@4139.4]
  assign _T_9664 = io_inAddr_27 == 5'h19; // @[Switch.scala 30:53:@4141.4]
  assign valid_25_27 = io_inValid_27 & _T_9664; // @[Switch.scala 30:36:@4142.4]
  assign _T_9667 = io_inAddr_28 == 5'h19; // @[Switch.scala 30:53:@4144.4]
  assign valid_25_28 = io_inValid_28 & _T_9667; // @[Switch.scala 30:36:@4145.4]
  assign _T_9670 = io_inAddr_29 == 5'h19; // @[Switch.scala 30:53:@4147.4]
  assign valid_25_29 = io_inValid_29 & _T_9670; // @[Switch.scala 30:36:@4148.4]
  assign _T_9673 = io_inAddr_30 == 5'h19; // @[Switch.scala 30:53:@4150.4]
  assign valid_25_30 = io_inValid_30 & _T_9673; // @[Switch.scala 30:36:@4151.4]
  assign _T_9676 = io_inAddr_31 == 5'h19; // @[Switch.scala 30:53:@4153.4]
  assign valid_25_31 = io_inValid_31 & _T_9676; // @[Switch.scala 30:36:@4154.4]
  assign _T_9710 = valid_25_30 ? 5'h1e : 5'h1f; // @[Mux.scala 31:69:@4156.4]
  assign _T_9711 = valid_25_29 ? 5'h1d : _T_9710; // @[Mux.scala 31:69:@4157.4]
  assign _T_9712 = valid_25_28 ? 5'h1c : _T_9711; // @[Mux.scala 31:69:@4158.4]
  assign _T_9713 = valid_25_27 ? 5'h1b : _T_9712; // @[Mux.scala 31:69:@4159.4]
  assign _T_9714 = valid_25_26 ? 5'h1a : _T_9713; // @[Mux.scala 31:69:@4160.4]
  assign _T_9715 = valid_25_25 ? 5'h19 : _T_9714; // @[Mux.scala 31:69:@4161.4]
  assign _T_9716 = valid_25_24 ? 5'h18 : _T_9715; // @[Mux.scala 31:69:@4162.4]
  assign _T_9717 = valid_25_23 ? 5'h17 : _T_9716; // @[Mux.scala 31:69:@4163.4]
  assign _T_9718 = valid_25_22 ? 5'h16 : _T_9717; // @[Mux.scala 31:69:@4164.4]
  assign _T_9719 = valid_25_21 ? 5'h15 : _T_9718; // @[Mux.scala 31:69:@4165.4]
  assign _T_9720 = valid_25_20 ? 5'h14 : _T_9719; // @[Mux.scala 31:69:@4166.4]
  assign _T_9721 = valid_25_19 ? 5'h13 : _T_9720; // @[Mux.scala 31:69:@4167.4]
  assign _T_9722 = valid_25_18 ? 5'h12 : _T_9721; // @[Mux.scala 31:69:@4168.4]
  assign _T_9723 = valid_25_17 ? 5'h11 : _T_9722; // @[Mux.scala 31:69:@4169.4]
  assign _T_9724 = valid_25_16 ? 5'h10 : _T_9723; // @[Mux.scala 31:69:@4170.4]
  assign _T_9725 = valid_25_15 ? 5'hf : _T_9724; // @[Mux.scala 31:69:@4171.4]
  assign _T_9726 = valid_25_14 ? 5'he : _T_9725; // @[Mux.scala 31:69:@4172.4]
  assign _T_9727 = valid_25_13 ? 5'hd : _T_9726; // @[Mux.scala 31:69:@4173.4]
  assign _T_9728 = valid_25_12 ? 5'hc : _T_9727; // @[Mux.scala 31:69:@4174.4]
  assign _T_9729 = valid_25_11 ? 5'hb : _T_9728; // @[Mux.scala 31:69:@4175.4]
  assign _T_9730 = valid_25_10 ? 5'ha : _T_9729; // @[Mux.scala 31:69:@4176.4]
  assign _T_9731 = valid_25_9 ? 5'h9 : _T_9730; // @[Mux.scala 31:69:@4177.4]
  assign _T_9732 = valid_25_8 ? 5'h8 : _T_9731; // @[Mux.scala 31:69:@4178.4]
  assign _T_9733 = valid_25_7 ? 5'h7 : _T_9732; // @[Mux.scala 31:69:@4179.4]
  assign _T_9734 = valid_25_6 ? 5'h6 : _T_9733; // @[Mux.scala 31:69:@4180.4]
  assign _T_9735 = valid_25_5 ? 5'h5 : _T_9734; // @[Mux.scala 31:69:@4181.4]
  assign _T_9736 = valid_25_4 ? 5'h4 : _T_9735; // @[Mux.scala 31:69:@4182.4]
  assign _T_9737 = valid_25_3 ? 5'h3 : _T_9736; // @[Mux.scala 31:69:@4183.4]
  assign _T_9738 = valid_25_2 ? 5'h2 : _T_9737; // @[Mux.scala 31:69:@4184.4]
  assign _T_9739 = valid_25_1 ? 5'h1 : _T_9738; // @[Mux.scala 31:69:@4185.4]
  assign select_25 = valid_25_0 ? 5'h0 : _T_9739; // @[Mux.scala 31:69:@4186.4]
  assign _GEN_801 = 5'h1 == select_25 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@4188.4]
  assign _GEN_802 = 5'h2 == select_25 ? io_inData_2 : _GEN_801; // @[Switch.scala 33:19:@4188.4]
  assign _GEN_803 = 5'h3 == select_25 ? io_inData_3 : _GEN_802; // @[Switch.scala 33:19:@4188.4]
  assign _GEN_804 = 5'h4 == select_25 ? io_inData_4 : _GEN_803; // @[Switch.scala 33:19:@4188.4]
  assign _GEN_805 = 5'h5 == select_25 ? io_inData_5 : _GEN_804; // @[Switch.scala 33:19:@4188.4]
  assign _GEN_806 = 5'h6 == select_25 ? io_inData_6 : _GEN_805; // @[Switch.scala 33:19:@4188.4]
  assign _GEN_807 = 5'h7 == select_25 ? io_inData_7 : _GEN_806; // @[Switch.scala 33:19:@4188.4]
  assign _GEN_808 = 5'h8 == select_25 ? io_inData_8 : _GEN_807; // @[Switch.scala 33:19:@4188.4]
  assign _GEN_809 = 5'h9 == select_25 ? io_inData_9 : _GEN_808; // @[Switch.scala 33:19:@4188.4]
  assign _GEN_810 = 5'ha == select_25 ? io_inData_10 : _GEN_809; // @[Switch.scala 33:19:@4188.4]
  assign _GEN_811 = 5'hb == select_25 ? io_inData_11 : _GEN_810; // @[Switch.scala 33:19:@4188.4]
  assign _GEN_812 = 5'hc == select_25 ? io_inData_12 : _GEN_811; // @[Switch.scala 33:19:@4188.4]
  assign _GEN_813 = 5'hd == select_25 ? io_inData_13 : _GEN_812; // @[Switch.scala 33:19:@4188.4]
  assign _GEN_814 = 5'he == select_25 ? io_inData_14 : _GEN_813; // @[Switch.scala 33:19:@4188.4]
  assign _GEN_815 = 5'hf == select_25 ? io_inData_15 : _GEN_814; // @[Switch.scala 33:19:@4188.4]
  assign _GEN_816 = 5'h10 == select_25 ? io_inData_16 : _GEN_815; // @[Switch.scala 33:19:@4188.4]
  assign _GEN_817 = 5'h11 == select_25 ? io_inData_17 : _GEN_816; // @[Switch.scala 33:19:@4188.4]
  assign _GEN_818 = 5'h12 == select_25 ? io_inData_18 : _GEN_817; // @[Switch.scala 33:19:@4188.4]
  assign _GEN_819 = 5'h13 == select_25 ? io_inData_19 : _GEN_818; // @[Switch.scala 33:19:@4188.4]
  assign _GEN_820 = 5'h14 == select_25 ? io_inData_20 : _GEN_819; // @[Switch.scala 33:19:@4188.4]
  assign _GEN_821 = 5'h15 == select_25 ? io_inData_21 : _GEN_820; // @[Switch.scala 33:19:@4188.4]
  assign _GEN_822 = 5'h16 == select_25 ? io_inData_22 : _GEN_821; // @[Switch.scala 33:19:@4188.4]
  assign _GEN_823 = 5'h17 == select_25 ? io_inData_23 : _GEN_822; // @[Switch.scala 33:19:@4188.4]
  assign _GEN_824 = 5'h18 == select_25 ? io_inData_24 : _GEN_823; // @[Switch.scala 33:19:@4188.4]
  assign _GEN_825 = 5'h19 == select_25 ? io_inData_25 : _GEN_824; // @[Switch.scala 33:19:@4188.4]
  assign _GEN_826 = 5'h1a == select_25 ? io_inData_26 : _GEN_825; // @[Switch.scala 33:19:@4188.4]
  assign _GEN_827 = 5'h1b == select_25 ? io_inData_27 : _GEN_826; // @[Switch.scala 33:19:@4188.4]
  assign _GEN_828 = 5'h1c == select_25 ? io_inData_28 : _GEN_827; // @[Switch.scala 33:19:@4188.4]
  assign _GEN_829 = 5'h1d == select_25 ? io_inData_29 : _GEN_828; // @[Switch.scala 33:19:@4188.4]
  assign _GEN_830 = 5'h1e == select_25 ? io_inData_30 : _GEN_829; // @[Switch.scala 33:19:@4188.4]
  assign _T_9748 = {valid_25_7,valid_25_6,valid_25_5,valid_25_4,valid_25_3,valid_25_2,valid_25_1,valid_25_0}; // @[Switch.scala 34:32:@4195.4]
  assign _T_9756 = {valid_25_15,valid_25_14,valid_25_13,valid_25_12,valid_25_11,valid_25_10,valid_25_9,valid_25_8,_T_9748}; // @[Switch.scala 34:32:@4203.4]
  assign _T_9763 = {valid_25_23,valid_25_22,valid_25_21,valid_25_20,valid_25_19,valid_25_18,valid_25_17,valid_25_16}; // @[Switch.scala 34:32:@4210.4]
  assign _T_9772 = {valid_25_31,valid_25_30,valid_25_29,valid_25_28,valid_25_27,valid_25_26,valid_25_25,valid_25_24,_T_9763,_T_9756}; // @[Switch.scala 34:32:@4219.4]
  assign _T_9776 = io_inAddr_0 == 5'h1a; // @[Switch.scala 30:53:@4222.4]
  assign valid_26_0 = io_inValid_0 & _T_9776; // @[Switch.scala 30:36:@4223.4]
  assign _T_9779 = io_inAddr_1 == 5'h1a; // @[Switch.scala 30:53:@4225.4]
  assign valid_26_1 = io_inValid_1 & _T_9779; // @[Switch.scala 30:36:@4226.4]
  assign _T_9782 = io_inAddr_2 == 5'h1a; // @[Switch.scala 30:53:@4228.4]
  assign valid_26_2 = io_inValid_2 & _T_9782; // @[Switch.scala 30:36:@4229.4]
  assign _T_9785 = io_inAddr_3 == 5'h1a; // @[Switch.scala 30:53:@4231.4]
  assign valid_26_3 = io_inValid_3 & _T_9785; // @[Switch.scala 30:36:@4232.4]
  assign _T_9788 = io_inAddr_4 == 5'h1a; // @[Switch.scala 30:53:@4234.4]
  assign valid_26_4 = io_inValid_4 & _T_9788; // @[Switch.scala 30:36:@4235.4]
  assign _T_9791 = io_inAddr_5 == 5'h1a; // @[Switch.scala 30:53:@4237.4]
  assign valid_26_5 = io_inValid_5 & _T_9791; // @[Switch.scala 30:36:@4238.4]
  assign _T_9794 = io_inAddr_6 == 5'h1a; // @[Switch.scala 30:53:@4240.4]
  assign valid_26_6 = io_inValid_6 & _T_9794; // @[Switch.scala 30:36:@4241.4]
  assign _T_9797 = io_inAddr_7 == 5'h1a; // @[Switch.scala 30:53:@4243.4]
  assign valid_26_7 = io_inValid_7 & _T_9797; // @[Switch.scala 30:36:@4244.4]
  assign _T_9800 = io_inAddr_8 == 5'h1a; // @[Switch.scala 30:53:@4246.4]
  assign valid_26_8 = io_inValid_8 & _T_9800; // @[Switch.scala 30:36:@4247.4]
  assign _T_9803 = io_inAddr_9 == 5'h1a; // @[Switch.scala 30:53:@4249.4]
  assign valid_26_9 = io_inValid_9 & _T_9803; // @[Switch.scala 30:36:@4250.4]
  assign _T_9806 = io_inAddr_10 == 5'h1a; // @[Switch.scala 30:53:@4252.4]
  assign valid_26_10 = io_inValid_10 & _T_9806; // @[Switch.scala 30:36:@4253.4]
  assign _T_9809 = io_inAddr_11 == 5'h1a; // @[Switch.scala 30:53:@4255.4]
  assign valid_26_11 = io_inValid_11 & _T_9809; // @[Switch.scala 30:36:@4256.4]
  assign _T_9812 = io_inAddr_12 == 5'h1a; // @[Switch.scala 30:53:@4258.4]
  assign valid_26_12 = io_inValid_12 & _T_9812; // @[Switch.scala 30:36:@4259.4]
  assign _T_9815 = io_inAddr_13 == 5'h1a; // @[Switch.scala 30:53:@4261.4]
  assign valid_26_13 = io_inValid_13 & _T_9815; // @[Switch.scala 30:36:@4262.4]
  assign _T_9818 = io_inAddr_14 == 5'h1a; // @[Switch.scala 30:53:@4264.4]
  assign valid_26_14 = io_inValid_14 & _T_9818; // @[Switch.scala 30:36:@4265.4]
  assign _T_9821 = io_inAddr_15 == 5'h1a; // @[Switch.scala 30:53:@4267.4]
  assign valid_26_15 = io_inValid_15 & _T_9821; // @[Switch.scala 30:36:@4268.4]
  assign _T_9824 = io_inAddr_16 == 5'h1a; // @[Switch.scala 30:53:@4270.4]
  assign valid_26_16 = io_inValid_16 & _T_9824; // @[Switch.scala 30:36:@4271.4]
  assign _T_9827 = io_inAddr_17 == 5'h1a; // @[Switch.scala 30:53:@4273.4]
  assign valid_26_17 = io_inValid_17 & _T_9827; // @[Switch.scala 30:36:@4274.4]
  assign _T_9830 = io_inAddr_18 == 5'h1a; // @[Switch.scala 30:53:@4276.4]
  assign valid_26_18 = io_inValid_18 & _T_9830; // @[Switch.scala 30:36:@4277.4]
  assign _T_9833 = io_inAddr_19 == 5'h1a; // @[Switch.scala 30:53:@4279.4]
  assign valid_26_19 = io_inValid_19 & _T_9833; // @[Switch.scala 30:36:@4280.4]
  assign _T_9836 = io_inAddr_20 == 5'h1a; // @[Switch.scala 30:53:@4282.4]
  assign valid_26_20 = io_inValid_20 & _T_9836; // @[Switch.scala 30:36:@4283.4]
  assign _T_9839 = io_inAddr_21 == 5'h1a; // @[Switch.scala 30:53:@4285.4]
  assign valid_26_21 = io_inValid_21 & _T_9839; // @[Switch.scala 30:36:@4286.4]
  assign _T_9842 = io_inAddr_22 == 5'h1a; // @[Switch.scala 30:53:@4288.4]
  assign valid_26_22 = io_inValid_22 & _T_9842; // @[Switch.scala 30:36:@4289.4]
  assign _T_9845 = io_inAddr_23 == 5'h1a; // @[Switch.scala 30:53:@4291.4]
  assign valid_26_23 = io_inValid_23 & _T_9845; // @[Switch.scala 30:36:@4292.4]
  assign _T_9848 = io_inAddr_24 == 5'h1a; // @[Switch.scala 30:53:@4294.4]
  assign valid_26_24 = io_inValid_24 & _T_9848; // @[Switch.scala 30:36:@4295.4]
  assign _T_9851 = io_inAddr_25 == 5'h1a; // @[Switch.scala 30:53:@4297.4]
  assign valid_26_25 = io_inValid_25 & _T_9851; // @[Switch.scala 30:36:@4298.4]
  assign _T_9854 = io_inAddr_26 == 5'h1a; // @[Switch.scala 30:53:@4300.4]
  assign valid_26_26 = io_inValid_26 & _T_9854; // @[Switch.scala 30:36:@4301.4]
  assign _T_9857 = io_inAddr_27 == 5'h1a; // @[Switch.scala 30:53:@4303.4]
  assign valid_26_27 = io_inValid_27 & _T_9857; // @[Switch.scala 30:36:@4304.4]
  assign _T_9860 = io_inAddr_28 == 5'h1a; // @[Switch.scala 30:53:@4306.4]
  assign valid_26_28 = io_inValid_28 & _T_9860; // @[Switch.scala 30:36:@4307.4]
  assign _T_9863 = io_inAddr_29 == 5'h1a; // @[Switch.scala 30:53:@4309.4]
  assign valid_26_29 = io_inValid_29 & _T_9863; // @[Switch.scala 30:36:@4310.4]
  assign _T_9866 = io_inAddr_30 == 5'h1a; // @[Switch.scala 30:53:@4312.4]
  assign valid_26_30 = io_inValid_30 & _T_9866; // @[Switch.scala 30:36:@4313.4]
  assign _T_9869 = io_inAddr_31 == 5'h1a; // @[Switch.scala 30:53:@4315.4]
  assign valid_26_31 = io_inValid_31 & _T_9869; // @[Switch.scala 30:36:@4316.4]
  assign _T_9903 = valid_26_30 ? 5'h1e : 5'h1f; // @[Mux.scala 31:69:@4318.4]
  assign _T_9904 = valid_26_29 ? 5'h1d : _T_9903; // @[Mux.scala 31:69:@4319.4]
  assign _T_9905 = valid_26_28 ? 5'h1c : _T_9904; // @[Mux.scala 31:69:@4320.4]
  assign _T_9906 = valid_26_27 ? 5'h1b : _T_9905; // @[Mux.scala 31:69:@4321.4]
  assign _T_9907 = valid_26_26 ? 5'h1a : _T_9906; // @[Mux.scala 31:69:@4322.4]
  assign _T_9908 = valid_26_25 ? 5'h19 : _T_9907; // @[Mux.scala 31:69:@4323.4]
  assign _T_9909 = valid_26_24 ? 5'h18 : _T_9908; // @[Mux.scala 31:69:@4324.4]
  assign _T_9910 = valid_26_23 ? 5'h17 : _T_9909; // @[Mux.scala 31:69:@4325.4]
  assign _T_9911 = valid_26_22 ? 5'h16 : _T_9910; // @[Mux.scala 31:69:@4326.4]
  assign _T_9912 = valid_26_21 ? 5'h15 : _T_9911; // @[Mux.scala 31:69:@4327.4]
  assign _T_9913 = valid_26_20 ? 5'h14 : _T_9912; // @[Mux.scala 31:69:@4328.4]
  assign _T_9914 = valid_26_19 ? 5'h13 : _T_9913; // @[Mux.scala 31:69:@4329.4]
  assign _T_9915 = valid_26_18 ? 5'h12 : _T_9914; // @[Mux.scala 31:69:@4330.4]
  assign _T_9916 = valid_26_17 ? 5'h11 : _T_9915; // @[Mux.scala 31:69:@4331.4]
  assign _T_9917 = valid_26_16 ? 5'h10 : _T_9916; // @[Mux.scala 31:69:@4332.4]
  assign _T_9918 = valid_26_15 ? 5'hf : _T_9917; // @[Mux.scala 31:69:@4333.4]
  assign _T_9919 = valid_26_14 ? 5'he : _T_9918; // @[Mux.scala 31:69:@4334.4]
  assign _T_9920 = valid_26_13 ? 5'hd : _T_9919; // @[Mux.scala 31:69:@4335.4]
  assign _T_9921 = valid_26_12 ? 5'hc : _T_9920; // @[Mux.scala 31:69:@4336.4]
  assign _T_9922 = valid_26_11 ? 5'hb : _T_9921; // @[Mux.scala 31:69:@4337.4]
  assign _T_9923 = valid_26_10 ? 5'ha : _T_9922; // @[Mux.scala 31:69:@4338.4]
  assign _T_9924 = valid_26_9 ? 5'h9 : _T_9923; // @[Mux.scala 31:69:@4339.4]
  assign _T_9925 = valid_26_8 ? 5'h8 : _T_9924; // @[Mux.scala 31:69:@4340.4]
  assign _T_9926 = valid_26_7 ? 5'h7 : _T_9925; // @[Mux.scala 31:69:@4341.4]
  assign _T_9927 = valid_26_6 ? 5'h6 : _T_9926; // @[Mux.scala 31:69:@4342.4]
  assign _T_9928 = valid_26_5 ? 5'h5 : _T_9927; // @[Mux.scala 31:69:@4343.4]
  assign _T_9929 = valid_26_4 ? 5'h4 : _T_9928; // @[Mux.scala 31:69:@4344.4]
  assign _T_9930 = valid_26_3 ? 5'h3 : _T_9929; // @[Mux.scala 31:69:@4345.4]
  assign _T_9931 = valid_26_2 ? 5'h2 : _T_9930; // @[Mux.scala 31:69:@4346.4]
  assign _T_9932 = valid_26_1 ? 5'h1 : _T_9931; // @[Mux.scala 31:69:@4347.4]
  assign select_26 = valid_26_0 ? 5'h0 : _T_9932; // @[Mux.scala 31:69:@4348.4]
  assign _GEN_833 = 5'h1 == select_26 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@4350.4]
  assign _GEN_834 = 5'h2 == select_26 ? io_inData_2 : _GEN_833; // @[Switch.scala 33:19:@4350.4]
  assign _GEN_835 = 5'h3 == select_26 ? io_inData_3 : _GEN_834; // @[Switch.scala 33:19:@4350.4]
  assign _GEN_836 = 5'h4 == select_26 ? io_inData_4 : _GEN_835; // @[Switch.scala 33:19:@4350.4]
  assign _GEN_837 = 5'h5 == select_26 ? io_inData_5 : _GEN_836; // @[Switch.scala 33:19:@4350.4]
  assign _GEN_838 = 5'h6 == select_26 ? io_inData_6 : _GEN_837; // @[Switch.scala 33:19:@4350.4]
  assign _GEN_839 = 5'h7 == select_26 ? io_inData_7 : _GEN_838; // @[Switch.scala 33:19:@4350.4]
  assign _GEN_840 = 5'h8 == select_26 ? io_inData_8 : _GEN_839; // @[Switch.scala 33:19:@4350.4]
  assign _GEN_841 = 5'h9 == select_26 ? io_inData_9 : _GEN_840; // @[Switch.scala 33:19:@4350.4]
  assign _GEN_842 = 5'ha == select_26 ? io_inData_10 : _GEN_841; // @[Switch.scala 33:19:@4350.4]
  assign _GEN_843 = 5'hb == select_26 ? io_inData_11 : _GEN_842; // @[Switch.scala 33:19:@4350.4]
  assign _GEN_844 = 5'hc == select_26 ? io_inData_12 : _GEN_843; // @[Switch.scala 33:19:@4350.4]
  assign _GEN_845 = 5'hd == select_26 ? io_inData_13 : _GEN_844; // @[Switch.scala 33:19:@4350.4]
  assign _GEN_846 = 5'he == select_26 ? io_inData_14 : _GEN_845; // @[Switch.scala 33:19:@4350.4]
  assign _GEN_847 = 5'hf == select_26 ? io_inData_15 : _GEN_846; // @[Switch.scala 33:19:@4350.4]
  assign _GEN_848 = 5'h10 == select_26 ? io_inData_16 : _GEN_847; // @[Switch.scala 33:19:@4350.4]
  assign _GEN_849 = 5'h11 == select_26 ? io_inData_17 : _GEN_848; // @[Switch.scala 33:19:@4350.4]
  assign _GEN_850 = 5'h12 == select_26 ? io_inData_18 : _GEN_849; // @[Switch.scala 33:19:@4350.4]
  assign _GEN_851 = 5'h13 == select_26 ? io_inData_19 : _GEN_850; // @[Switch.scala 33:19:@4350.4]
  assign _GEN_852 = 5'h14 == select_26 ? io_inData_20 : _GEN_851; // @[Switch.scala 33:19:@4350.4]
  assign _GEN_853 = 5'h15 == select_26 ? io_inData_21 : _GEN_852; // @[Switch.scala 33:19:@4350.4]
  assign _GEN_854 = 5'h16 == select_26 ? io_inData_22 : _GEN_853; // @[Switch.scala 33:19:@4350.4]
  assign _GEN_855 = 5'h17 == select_26 ? io_inData_23 : _GEN_854; // @[Switch.scala 33:19:@4350.4]
  assign _GEN_856 = 5'h18 == select_26 ? io_inData_24 : _GEN_855; // @[Switch.scala 33:19:@4350.4]
  assign _GEN_857 = 5'h19 == select_26 ? io_inData_25 : _GEN_856; // @[Switch.scala 33:19:@4350.4]
  assign _GEN_858 = 5'h1a == select_26 ? io_inData_26 : _GEN_857; // @[Switch.scala 33:19:@4350.4]
  assign _GEN_859 = 5'h1b == select_26 ? io_inData_27 : _GEN_858; // @[Switch.scala 33:19:@4350.4]
  assign _GEN_860 = 5'h1c == select_26 ? io_inData_28 : _GEN_859; // @[Switch.scala 33:19:@4350.4]
  assign _GEN_861 = 5'h1d == select_26 ? io_inData_29 : _GEN_860; // @[Switch.scala 33:19:@4350.4]
  assign _GEN_862 = 5'h1e == select_26 ? io_inData_30 : _GEN_861; // @[Switch.scala 33:19:@4350.4]
  assign _T_9941 = {valid_26_7,valid_26_6,valid_26_5,valid_26_4,valid_26_3,valid_26_2,valid_26_1,valid_26_0}; // @[Switch.scala 34:32:@4357.4]
  assign _T_9949 = {valid_26_15,valid_26_14,valid_26_13,valid_26_12,valid_26_11,valid_26_10,valid_26_9,valid_26_8,_T_9941}; // @[Switch.scala 34:32:@4365.4]
  assign _T_9956 = {valid_26_23,valid_26_22,valid_26_21,valid_26_20,valid_26_19,valid_26_18,valid_26_17,valid_26_16}; // @[Switch.scala 34:32:@4372.4]
  assign _T_9965 = {valid_26_31,valid_26_30,valid_26_29,valid_26_28,valid_26_27,valid_26_26,valid_26_25,valid_26_24,_T_9956,_T_9949}; // @[Switch.scala 34:32:@4381.4]
  assign _T_9969 = io_inAddr_0 == 5'h1b; // @[Switch.scala 30:53:@4384.4]
  assign valid_27_0 = io_inValid_0 & _T_9969; // @[Switch.scala 30:36:@4385.4]
  assign _T_9972 = io_inAddr_1 == 5'h1b; // @[Switch.scala 30:53:@4387.4]
  assign valid_27_1 = io_inValid_1 & _T_9972; // @[Switch.scala 30:36:@4388.4]
  assign _T_9975 = io_inAddr_2 == 5'h1b; // @[Switch.scala 30:53:@4390.4]
  assign valid_27_2 = io_inValid_2 & _T_9975; // @[Switch.scala 30:36:@4391.4]
  assign _T_9978 = io_inAddr_3 == 5'h1b; // @[Switch.scala 30:53:@4393.4]
  assign valid_27_3 = io_inValid_3 & _T_9978; // @[Switch.scala 30:36:@4394.4]
  assign _T_9981 = io_inAddr_4 == 5'h1b; // @[Switch.scala 30:53:@4396.4]
  assign valid_27_4 = io_inValid_4 & _T_9981; // @[Switch.scala 30:36:@4397.4]
  assign _T_9984 = io_inAddr_5 == 5'h1b; // @[Switch.scala 30:53:@4399.4]
  assign valid_27_5 = io_inValid_5 & _T_9984; // @[Switch.scala 30:36:@4400.4]
  assign _T_9987 = io_inAddr_6 == 5'h1b; // @[Switch.scala 30:53:@4402.4]
  assign valid_27_6 = io_inValid_6 & _T_9987; // @[Switch.scala 30:36:@4403.4]
  assign _T_9990 = io_inAddr_7 == 5'h1b; // @[Switch.scala 30:53:@4405.4]
  assign valid_27_7 = io_inValid_7 & _T_9990; // @[Switch.scala 30:36:@4406.4]
  assign _T_9993 = io_inAddr_8 == 5'h1b; // @[Switch.scala 30:53:@4408.4]
  assign valid_27_8 = io_inValid_8 & _T_9993; // @[Switch.scala 30:36:@4409.4]
  assign _T_9996 = io_inAddr_9 == 5'h1b; // @[Switch.scala 30:53:@4411.4]
  assign valid_27_9 = io_inValid_9 & _T_9996; // @[Switch.scala 30:36:@4412.4]
  assign _T_9999 = io_inAddr_10 == 5'h1b; // @[Switch.scala 30:53:@4414.4]
  assign valid_27_10 = io_inValid_10 & _T_9999; // @[Switch.scala 30:36:@4415.4]
  assign _T_10002 = io_inAddr_11 == 5'h1b; // @[Switch.scala 30:53:@4417.4]
  assign valid_27_11 = io_inValid_11 & _T_10002; // @[Switch.scala 30:36:@4418.4]
  assign _T_10005 = io_inAddr_12 == 5'h1b; // @[Switch.scala 30:53:@4420.4]
  assign valid_27_12 = io_inValid_12 & _T_10005; // @[Switch.scala 30:36:@4421.4]
  assign _T_10008 = io_inAddr_13 == 5'h1b; // @[Switch.scala 30:53:@4423.4]
  assign valid_27_13 = io_inValid_13 & _T_10008; // @[Switch.scala 30:36:@4424.4]
  assign _T_10011 = io_inAddr_14 == 5'h1b; // @[Switch.scala 30:53:@4426.4]
  assign valid_27_14 = io_inValid_14 & _T_10011; // @[Switch.scala 30:36:@4427.4]
  assign _T_10014 = io_inAddr_15 == 5'h1b; // @[Switch.scala 30:53:@4429.4]
  assign valid_27_15 = io_inValid_15 & _T_10014; // @[Switch.scala 30:36:@4430.4]
  assign _T_10017 = io_inAddr_16 == 5'h1b; // @[Switch.scala 30:53:@4432.4]
  assign valid_27_16 = io_inValid_16 & _T_10017; // @[Switch.scala 30:36:@4433.4]
  assign _T_10020 = io_inAddr_17 == 5'h1b; // @[Switch.scala 30:53:@4435.4]
  assign valid_27_17 = io_inValid_17 & _T_10020; // @[Switch.scala 30:36:@4436.4]
  assign _T_10023 = io_inAddr_18 == 5'h1b; // @[Switch.scala 30:53:@4438.4]
  assign valid_27_18 = io_inValid_18 & _T_10023; // @[Switch.scala 30:36:@4439.4]
  assign _T_10026 = io_inAddr_19 == 5'h1b; // @[Switch.scala 30:53:@4441.4]
  assign valid_27_19 = io_inValid_19 & _T_10026; // @[Switch.scala 30:36:@4442.4]
  assign _T_10029 = io_inAddr_20 == 5'h1b; // @[Switch.scala 30:53:@4444.4]
  assign valid_27_20 = io_inValid_20 & _T_10029; // @[Switch.scala 30:36:@4445.4]
  assign _T_10032 = io_inAddr_21 == 5'h1b; // @[Switch.scala 30:53:@4447.4]
  assign valid_27_21 = io_inValid_21 & _T_10032; // @[Switch.scala 30:36:@4448.4]
  assign _T_10035 = io_inAddr_22 == 5'h1b; // @[Switch.scala 30:53:@4450.4]
  assign valid_27_22 = io_inValid_22 & _T_10035; // @[Switch.scala 30:36:@4451.4]
  assign _T_10038 = io_inAddr_23 == 5'h1b; // @[Switch.scala 30:53:@4453.4]
  assign valid_27_23 = io_inValid_23 & _T_10038; // @[Switch.scala 30:36:@4454.4]
  assign _T_10041 = io_inAddr_24 == 5'h1b; // @[Switch.scala 30:53:@4456.4]
  assign valid_27_24 = io_inValid_24 & _T_10041; // @[Switch.scala 30:36:@4457.4]
  assign _T_10044 = io_inAddr_25 == 5'h1b; // @[Switch.scala 30:53:@4459.4]
  assign valid_27_25 = io_inValid_25 & _T_10044; // @[Switch.scala 30:36:@4460.4]
  assign _T_10047 = io_inAddr_26 == 5'h1b; // @[Switch.scala 30:53:@4462.4]
  assign valid_27_26 = io_inValid_26 & _T_10047; // @[Switch.scala 30:36:@4463.4]
  assign _T_10050 = io_inAddr_27 == 5'h1b; // @[Switch.scala 30:53:@4465.4]
  assign valid_27_27 = io_inValid_27 & _T_10050; // @[Switch.scala 30:36:@4466.4]
  assign _T_10053 = io_inAddr_28 == 5'h1b; // @[Switch.scala 30:53:@4468.4]
  assign valid_27_28 = io_inValid_28 & _T_10053; // @[Switch.scala 30:36:@4469.4]
  assign _T_10056 = io_inAddr_29 == 5'h1b; // @[Switch.scala 30:53:@4471.4]
  assign valid_27_29 = io_inValid_29 & _T_10056; // @[Switch.scala 30:36:@4472.4]
  assign _T_10059 = io_inAddr_30 == 5'h1b; // @[Switch.scala 30:53:@4474.4]
  assign valid_27_30 = io_inValid_30 & _T_10059; // @[Switch.scala 30:36:@4475.4]
  assign _T_10062 = io_inAddr_31 == 5'h1b; // @[Switch.scala 30:53:@4477.4]
  assign valid_27_31 = io_inValid_31 & _T_10062; // @[Switch.scala 30:36:@4478.4]
  assign _T_10096 = valid_27_30 ? 5'h1e : 5'h1f; // @[Mux.scala 31:69:@4480.4]
  assign _T_10097 = valid_27_29 ? 5'h1d : _T_10096; // @[Mux.scala 31:69:@4481.4]
  assign _T_10098 = valid_27_28 ? 5'h1c : _T_10097; // @[Mux.scala 31:69:@4482.4]
  assign _T_10099 = valid_27_27 ? 5'h1b : _T_10098; // @[Mux.scala 31:69:@4483.4]
  assign _T_10100 = valid_27_26 ? 5'h1a : _T_10099; // @[Mux.scala 31:69:@4484.4]
  assign _T_10101 = valid_27_25 ? 5'h19 : _T_10100; // @[Mux.scala 31:69:@4485.4]
  assign _T_10102 = valid_27_24 ? 5'h18 : _T_10101; // @[Mux.scala 31:69:@4486.4]
  assign _T_10103 = valid_27_23 ? 5'h17 : _T_10102; // @[Mux.scala 31:69:@4487.4]
  assign _T_10104 = valid_27_22 ? 5'h16 : _T_10103; // @[Mux.scala 31:69:@4488.4]
  assign _T_10105 = valid_27_21 ? 5'h15 : _T_10104; // @[Mux.scala 31:69:@4489.4]
  assign _T_10106 = valid_27_20 ? 5'h14 : _T_10105; // @[Mux.scala 31:69:@4490.4]
  assign _T_10107 = valid_27_19 ? 5'h13 : _T_10106; // @[Mux.scala 31:69:@4491.4]
  assign _T_10108 = valid_27_18 ? 5'h12 : _T_10107; // @[Mux.scala 31:69:@4492.4]
  assign _T_10109 = valid_27_17 ? 5'h11 : _T_10108; // @[Mux.scala 31:69:@4493.4]
  assign _T_10110 = valid_27_16 ? 5'h10 : _T_10109; // @[Mux.scala 31:69:@4494.4]
  assign _T_10111 = valid_27_15 ? 5'hf : _T_10110; // @[Mux.scala 31:69:@4495.4]
  assign _T_10112 = valid_27_14 ? 5'he : _T_10111; // @[Mux.scala 31:69:@4496.4]
  assign _T_10113 = valid_27_13 ? 5'hd : _T_10112; // @[Mux.scala 31:69:@4497.4]
  assign _T_10114 = valid_27_12 ? 5'hc : _T_10113; // @[Mux.scala 31:69:@4498.4]
  assign _T_10115 = valid_27_11 ? 5'hb : _T_10114; // @[Mux.scala 31:69:@4499.4]
  assign _T_10116 = valid_27_10 ? 5'ha : _T_10115; // @[Mux.scala 31:69:@4500.4]
  assign _T_10117 = valid_27_9 ? 5'h9 : _T_10116; // @[Mux.scala 31:69:@4501.4]
  assign _T_10118 = valid_27_8 ? 5'h8 : _T_10117; // @[Mux.scala 31:69:@4502.4]
  assign _T_10119 = valid_27_7 ? 5'h7 : _T_10118; // @[Mux.scala 31:69:@4503.4]
  assign _T_10120 = valid_27_6 ? 5'h6 : _T_10119; // @[Mux.scala 31:69:@4504.4]
  assign _T_10121 = valid_27_5 ? 5'h5 : _T_10120; // @[Mux.scala 31:69:@4505.4]
  assign _T_10122 = valid_27_4 ? 5'h4 : _T_10121; // @[Mux.scala 31:69:@4506.4]
  assign _T_10123 = valid_27_3 ? 5'h3 : _T_10122; // @[Mux.scala 31:69:@4507.4]
  assign _T_10124 = valid_27_2 ? 5'h2 : _T_10123; // @[Mux.scala 31:69:@4508.4]
  assign _T_10125 = valid_27_1 ? 5'h1 : _T_10124; // @[Mux.scala 31:69:@4509.4]
  assign select_27 = valid_27_0 ? 5'h0 : _T_10125; // @[Mux.scala 31:69:@4510.4]
  assign _GEN_865 = 5'h1 == select_27 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@4512.4]
  assign _GEN_866 = 5'h2 == select_27 ? io_inData_2 : _GEN_865; // @[Switch.scala 33:19:@4512.4]
  assign _GEN_867 = 5'h3 == select_27 ? io_inData_3 : _GEN_866; // @[Switch.scala 33:19:@4512.4]
  assign _GEN_868 = 5'h4 == select_27 ? io_inData_4 : _GEN_867; // @[Switch.scala 33:19:@4512.4]
  assign _GEN_869 = 5'h5 == select_27 ? io_inData_5 : _GEN_868; // @[Switch.scala 33:19:@4512.4]
  assign _GEN_870 = 5'h6 == select_27 ? io_inData_6 : _GEN_869; // @[Switch.scala 33:19:@4512.4]
  assign _GEN_871 = 5'h7 == select_27 ? io_inData_7 : _GEN_870; // @[Switch.scala 33:19:@4512.4]
  assign _GEN_872 = 5'h8 == select_27 ? io_inData_8 : _GEN_871; // @[Switch.scala 33:19:@4512.4]
  assign _GEN_873 = 5'h9 == select_27 ? io_inData_9 : _GEN_872; // @[Switch.scala 33:19:@4512.4]
  assign _GEN_874 = 5'ha == select_27 ? io_inData_10 : _GEN_873; // @[Switch.scala 33:19:@4512.4]
  assign _GEN_875 = 5'hb == select_27 ? io_inData_11 : _GEN_874; // @[Switch.scala 33:19:@4512.4]
  assign _GEN_876 = 5'hc == select_27 ? io_inData_12 : _GEN_875; // @[Switch.scala 33:19:@4512.4]
  assign _GEN_877 = 5'hd == select_27 ? io_inData_13 : _GEN_876; // @[Switch.scala 33:19:@4512.4]
  assign _GEN_878 = 5'he == select_27 ? io_inData_14 : _GEN_877; // @[Switch.scala 33:19:@4512.4]
  assign _GEN_879 = 5'hf == select_27 ? io_inData_15 : _GEN_878; // @[Switch.scala 33:19:@4512.4]
  assign _GEN_880 = 5'h10 == select_27 ? io_inData_16 : _GEN_879; // @[Switch.scala 33:19:@4512.4]
  assign _GEN_881 = 5'h11 == select_27 ? io_inData_17 : _GEN_880; // @[Switch.scala 33:19:@4512.4]
  assign _GEN_882 = 5'h12 == select_27 ? io_inData_18 : _GEN_881; // @[Switch.scala 33:19:@4512.4]
  assign _GEN_883 = 5'h13 == select_27 ? io_inData_19 : _GEN_882; // @[Switch.scala 33:19:@4512.4]
  assign _GEN_884 = 5'h14 == select_27 ? io_inData_20 : _GEN_883; // @[Switch.scala 33:19:@4512.4]
  assign _GEN_885 = 5'h15 == select_27 ? io_inData_21 : _GEN_884; // @[Switch.scala 33:19:@4512.4]
  assign _GEN_886 = 5'h16 == select_27 ? io_inData_22 : _GEN_885; // @[Switch.scala 33:19:@4512.4]
  assign _GEN_887 = 5'h17 == select_27 ? io_inData_23 : _GEN_886; // @[Switch.scala 33:19:@4512.4]
  assign _GEN_888 = 5'h18 == select_27 ? io_inData_24 : _GEN_887; // @[Switch.scala 33:19:@4512.4]
  assign _GEN_889 = 5'h19 == select_27 ? io_inData_25 : _GEN_888; // @[Switch.scala 33:19:@4512.4]
  assign _GEN_890 = 5'h1a == select_27 ? io_inData_26 : _GEN_889; // @[Switch.scala 33:19:@4512.4]
  assign _GEN_891 = 5'h1b == select_27 ? io_inData_27 : _GEN_890; // @[Switch.scala 33:19:@4512.4]
  assign _GEN_892 = 5'h1c == select_27 ? io_inData_28 : _GEN_891; // @[Switch.scala 33:19:@4512.4]
  assign _GEN_893 = 5'h1d == select_27 ? io_inData_29 : _GEN_892; // @[Switch.scala 33:19:@4512.4]
  assign _GEN_894 = 5'h1e == select_27 ? io_inData_30 : _GEN_893; // @[Switch.scala 33:19:@4512.4]
  assign _T_10134 = {valid_27_7,valid_27_6,valid_27_5,valid_27_4,valid_27_3,valid_27_2,valid_27_1,valid_27_0}; // @[Switch.scala 34:32:@4519.4]
  assign _T_10142 = {valid_27_15,valid_27_14,valid_27_13,valid_27_12,valid_27_11,valid_27_10,valid_27_9,valid_27_8,_T_10134}; // @[Switch.scala 34:32:@4527.4]
  assign _T_10149 = {valid_27_23,valid_27_22,valid_27_21,valid_27_20,valid_27_19,valid_27_18,valid_27_17,valid_27_16}; // @[Switch.scala 34:32:@4534.4]
  assign _T_10158 = {valid_27_31,valid_27_30,valid_27_29,valid_27_28,valid_27_27,valid_27_26,valid_27_25,valid_27_24,_T_10149,_T_10142}; // @[Switch.scala 34:32:@4543.4]
  assign _T_10162 = io_inAddr_0 == 5'h1c; // @[Switch.scala 30:53:@4546.4]
  assign valid_28_0 = io_inValid_0 & _T_10162; // @[Switch.scala 30:36:@4547.4]
  assign _T_10165 = io_inAddr_1 == 5'h1c; // @[Switch.scala 30:53:@4549.4]
  assign valid_28_1 = io_inValid_1 & _T_10165; // @[Switch.scala 30:36:@4550.4]
  assign _T_10168 = io_inAddr_2 == 5'h1c; // @[Switch.scala 30:53:@4552.4]
  assign valid_28_2 = io_inValid_2 & _T_10168; // @[Switch.scala 30:36:@4553.4]
  assign _T_10171 = io_inAddr_3 == 5'h1c; // @[Switch.scala 30:53:@4555.4]
  assign valid_28_3 = io_inValid_3 & _T_10171; // @[Switch.scala 30:36:@4556.4]
  assign _T_10174 = io_inAddr_4 == 5'h1c; // @[Switch.scala 30:53:@4558.4]
  assign valid_28_4 = io_inValid_4 & _T_10174; // @[Switch.scala 30:36:@4559.4]
  assign _T_10177 = io_inAddr_5 == 5'h1c; // @[Switch.scala 30:53:@4561.4]
  assign valid_28_5 = io_inValid_5 & _T_10177; // @[Switch.scala 30:36:@4562.4]
  assign _T_10180 = io_inAddr_6 == 5'h1c; // @[Switch.scala 30:53:@4564.4]
  assign valid_28_6 = io_inValid_6 & _T_10180; // @[Switch.scala 30:36:@4565.4]
  assign _T_10183 = io_inAddr_7 == 5'h1c; // @[Switch.scala 30:53:@4567.4]
  assign valid_28_7 = io_inValid_7 & _T_10183; // @[Switch.scala 30:36:@4568.4]
  assign _T_10186 = io_inAddr_8 == 5'h1c; // @[Switch.scala 30:53:@4570.4]
  assign valid_28_8 = io_inValid_8 & _T_10186; // @[Switch.scala 30:36:@4571.4]
  assign _T_10189 = io_inAddr_9 == 5'h1c; // @[Switch.scala 30:53:@4573.4]
  assign valid_28_9 = io_inValid_9 & _T_10189; // @[Switch.scala 30:36:@4574.4]
  assign _T_10192 = io_inAddr_10 == 5'h1c; // @[Switch.scala 30:53:@4576.4]
  assign valid_28_10 = io_inValid_10 & _T_10192; // @[Switch.scala 30:36:@4577.4]
  assign _T_10195 = io_inAddr_11 == 5'h1c; // @[Switch.scala 30:53:@4579.4]
  assign valid_28_11 = io_inValid_11 & _T_10195; // @[Switch.scala 30:36:@4580.4]
  assign _T_10198 = io_inAddr_12 == 5'h1c; // @[Switch.scala 30:53:@4582.4]
  assign valid_28_12 = io_inValid_12 & _T_10198; // @[Switch.scala 30:36:@4583.4]
  assign _T_10201 = io_inAddr_13 == 5'h1c; // @[Switch.scala 30:53:@4585.4]
  assign valid_28_13 = io_inValid_13 & _T_10201; // @[Switch.scala 30:36:@4586.4]
  assign _T_10204 = io_inAddr_14 == 5'h1c; // @[Switch.scala 30:53:@4588.4]
  assign valid_28_14 = io_inValid_14 & _T_10204; // @[Switch.scala 30:36:@4589.4]
  assign _T_10207 = io_inAddr_15 == 5'h1c; // @[Switch.scala 30:53:@4591.4]
  assign valid_28_15 = io_inValid_15 & _T_10207; // @[Switch.scala 30:36:@4592.4]
  assign _T_10210 = io_inAddr_16 == 5'h1c; // @[Switch.scala 30:53:@4594.4]
  assign valid_28_16 = io_inValid_16 & _T_10210; // @[Switch.scala 30:36:@4595.4]
  assign _T_10213 = io_inAddr_17 == 5'h1c; // @[Switch.scala 30:53:@4597.4]
  assign valid_28_17 = io_inValid_17 & _T_10213; // @[Switch.scala 30:36:@4598.4]
  assign _T_10216 = io_inAddr_18 == 5'h1c; // @[Switch.scala 30:53:@4600.4]
  assign valid_28_18 = io_inValid_18 & _T_10216; // @[Switch.scala 30:36:@4601.4]
  assign _T_10219 = io_inAddr_19 == 5'h1c; // @[Switch.scala 30:53:@4603.4]
  assign valid_28_19 = io_inValid_19 & _T_10219; // @[Switch.scala 30:36:@4604.4]
  assign _T_10222 = io_inAddr_20 == 5'h1c; // @[Switch.scala 30:53:@4606.4]
  assign valid_28_20 = io_inValid_20 & _T_10222; // @[Switch.scala 30:36:@4607.4]
  assign _T_10225 = io_inAddr_21 == 5'h1c; // @[Switch.scala 30:53:@4609.4]
  assign valid_28_21 = io_inValid_21 & _T_10225; // @[Switch.scala 30:36:@4610.4]
  assign _T_10228 = io_inAddr_22 == 5'h1c; // @[Switch.scala 30:53:@4612.4]
  assign valid_28_22 = io_inValid_22 & _T_10228; // @[Switch.scala 30:36:@4613.4]
  assign _T_10231 = io_inAddr_23 == 5'h1c; // @[Switch.scala 30:53:@4615.4]
  assign valid_28_23 = io_inValid_23 & _T_10231; // @[Switch.scala 30:36:@4616.4]
  assign _T_10234 = io_inAddr_24 == 5'h1c; // @[Switch.scala 30:53:@4618.4]
  assign valid_28_24 = io_inValid_24 & _T_10234; // @[Switch.scala 30:36:@4619.4]
  assign _T_10237 = io_inAddr_25 == 5'h1c; // @[Switch.scala 30:53:@4621.4]
  assign valid_28_25 = io_inValid_25 & _T_10237; // @[Switch.scala 30:36:@4622.4]
  assign _T_10240 = io_inAddr_26 == 5'h1c; // @[Switch.scala 30:53:@4624.4]
  assign valid_28_26 = io_inValid_26 & _T_10240; // @[Switch.scala 30:36:@4625.4]
  assign _T_10243 = io_inAddr_27 == 5'h1c; // @[Switch.scala 30:53:@4627.4]
  assign valid_28_27 = io_inValid_27 & _T_10243; // @[Switch.scala 30:36:@4628.4]
  assign _T_10246 = io_inAddr_28 == 5'h1c; // @[Switch.scala 30:53:@4630.4]
  assign valid_28_28 = io_inValid_28 & _T_10246; // @[Switch.scala 30:36:@4631.4]
  assign _T_10249 = io_inAddr_29 == 5'h1c; // @[Switch.scala 30:53:@4633.4]
  assign valid_28_29 = io_inValid_29 & _T_10249; // @[Switch.scala 30:36:@4634.4]
  assign _T_10252 = io_inAddr_30 == 5'h1c; // @[Switch.scala 30:53:@4636.4]
  assign valid_28_30 = io_inValid_30 & _T_10252; // @[Switch.scala 30:36:@4637.4]
  assign _T_10255 = io_inAddr_31 == 5'h1c; // @[Switch.scala 30:53:@4639.4]
  assign valid_28_31 = io_inValid_31 & _T_10255; // @[Switch.scala 30:36:@4640.4]
  assign _T_10289 = valid_28_30 ? 5'h1e : 5'h1f; // @[Mux.scala 31:69:@4642.4]
  assign _T_10290 = valid_28_29 ? 5'h1d : _T_10289; // @[Mux.scala 31:69:@4643.4]
  assign _T_10291 = valid_28_28 ? 5'h1c : _T_10290; // @[Mux.scala 31:69:@4644.4]
  assign _T_10292 = valid_28_27 ? 5'h1b : _T_10291; // @[Mux.scala 31:69:@4645.4]
  assign _T_10293 = valid_28_26 ? 5'h1a : _T_10292; // @[Mux.scala 31:69:@4646.4]
  assign _T_10294 = valid_28_25 ? 5'h19 : _T_10293; // @[Mux.scala 31:69:@4647.4]
  assign _T_10295 = valid_28_24 ? 5'h18 : _T_10294; // @[Mux.scala 31:69:@4648.4]
  assign _T_10296 = valid_28_23 ? 5'h17 : _T_10295; // @[Mux.scala 31:69:@4649.4]
  assign _T_10297 = valid_28_22 ? 5'h16 : _T_10296; // @[Mux.scala 31:69:@4650.4]
  assign _T_10298 = valid_28_21 ? 5'h15 : _T_10297; // @[Mux.scala 31:69:@4651.4]
  assign _T_10299 = valid_28_20 ? 5'h14 : _T_10298; // @[Mux.scala 31:69:@4652.4]
  assign _T_10300 = valid_28_19 ? 5'h13 : _T_10299; // @[Mux.scala 31:69:@4653.4]
  assign _T_10301 = valid_28_18 ? 5'h12 : _T_10300; // @[Mux.scala 31:69:@4654.4]
  assign _T_10302 = valid_28_17 ? 5'h11 : _T_10301; // @[Mux.scala 31:69:@4655.4]
  assign _T_10303 = valid_28_16 ? 5'h10 : _T_10302; // @[Mux.scala 31:69:@4656.4]
  assign _T_10304 = valid_28_15 ? 5'hf : _T_10303; // @[Mux.scala 31:69:@4657.4]
  assign _T_10305 = valid_28_14 ? 5'he : _T_10304; // @[Mux.scala 31:69:@4658.4]
  assign _T_10306 = valid_28_13 ? 5'hd : _T_10305; // @[Mux.scala 31:69:@4659.4]
  assign _T_10307 = valid_28_12 ? 5'hc : _T_10306; // @[Mux.scala 31:69:@4660.4]
  assign _T_10308 = valid_28_11 ? 5'hb : _T_10307; // @[Mux.scala 31:69:@4661.4]
  assign _T_10309 = valid_28_10 ? 5'ha : _T_10308; // @[Mux.scala 31:69:@4662.4]
  assign _T_10310 = valid_28_9 ? 5'h9 : _T_10309; // @[Mux.scala 31:69:@4663.4]
  assign _T_10311 = valid_28_8 ? 5'h8 : _T_10310; // @[Mux.scala 31:69:@4664.4]
  assign _T_10312 = valid_28_7 ? 5'h7 : _T_10311; // @[Mux.scala 31:69:@4665.4]
  assign _T_10313 = valid_28_6 ? 5'h6 : _T_10312; // @[Mux.scala 31:69:@4666.4]
  assign _T_10314 = valid_28_5 ? 5'h5 : _T_10313; // @[Mux.scala 31:69:@4667.4]
  assign _T_10315 = valid_28_4 ? 5'h4 : _T_10314; // @[Mux.scala 31:69:@4668.4]
  assign _T_10316 = valid_28_3 ? 5'h3 : _T_10315; // @[Mux.scala 31:69:@4669.4]
  assign _T_10317 = valid_28_2 ? 5'h2 : _T_10316; // @[Mux.scala 31:69:@4670.4]
  assign _T_10318 = valid_28_1 ? 5'h1 : _T_10317; // @[Mux.scala 31:69:@4671.4]
  assign select_28 = valid_28_0 ? 5'h0 : _T_10318; // @[Mux.scala 31:69:@4672.4]
  assign _GEN_897 = 5'h1 == select_28 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@4674.4]
  assign _GEN_898 = 5'h2 == select_28 ? io_inData_2 : _GEN_897; // @[Switch.scala 33:19:@4674.4]
  assign _GEN_899 = 5'h3 == select_28 ? io_inData_3 : _GEN_898; // @[Switch.scala 33:19:@4674.4]
  assign _GEN_900 = 5'h4 == select_28 ? io_inData_4 : _GEN_899; // @[Switch.scala 33:19:@4674.4]
  assign _GEN_901 = 5'h5 == select_28 ? io_inData_5 : _GEN_900; // @[Switch.scala 33:19:@4674.4]
  assign _GEN_902 = 5'h6 == select_28 ? io_inData_6 : _GEN_901; // @[Switch.scala 33:19:@4674.4]
  assign _GEN_903 = 5'h7 == select_28 ? io_inData_7 : _GEN_902; // @[Switch.scala 33:19:@4674.4]
  assign _GEN_904 = 5'h8 == select_28 ? io_inData_8 : _GEN_903; // @[Switch.scala 33:19:@4674.4]
  assign _GEN_905 = 5'h9 == select_28 ? io_inData_9 : _GEN_904; // @[Switch.scala 33:19:@4674.4]
  assign _GEN_906 = 5'ha == select_28 ? io_inData_10 : _GEN_905; // @[Switch.scala 33:19:@4674.4]
  assign _GEN_907 = 5'hb == select_28 ? io_inData_11 : _GEN_906; // @[Switch.scala 33:19:@4674.4]
  assign _GEN_908 = 5'hc == select_28 ? io_inData_12 : _GEN_907; // @[Switch.scala 33:19:@4674.4]
  assign _GEN_909 = 5'hd == select_28 ? io_inData_13 : _GEN_908; // @[Switch.scala 33:19:@4674.4]
  assign _GEN_910 = 5'he == select_28 ? io_inData_14 : _GEN_909; // @[Switch.scala 33:19:@4674.4]
  assign _GEN_911 = 5'hf == select_28 ? io_inData_15 : _GEN_910; // @[Switch.scala 33:19:@4674.4]
  assign _GEN_912 = 5'h10 == select_28 ? io_inData_16 : _GEN_911; // @[Switch.scala 33:19:@4674.4]
  assign _GEN_913 = 5'h11 == select_28 ? io_inData_17 : _GEN_912; // @[Switch.scala 33:19:@4674.4]
  assign _GEN_914 = 5'h12 == select_28 ? io_inData_18 : _GEN_913; // @[Switch.scala 33:19:@4674.4]
  assign _GEN_915 = 5'h13 == select_28 ? io_inData_19 : _GEN_914; // @[Switch.scala 33:19:@4674.4]
  assign _GEN_916 = 5'h14 == select_28 ? io_inData_20 : _GEN_915; // @[Switch.scala 33:19:@4674.4]
  assign _GEN_917 = 5'h15 == select_28 ? io_inData_21 : _GEN_916; // @[Switch.scala 33:19:@4674.4]
  assign _GEN_918 = 5'h16 == select_28 ? io_inData_22 : _GEN_917; // @[Switch.scala 33:19:@4674.4]
  assign _GEN_919 = 5'h17 == select_28 ? io_inData_23 : _GEN_918; // @[Switch.scala 33:19:@4674.4]
  assign _GEN_920 = 5'h18 == select_28 ? io_inData_24 : _GEN_919; // @[Switch.scala 33:19:@4674.4]
  assign _GEN_921 = 5'h19 == select_28 ? io_inData_25 : _GEN_920; // @[Switch.scala 33:19:@4674.4]
  assign _GEN_922 = 5'h1a == select_28 ? io_inData_26 : _GEN_921; // @[Switch.scala 33:19:@4674.4]
  assign _GEN_923 = 5'h1b == select_28 ? io_inData_27 : _GEN_922; // @[Switch.scala 33:19:@4674.4]
  assign _GEN_924 = 5'h1c == select_28 ? io_inData_28 : _GEN_923; // @[Switch.scala 33:19:@4674.4]
  assign _GEN_925 = 5'h1d == select_28 ? io_inData_29 : _GEN_924; // @[Switch.scala 33:19:@4674.4]
  assign _GEN_926 = 5'h1e == select_28 ? io_inData_30 : _GEN_925; // @[Switch.scala 33:19:@4674.4]
  assign _T_10327 = {valid_28_7,valid_28_6,valid_28_5,valid_28_4,valid_28_3,valid_28_2,valid_28_1,valid_28_0}; // @[Switch.scala 34:32:@4681.4]
  assign _T_10335 = {valid_28_15,valid_28_14,valid_28_13,valid_28_12,valid_28_11,valid_28_10,valid_28_9,valid_28_8,_T_10327}; // @[Switch.scala 34:32:@4689.4]
  assign _T_10342 = {valid_28_23,valid_28_22,valid_28_21,valid_28_20,valid_28_19,valid_28_18,valid_28_17,valid_28_16}; // @[Switch.scala 34:32:@4696.4]
  assign _T_10351 = {valid_28_31,valid_28_30,valid_28_29,valid_28_28,valid_28_27,valid_28_26,valid_28_25,valid_28_24,_T_10342,_T_10335}; // @[Switch.scala 34:32:@4705.4]
  assign _T_10355 = io_inAddr_0 == 5'h1d; // @[Switch.scala 30:53:@4708.4]
  assign valid_29_0 = io_inValid_0 & _T_10355; // @[Switch.scala 30:36:@4709.4]
  assign _T_10358 = io_inAddr_1 == 5'h1d; // @[Switch.scala 30:53:@4711.4]
  assign valid_29_1 = io_inValid_1 & _T_10358; // @[Switch.scala 30:36:@4712.4]
  assign _T_10361 = io_inAddr_2 == 5'h1d; // @[Switch.scala 30:53:@4714.4]
  assign valid_29_2 = io_inValid_2 & _T_10361; // @[Switch.scala 30:36:@4715.4]
  assign _T_10364 = io_inAddr_3 == 5'h1d; // @[Switch.scala 30:53:@4717.4]
  assign valid_29_3 = io_inValid_3 & _T_10364; // @[Switch.scala 30:36:@4718.4]
  assign _T_10367 = io_inAddr_4 == 5'h1d; // @[Switch.scala 30:53:@4720.4]
  assign valid_29_4 = io_inValid_4 & _T_10367; // @[Switch.scala 30:36:@4721.4]
  assign _T_10370 = io_inAddr_5 == 5'h1d; // @[Switch.scala 30:53:@4723.4]
  assign valid_29_5 = io_inValid_5 & _T_10370; // @[Switch.scala 30:36:@4724.4]
  assign _T_10373 = io_inAddr_6 == 5'h1d; // @[Switch.scala 30:53:@4726.4]
  assign valid_29_6 = io_inValid_6 & _T_10373; // @[Switch.scala 30:36:@4727.4]
  assign _T_10376 = io_inAddr_7 == 5'h1d; // @[Switch.scala 30:53:@4729.4]
  assign valid_29_7 = io_inValid_7 & _T_10376; // @[Switch.scala 30:36:@4730.4]
  assign _T_10379 = io_inAddr_8 == 5'h1d; // @[Switch.scala 30:53:@4732.4]
  assign valid_29_8 = io_inValid_8 & _T_10379; // @[Switch.scala 30:36:@4733.4]
  assign _T_10382 = io_inAddr_9 == 5'h1d; // @[Switch.scala 30:53:@4735.4]
  assign valid_29_9 = io_inValid_9 & _T_10382; // @[Switch.scala 30:36:@4736.4]
  assign _T_10385 = io_inAddr_10 == 5'h1d; // @[Switch.scala 30:53:@4738.4]
  assign valid_29_10 = io_inValid_10 & _T_10385; // @[Switch.scala 30:36:@4739.4]
  assign _T_10388 = io_inAddr_11 == 5'h1d; // @[Switch.scala 30:53:@4741.4]
  assign valid_29_11 = io_inValid_11 & _T_10388; // @[Switch.scala 30:36:@4742.4]
  assign _T_10391 = io_inAddr_12 == 5'h1d; // @[Switch.scala 30:53:@4744.4]
  assign valid_29_12 = io_inValid_12 & _T_10391; // @[Switch.scala 30:36:@4745.4]
  assign _T_10394 = io_inAddr_13 == 5'h1d; // @[Switch.scala 30:53:@4747.4]
  assign valid_29_13 = io_inValid_13 & _T_10394; // @[Switch.scala 30:36:@4748.4]
  assign _T_10397 = io_inAddr_14 == 5'h1d; // @[Switch.scala 30:53:@4750.4]
  assign valid_29_14 = io_inValid_14 & _T_10397; // @[Switch.scala 30:36:@4751.4]
  assign _T_10400 = io_inAddr_15 == 5'h1d; // @[Switch.scala 30:53:@4753.4]
  assign valid_29_15 = io_inValid_15 & _T_10400; // @[Switch.scala 30:36:@4754.4]
  assign _T_10403 = io_inAddr_16 == 5'h1d; // @[Switch.scala 30:53:@4756.4]
  assign valid_29_16 = io_inValid_16 & _T_10403; // @[Switch.scala 30:36:@4757.4]
  assign _T_10406 = io_inAddr_17 == 5'h1d; // @[Switch.scala 30:53:@4759.4]
  assign valid_29_17 = io_inValid_17 & _T_10406; // @[Switch.scala 30:36:@4760.4]
  assign _T_10409 = io_inAddr_18 == 5'h1d; // @[Switch.scala 30:53:@4762.4]
  assign valid_29_18 = io_inValid_18 & _T_10409; // @[Switch.scala 30:36:@4763.4]
  assign _T_10412 = io_inAddr_19 == 5'h1d; // @[Switch.scala 30:53:@4765.4]
  assign valid_29_19 = io_inValid_19 & _T_10412; // @[Switch.scala 30:36:@4766.4]
  assign _T_10415 = io_inAddr_20 == 5'h1d; // @[Switch.scala 30:53:@4768.4]
  assign valid_29_20 = io_inValid_20 & _T_10415; // @[Switch.scala 30:36:@4769.4]
  assign _T_10418 = io_inAddr_21 == 5'h1d; // @[Switch.scala 30:53:@4771.4]
  assign valid_29_21 = io_inValid_21 & _T_10418; // @[Switch.scala 30:36:@4772.4]
  assign _T_10421 = io_inAddr_22 == 5'h1d; // @[Switch.scala 30:53:@4774.4]
  assign valid_29_22 = io_inValid_22 & _T_10421; // @[Switch.scala 30:36:@4775.4]
  assign _T_10424 = io_inAddr_23 == 5'h1d; // @[Switch.scala 30:53:@4777.4]
  assign valid_29_23 = io_inValid_23 & _T_10424; // @[Switch.scala 30:36:@4778.4]
  assign _T_10427 = io_inAddr_24 == 5'h1d; // @[Switch.scala 30:53:@4780.4]
  assign valid_29_24 = io_inValid_24 & _T_10427; // @[Switch.scala 30:36:@4781.4]
  assign _T_10430 = io_inAddr_25 == 5'h1d; // @[Switch.scala 30:53:@4783.4]
  assign valid_29_25 = io_inValid_25 & _T_10430; // @[Switch.scala 30:36:@4784.4]
  assign _T_10433 = io_inAddr_26 == 5'h1d; // @[Switch.scala 30:53:@4786.4]
  assign valid_29_26 = io_inValid_26 & _T_10433; // @[Switch.scala 30:36:@4787.4]
  assign _T_10436 = io_inAddr_27 == 5'h1d; // @[Switch.scala 30:53:@4789.4]
  assign valid_29_27 = io_inValid_27 & _T_10436; // @[Switch.scala 30:36:@4790.4]
  assign _T_10439 = io_inAddr_28 == 5'h1d; // @[Switch.scala 30:53:@4792.4]
  assign valid_29_28 = io_inValid_28 & _T_10439; // @[Switch.scala 30:36:@4793.4]
  assign _T_10442 = io_inAddr_29 == 5'h1d; // @[Switch.scala 30:53:@4795.4]
  assign valid_29_29 = io_inValid_29 & _T_10442; // @[Switch.scala 30:36:@4796.4]
  assign _T_10445 = io_inAddr_30 == 5'h1d; // @[Switch.scala 30:53:@4798.4]
  assign valid_29_30 = io_inValid_30 & _T_10445; // @[Switch.scala 30:36:@4799.4]
  assign _T_10448 = io_inAddr_31 == 5'h1d; // @[Switch.scala 30:53:@4801.4]
  assign valid_29_31 = io_inValid_31 & _T_10448; // @[Switch.scala 30:36:@4802.4]
  assign _T_10482 = valid_29_30 ? 5'h1e : 5'h1f; // @[Mux.scala 31:69:@4804.4]
  assign _T_10483 = valid_29_29 ? 5'h1d : _T_10482; // @[Mux.scala 31:69:@4805.4]
  assign _T_10484 = valid_29_28 ? 5'h1c : _T_10483; // @[Mux.scala 31:69:@4806.4]
  assign _T_10485 = valid_29_27 ? 5'h1b : _T_10484; // @[Mux.scala 31:69:@4807.4]
  assign _T_10486 = valid_29_26 ? 5'h1a : _T_10485; // @[Mux.scala 31:69:@4808.4]
  assign _T_10487 = valid_29_25 ? 5'h19 : _T_10486; // @[Mux.scala 31:69:@4809.4]
  assign _T_10488 = valid_29_24 ? 5'h18 : _T_10487; // @[Mux.scala 31:69:@4810.4]
  assign _T_10489 = valid_29_23 ? 5'h17 : _T_10488; // @[Mux.scala 31:69:@4811.4]
  assign _T_10490 = valid_29_22 ? 5'h16 : _T_10489; // @[Mux.scala 31:69:@4812.4]
  assign _T_10491 = valid_29_21 ? 5'h15 : _T_10490; // @[Mux.scala 31:69:@4813.4]
  assign _T_10492 = valid_29_20 ? 5'h14 : _T_10491; // @[Mux.scala 31:69:@4814.4]
  assign _T_10493 = valid_29_19 ? 5'h13 : _T_10492; // @[Mux.scala 31:69:@4815.4]
  assign _T_10494 = valid_29_18 ? 5'h12 : _T_10493; // @[Mux.scala 31:69:@4816.4]
  assign _T_10495 = valid_29_17 ? 5'h11 : _T_10494; // @[Mux.scala 31:69:@4817.4]
  assign _T_10496 = valid_29_16 ? 5'h10 : _T_10495; // @[Mux.scala 31:69:@4818.4]
  assign _T_10497 = valid_29_15 ? 5'hf : _T_10496; // @[Mux.scala 31:69:@4819.4]
  assign _T_10498 = valid_29_14 ? 5'he : _T_10497; // @[Mux.scala 31:69:@4820.4]
  assign _T_10499 = valid_29_13 ? 5'hd : _T_10498; // @[Mux.scala 31:69:@4821.4]
  assign _T_10500 = valid_29_12 ? 5'hc : _T_10499; // @[Mux.scala 31:69:@4822.4]
  assign _T_10501 = valid_29_11 ? 5'hb : _T_10500; // @[Mux.scala 31:69:@4823.4]
  assign _T_10502 = valid_29_10 ? 5'ha : _T_10501; // @[Mux.scala 31:69:@4824.4]
  assign _T_10503 = valid_29_9 ? 5'h9 : _T_10502; // @[Mux.scala 31:69:@4825.4]
  assign _T_10504 = valid_29_8 ? 5'h8 : _T_10503; // @[Mux.scala 31:69:@4826.4]
  assign _T_10505 = valid_29_7 ? 5'h7 : _T_10504; // @[Mux.scala 31:69:@4827.4]
  assign _T_10506 = valid_29_6 ? 5'h6 : _T_10505; // @[Mux.scala 31:69:@4828.4]
  assign _T_10507 = valid_29_5 ? 5'h5 : _T_10506; // @[Mux.scala 31:69:@4829.4]
  assign _T_10508 = valid_29_4 ? 5'h4 : _T_10507; // @[Mux.scala 31:69:@4830.4]
  assign _T_10509 = valid_29_3 ? 5'h3 : _T_10508; // @[Mux.scala 31:69:@4831.4]
  assign _T_10510 = valid_29_2 ? 5'h2 : _T_10509; // @[Mux.scala 31:69:@4832.4]
  assign _T_10511 = valid_29_1 ? 5'h1 : _T_10510; // @[Mux.scala 31:69:@4833.4]
  assign select_29 = valid_29_0 ? 5'h0 : _T_10511; // @[Mux.scala 31:69:@4834.4]
  assign _GEN_929 = 5'h1 == select_29 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@4836.4]
  assign _GEN_930 = 5'h2 == select_29 ? io_inData_2 : _GEN_929; // @[Switch.scala 33:19:@4836.4]
  assign _GEN_931 = 5'h3 == select_29 ? io_inData_3 : _GEN_930; // @[Switch.scala 33:19:@4836.4]
  assign _GEN_932 = 5'h4 == select_29 ? io_inData_4 : _GEN_931; // @[Switch.scala 33:19:@4836.4]
  assign _GEN_933 = 5'h5 == select_29 ? io_inData_5 : _GEN_932; // @[Switch.scala 33:19:@4836.4]
  assign _GEN_934 = 5'h6 == select_29 ? io_inData_6 : _GEN_933; // @[Switch.scala 33:19:@4836.4]
  assign _GEN_935 = 5'h7 == select_29 ? io_inData_7 : _GEN_934; // @[Switch.scala 33:19:@4836.4]
  assign _GEN_936 = 5'h8 == select_29 ? io_inData_8 : _GEN_935; // @[Switch.scala 33:19:@4836.4]
  assign _GEN_937 = 5'h9 == select_29 ? io_inData_9 : _GEN_936; // @[Switch.scala 33:19:@4836.4]
  assign _GEN_938 = 5'ha == select_29 ? io_inData_10 : _GEN_937; // @[Switch.scala 33:19:@4836.4]
  assign _GEN_939 = 5'hb == select_29 ? io_inData_11 : _GEN_938; // @[Switch.scala 33:19:@4836.4]
  assign _GEN_940 = 5'hc == select_29 ? io_inData_12 : _GEN_939; // @[Switch.scala 33:19:@4836.4]
  assign _GEN_941 = 5'hd == select_29 ? io_inData_13 : _GEN_940; // @[Switch.scala 33:19:@4836.4]
  assign _GEN_942 = 5'he == select_29 ? io_inData_14 : _GEN_941; // @[Switch.scala 33:19:@4836.4]
  assign _GEN_943 = 5'hf == select_29 ? io_inData_15 : _GEN_942; // @[Switch.scala 33:19:@4836.4]
  assign _GEN_944 = 5'h10 == select_29 ? io_inData_16 : _GEN_943; // @[Switch.scala 33:19:@4836.4]
  assign _GEN_945 = 5'h11 == select_29 ? io_inData_17 : _GEN_944; // @[Switch.scala 33:19:@4836.4]
  assign _GEN_946 = 5'h12 == select_29 ? io_inData_18 : _GEN_945; // @[Switch.scala 33:19:@4836.4]
  assign _GEN_947 = 5'h13 == select_29 ? io_inData_19 : _GEN_946; // @[Switch.scala 33:19:@4836.4]
  assign _GEN_948 = 5'h14 == select_29 ? io_inData_20 : _GEN_947; // @[Switch.scala 33:19:@4836.4]
  assign _GEN_949 = 5'h15 == select_29 ? io_inData_21 : _GEN_948; // @[Switch.scala 33:19:@4836.4]
  assign _GEN_950 = 5'h16 == select_29 ? io_inData_22 : _GEN_949; // @[Switch.scala 33:19:@4836.4]
  assign _GEN_951 = 5'h17 == select_29 ? io_inData_23 : _GEN_950; // @[Switch.scala 33:19:@4836.4]
  assign _GEN_952 = 5'h18 == select_29 ? io_inData_24 : _GEN_951; // @[Switch.scala 33:19:@4836.4]
  assign _GEN_953 = 5'h19 == select_29 ? io_inData_25 : _GEN_952; // @[Switch.scala 33:19:@4836.4]
  assign _GEN_954 = 5'h1a == select_29 ? io_inData_26 : _GEN_953; // @[Switch.scala 33:19:@4836.4]
  assign _GEN_955 = 5'h1b == select_29 ? io_inData_27 : _GEN_954; // @[Switch.scala 33:19:@4836.4]
  assign _GEN_956 = 5'h1c == select_29 ? io_inData_28 : _GEN_955; // @[Switch.scala 33:19:@4836.4]
  assign _GEN_957 = 5'h1d == select_29 ? io_inData_29 : _GEN_956; // @[Switch.scala 33:19:@4836.4]
  assign _GEN_958 = 5'h1e == select_29 ? io_inData_30 : _GEN_957; // @[Switch.scala 33:19:@4836.4]
  assign _T_10520 = {valid_29_7,valid_29_6,valid_29_5,valid_29_4,valid_29_3,valid_29_2,valid_29_1,valid_29_0}; // @[Switch.scala 34:32:@4843.4]
  assign _T_10528 = {valid_29_15,valid_29_14,valid_29_13,valid_29_12,valid_29_11,valid_29_10,valid_29_9,valid_29_8,_T_10520}; // @[Switch.scala 34:32:@4851.4]
  assign _T_10535 = {valid_29_23,valid_29_22,valid_29_21,valid_29_20,valid_29_19,valid_29_18,valid_29_17,valid_29_16}; // @[Switch.scala 34:32:@4858.4]
  assign _T_10544 = {valid_29_31,valid_29_30,valid_29_29,valid_29_28,valid_29_27,valid_29_26,valid_29_25,valid_29_24,_T_10535,_T_10528}; // @[Switch.scala 34:32:@4867.4]
  assign _T_10548 = io_inAddr_0 == 5'h1e; // @[Switch.scala 30:53:@4870.4]
  assign valid_30_0 = io_inValid_0 & _T_10548; // @[Switch.scala 30:36:@4871.4]
  assign _T_10551 = io_inAddr_1 == 5'h1e; // @[Switch.scala 30:53:@4873.4]
  assign valid_30_1 = io_inValid_1 & _T_10551; // @[Switch.scala 30:36:@4874.4]
  assign _T_10554 = io_inAddr_2 == 5'h1e; // @[Switch.scala 30:53:@4876.4]
  assign valid_30_2 = io_inValid_2 & _T_10554; // @[Switch.scala 30:36:@4877.4]
  assign _T_10557 = io_inAddr_3 == 5'h1e; // @[Switch.scala 30:53:@4879.4]
  assign valid_30_3 = io_inValid_3 & _T_10557; // @[Switch.scala 30:36:@4880.4]
  assign _T_10560 = io_inAddr_4 == 5'h1e; // @[Switch.scala 30:53:@4882.4]
  assign valid_30_4 = io_inValid_4 & _T_10560; // @[Switch.scala 30:36:@4883.4]
  assign _T_10563 = io_inAddr_5 == 5'h1e; // @[Switch.scala 30:53:@4885.4]
  assign valid_30_5 = io_inValid_5 & _T_10563; // @[Switch.scala 30:36:@4886.4]
  assign _T_10566 = io_inAddr_6 == 5'h1e; // @[Switch.scala 30:53:@4888.4]
  assign valid_30_6 = io_inValid_6 & _T_10566; // @[Switch.scala 30:36:@4889.4]
  assign _T_10569 = io_inAddr_7 == 5'h1e; // @[Switch.scala 30:53:@4891.4]
  assign valid_30_7 = io_inValid_7 & _T_10569; // @[Switch.scala 30:36:@4892.4]
  assign _T_10572 = io_inAddr_8 == 5'h1e; // @[Switch.scala 30:53:@4894.4]
  assign valid_30_8 = io_inValid_8 & _T_10572; // @[Switch.scala 30:36:@4895.4]
  assign _T_10575 = io_inAddr_9 == 5'h1e; // @[Switch.scala 30:53:@4897.4]
  assign valid_30_9 = io_inValid_9 & _T_10575; // @[Switch.scala 30:36:@4898.4]
  assign _T_10578 = io_inAddr_10 == 5'h1e; // @[Switch.scala 30:53:@4900.4]
  assign valid_30_10 = io_inValid_10 & _T_10578; // @[Switch.scala 30:36:@4901.4]
  assign _T_10581 = io_inAddr_11 == 5'h1e; // @[Switch.scala 30:53:@4903.4]
  assign valid_30_11 = io_inValid_11 & _T_10581; // @[Switch.scala 30:36:@4904.4]
  assign _T_10584 = io_inAddr_12 == 5'h1e; // @[Switch.scala 30:53:@4906.4]
  assign valid_30_12 = io_inValid_12 & _T_10584; // @[Switch.scala 30:36:@4907.4]
  assign _T_10587 = io_inAddr_13 == 5'h1e; // @[Switch.scala 30:53:@4909.4]
  assign valid_30_13 = io_inValid_13 & _T_10587; // @[Switch.scala 30:36:@4910.4]
  assign _T_10590 = io_inAddr_14 == 5'h1e; // @[Switch.scala 30:53:@4912.4]
  assign valid_30_14 = io_inValid_14 & _T_10590; // @[Switch.scala 30:36:@4913.4]
  assign _T_10593 = io_inAddr_15 == 5'h1e; // @[Switch.scala 30:53:@4915.4]
  assign valid_30_15 = io_inValid_15 & _T_10593; // @[Switch.scala 30:36:@4916.4]
  assign _T_10596 = io_inAddr_16 == 5'h1e; // @[Switch.scala 30:53:@4918.4]
  assign valid_30_16 = io_inValid_16 & _T_10596; // @[Switch.scala 30:36:@4919.4]
  assign _T_10599 = io_inAddr_17 == 5'h1e; // @[Switch.scala 30:53:@4921.4]
  assign valid_30_17 = io_inValid_17 & _T_10599; // @[Switch.scala 30:36:@4922.4]
  assign _T_10602 = io_inAddr_18 == 5'h1e; // @[Switch.scala 30:53:@4924.4]
  assign valid_30_18 = io_inValid_18 & _T_10602; // @[Switch.scala 30:36:@4925.4]
  assign _T_10605 = io_inAddr_19 == 5'h1e; // @[Switch.scala 30:53:@4927.4]
  assign valid_30_19 = io_inValid_19 & _T_10605; // @[Switch.scala 30:36:@4928.4]
  assign _T_10608 = io_inAddr_20 == 5'h1e; // @[Switch.scala 30:53:@4930.4]
  assign valid_30_20 = io_inValid_20 & _T_10608; // @[Switch.scala 30:36:@4931.4]
  assign _T_10611 = io_inAddr_21 == 5'h1e; // @[Switch.scala 30:53:@4933.4]
  assign valid_30_21 = io_inValid_21 & _T_10611; // @[Switch.scala 30:36:@4934.4]
  assign _T_10614 = io_inAddr_22 == 5'h1e; // @[Switch.scala 30:53:@4936.4]
  assign valid_30_22 = io_inValid_22 & _T_10614; // @[Switch.scala 30:36:@4937.4]
  assign _T_10617 = io_inAddr_23 == 5'h1e; // @[Switch.scala 30:53:@4939.4]
  assign valid_30_23 = io_inValid_23 & _T_10617; // @[Switch.scala 30:36:@4940.4]
  assign _T_10620 = io_inAddr_24 == 5'h1e; // @[Switch.scala 30:53:@4942.4]
  assign valid_30_24 = io_inValid_24 & _T_10620; // @[Switch.scala 30:36:@4943.4]
  assign _T_10623 = io_inAddr_25 == 5'h1e; // @[Switch.scala 30:53:@4945.4]
  assign valid_30_25 = io_inValid_25 & _T_10623; // @[Switch.scala 30:36:@4946.4]
  assign _T_10626 = io_inAddr_26 == 5'h1e; // @[Switch.scala 30:53:@4948.4]
  assign valid_30_26 = io_inValid_26 & _T_10626; // @[Switch.scala 30:36:@4949.4]
  assign _T_10629 = io_inAddr_27 == 5'h1e; // @[Switch.scala 30:53:@4951.4]
  assign valid_30_27 = io_inValid_27 & _T_10629; // @[Switch.scala 30:36:@4952.4]
  assign _T_10632 = io_inAddr_28 == 5'h1e; // @[Switch.scala 30:53:@4954.4]
  assign valid_30_28 = io_inValid_28 & _T_10632; // @[Switch.scala 30:36:@4955.4]
  assign _T_10635 = io_inAddr_29 == 5'h1e; // @[Switch.scala 30:53:@4957.4]
  assign valid_30_29 = io_inValid_29 & _T_10635; // @[Switch.scala 30:36:@4958.4]
  assign _T_10638 = io_inAddr_30 == 5'h1e; // @[Switch.scala 30:53:@4960.4]
  assign valid_30_30 = io_inValid_30 & _T_10638; // @[Switch.scala 30:36:@4961.4]
  assign _T_10641 = io_inAddr_31 == 5'h1e; // @[Switch.scala 30:53:@4963.4]
  assign valid_30_31 = io_inValid_31 & _T_10641; // @[Switch.scala 30:36:@4964.4]
  assign _T_10675 = valid_30_30 ? 5'h1e : 5'h1f; // @[Mux.scala 31:69:@4966.4]
  assign _T_10676 = valid_30_29 ? 5'h1d : _T_10675; // @[Mux.scala 31:69:@4967.4]
  assign _T_10677 = valid_30_28 ? 5'h1c : _T_10676; // @[Mux.scala 31:69:@4968.4]
  assign _T_10678 = valid_30_27 ? 5'h1b : _T_10677; // @[Mux.scala 31:69:@4969.4]
  assign _T_10679 = valid_30_26 ? 5'h1a : _T_10678; // @[Mux.scala 31:69:@4970.4]
  assign _T_10680 = valid_30_25 ? 5'h19 : _T_10679; // @[Mux.scala 31:69:@4971.4]
  assign _T_10681 = valid_30_24 ? 5'h18 : _T_10680; // @[Mux.scala 31:69:@4972.4]
  assign _T_10682 = valid_30_23 ? 5'h17 : _T_10681; // @[Mux.scala 31:69:@4973.4]
  assign _T_10683 = valid_30_22 ? 5'h16 : _T_10682; // @[Mux.scala 31:69:@4974.4]
  assign _T_10684 = valid_30_21 ? 5'h15 : _T_10683; // @[Mux.scala 31:69:@4975.4]
  assign _T_10685 = valid_30_20 ? 5'h14 : _T_10684; // @[Mux.scala 31:69:@4976.4]
  assign _T_10686 = valid_30_19 ? 5'h13 : _T_10685; // @[Mux.scala 31:69:@4977.4]
  assign _T_10687 = valid_30_18 ? 5'h12 : _T_10686; // @[Mux.scala 31:69:@4978.4]
  assign _T_10688 = valid_30_17 ? 5'h11 : _T_10687; // @[Mux.scala 31:69:@4979.4]
  assign _T_10689 = valid_30_16 ? 5'h10 : _T_10688; // @[Mux.scala 31:69:@4980.4]
  assign _T_10690 = valid_30_15 ? 5'hf : _T_10689; // @[Mux.scala 31:69:@4981.4]
  assign _T_10691 = valid_30_14 ? 5'he : _T_10690; // @[Mux.scala 31:69:@4982.4]
  assign _T_10692 = valid_30_13 ? 5'hd : _T_10691; // @[Mux.scala 31:69:@4983.4]
  assign _T_10693 = valid_30_12 ? 5'hc : _T_10692; // @[Mux.scala 31:69:@4984.4]
  assign _T_10694 = valid_30_11 ? 5'hb : _T_10693; // @[Mux.scala 31:69:@4985.4]
  assign _T_10695 = valid_30_10 ? 5'ha : _T_10694; // @[Mux.scala 31:69:@4986.4]
  assign _T_10696 = valid_30_9 ? 5'h9 : _T_10695; // @[Mux.scala 31:69:@4987.4]
  assign _T_10697 = valid_30_8 ? 5'h8 : _T_10696; // @[Mux.scala 31:69:@4988.4]
  assign _T_10698 = valid_30_7 ? 5'h7 : _T_10697; // @[Mux.scala 31:69:@4989.4]
  assign _T_10699 = valid_30_6 ? 5'h6 : _T_10698; // @[Mux.scala 31:69:@4990.4]
  assign _T_10700 = valid_30_5 ? 5'h5 : _T_10699; // @[Mux.scala 31:69:@4991.4]
  assign _T_10701 = valid_30_4 ? 5'h4 : _T_10700; // @[Mux.scala 31:69:@4992.4]
  assign _T_10702 = valid_30_3 ? 5'h3 : _T_10701; // @[Mux.scala 31:69:@4993.4]
  assign _T_10703 = valid_30_2 ? 5'h2 : _T_10702; // @[Mux.scala 31:69:@4994.4]
  assign _T_10704 = valid_30_1 ? 5'h1 : _T_10703; // @[Mux.scala 31:69:@4995.4]
  assign select_30 = valid_30_0 ? 5'h0 : _T_10704; // @[Mux.scala 31:69:@4996.4]
  assign _GEN_961 = 5'h1 == select_30 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@4998.4]
  assign _GEN_962 = 5'h2 == select_30 ? io_inData_2 : _GEN_961; // @[Switch.scala 33:19:@4998.4]
  assign _GEN_963 = 5'h3 == select_30 ? io_inData_3 : _GEN_962; // @[Switch.scala 33:19:@4998.4]
  assign _GEN_964 = 5'h4 == select_30 ? io_inData_4 : _GEN_963; // @[Switch.scala 33:19:@4998.4]
  assign _GEN_965 = 5'h5 == select_30 ? io_inData_5 : _GEN_964; // @[Switch.scala 33:19:@4998.4]
  assign _GEN_966 = 5'h6 == select_30 ? io_inData_6 : _GEN_965; // @[Switch.scala 33:19:@4998.4]
  assign _GEN_967 = 5'h7 == select_30 ? io_inData_7 : _GEN_966; // @[Switch.scala 33:19:@4998.4]
  assign _GEN_968 = 5'h8 == select_30 ? io_inData_8 : _GEN_967; // @[Switch.scala 33:19:@4998.4]
  assign _GEN_969 = 5'h9 == select_30 ? io_inData_9 : _GEN_968; // @[Switch.scala 33:19:@4998.4]
  assign _GEN_970 = 5'ha == select_30 ? io_inData_10 : _GEN_969; // @[Switch.scala 33:19:@4998.4]
  assign _GEN_971 = 5'hb == select_30 ? io_inData_11 : _GEN_970; // @[Switch.scala 33:19:@4998.4]
  assign _GEN_972 = 5'hc == select_30 ? io_inData_12 : _GEN_971; // @[Switch.scala 33:19:@4998.4]
  assign _GEN_973 = 5'hd == select_30 ? io_inData_13 : _GEN_972; // @[Switch.scala 33:19:@4998.4]
  assign _GEN_974 = 5'he == select_30 ? io_inData_14 : _GEN_973; // @[Switch.scala 33:19:@4998.4]
  assign _GEN_975 = 5'hf == select_30 ? io_inData_15 : _GEN_974; // @[Switch.scala 33:19:@4998.4]
  assign _GEN_976 = 5'h10 == select_30 ? io_inData_16 : _GEN_975; // @[Switch.scala 33:19:@4998.4]
  assign _GEN_977 = 5'h11 == select_30 ? io_inData_17 : _GEN_976; // @[Switch.scala 33:19:@4998.4]
  assign _GEN_978 = 5'h12 == select_30 ? io_inData_18 : _GEN_977; // @[Switch.scala 33:19:@4998.4]
  assign _GEN_979 = 5'h13 == select_30 ? io_inData_19 : _GEN_978; // @[Switch.scala 33:19:@4998.4]
  assign _GEN_980 = 5'h14 == select_30 ? io_inData_20 : _GEN_979; // @[Switch.scala 33:19:@4998.4]
  assign _GEN_981 = 5'h15 == select_30 ? io_inData_21 : _GEN_980; // @[Switch.scala 33:19:@4998.4]
  assign _GEN_982 = 5'h16 == select_30 ? io_inData_22 : _GEN_981; // @[Switch.scala 33:19:@4998.4]
  assign _GEN_983 = 5'h17 == select_30 ? io_inData_23 : _GEN_982; // @[Switch.scala 33:19:@4998.4]
  assign _GEN_984 = 5'h18 == select_30 ? io_inData_24 : _GEN_983; // @[Switch.scala 33:19:@4998.4]
  assign _GEN_985 = 5'h19 == select_30 ? io_inData_25 : _GEN_984; // @[Switch.scala 33:19:@4998.4]
  assign _GEN_986 = 5'h1a == select_30 ? io_inData_26 : _GEN_985; // @[Switch.scala 33:19:@4998.4]
  assign _GEN_987 = 5'h1b == select_30 ? io_inData_27 : _GEN_986; // @[Switch.scala 33:19:@4998.4]
  assign _GEN_988 = 5'h1c == select_30 ? io_inData_28 : _GEN_987; // @[Switch.scala 33:19:@4998.4]
  assign _GEN_989 = 5'h1d == select_30 ? io_inData_29 : _GEN_988; // @[Switch.scala 33:19:@4998.4]
  assign _GEN_990 = 5'h1e == select_30 ? io_inData_30 : _GEN_989; // @[Switch.scala 33:19:@4998.4]
  assign _T_10713 = {valid_30_7,valid_30_6,valid_30_5,valid_30_4,valid_30_3,valid_30_2,valid_30_1,valid_30_0}; // @[Switch.scala 34:32:@5005.4]
  assign _T_10721 = {valid_30_15,valid_30_14,valid_30_13,valid_30_12,valid_30_11,valid_30_10,valid_30_9,valid_30_8,_T_10713}; // @[Switch.scala 34:32:@5013.4]
  assign _T_10728 = {valid_30_23,valid_30_22,valid_30_21,valid_30_20,valid_30_19,valid_30_18,valid_30_17,valid_30_16}; // @[Switch.scala 34:32:@5020.4]
  assign _T_10737 = {valid_30_31,valid_30_30,valid_30_29,valid_30_28,valid_30_27,valid_30_26,valid_30_25,valid_30_24,_T_10728,_T_10721}; // @[Switch.scala 34:32:@5029.4]
  assign _T_10741 = io_inAddr_0 == 5'h1f; // @[Switch.scala 30:53:@5032.4]
  assign valid_31_0 = io_inValid_0 & _T_10741; // @[Switch.scala 30:36:@5033.4]
  assign _T_10744 = io_inAddr_1 == 5'h1f; // @[Switch.scala 30:53:@5035.4]
  assign valid_31_1 = io_inValid_1 & _T_10744; // @[Switch.scala 30:36:@5036.4]
  assign _T_10747 = io_inAddr_2 == 5'h1f; // @[Switch.scala 30:53:@5038.4]
  assign valid_31_2 = io_inValid_2 & _T_10747; // @[Switch.scala 30:36:@5039.4]
  assign _T_10750 = io_inAddr_3 == 5'h1f; // @[Switch.scala 30:53:@5041.4]
  assign valid_31_3 = io_inValid_3 & _T_10750; // @[Switch.scala 30:36:@5042.4]
  assign _T_10753 = io_inAddr_4 == 5'h1f; // @[Switch.scala 30:53:@5044.4]
  assign valid_31_4 = io_inValid_4 & _T_10753; // @[Switch.scala 30:36:@5045.4]
  assign _T_10756 = io_inAddr_5 == 5'h1f; // @[Switch.scala 30:53:@5047.4]
  assign valid_31_5 = io_inValid_5 & _T_10756; // @[Switch.scala 30:36:@5048.4]
  assign _T_10759 = io_inAddr_6 == 5'h1f; // @[Switch.scala 30:53:@5050.4]
  assign valid_31_6 = io_inValid_6 & _T_10759; // @[Switch.scala 30:36:@5051.4]
  assign _T_10762 = io_inAddr_7 == 5'h1f; // @[Switch.scala 30:53:@5053.4]
  assign valid_31_7 = io_inValid_7 & _T_10762; // @[Switch.scala 30:36:@5054.4]
  assign _T_10765 = io_inAddr_8 == 5'h1f; // @[Switch.scala 30:53:@5056.4]
  assign valid_31_8 = io_inValid_8 & _T_10765; // @[Switch.scala 30:36:@5057.4]
  assign _T_10768 = io_inAddr_9 == 5'h1f; // @[Switch.scala 30:53:@5059.4]
  assign valid_31_9 = io_inValid_9 & _T_10768; // @[Switch.scala 30:36:@5060.4]
  assign _T_10771 = io_inAddr_10 == 5'h1f; // @[Switch.scala 30:53:@5062.4]
  assign valid_31_10 = io_inValid_10 & _T_10771; // @[Switch.scala 30:36:@5063.4]
  assign _T_10774 = io_inAddr_11 == 5'h1f; // @[Switch.scala 30:53:@5065.4]
  assign valid_31_11 = io_inValid_11 & _T_10774; // @[Switch.scala 30:36:@5066.4]
  assign _T_10777 = io_inAddr_12 == 5'h1f; // @[Switch.scala 30:53:@5068.4]
  assign valid_31_12 = io_inValid_12 & _T_10777; // @[Switch.scala 30:36:@5069.4]
  assign _T_10780 = io_inAddr_13 == 5'h1f; // @[Switch.scala 30:53:@5071.4]
  assign valid_31_13 = io_inValid_13 & _T_10780; // @[Switch.scala 30:36:@5072.4]
  assign _T_10783 = io_inAddr_14 == 5'h1f; // @[Switch.scala 30:53:@5074.4]
  assign valid_31_14 = io_inValid_14 & _T_10783; // @[Switch.scala 30:36:@5075.4]
  assign _T_10786 = io_inAddr_15 == 5'h1f; // @[Switch.scala 30:53:@5077.4]
  assign valid_31_15 = io_inValid_15 & _T_10786; // @[Switch.scala 30:36:@5078.4]
  assign _T_10789 = io_inAddr_16 == 5'h1f; // @[Switch.scala 30:53:@5080.4]
  assign valid_31_16 = io_inValid_16 & _T_10789; // @[Switch.scala 30:36:@5081.4]
  assign _T_10792 = io_inAddr_17 == 5'h1f; // @[Switch.scala 30:53:@5083.4]
  assign valid_31_17 = io_inValid_17 & _T_10792; // @[Switch.scala 30:36:@5084.4]
  assign _T_10795 = io_inAddr_18 == 5'h1f; // @[Switch.scala 30:53:@5086.4]
  assign valid_31_18 = io_inValid_18 & _T_10795; // @[Switch.scala 30:36:@5087.4]
  assign _T_10798 = io_inAddr_19 == 5'h1f; // @[Switch.scala 30:53:@5089.4]
  assign valid_31_19 = io_inValid_19 & _T_10798; // @[Switch.scala 30:36:@5090.4]
  assign _T_10801 = io_inAddr_20 == 5'h1f; // @[Switch.scala 30:53:@5092.4]
  assign valid_31_20 = io_inValid_20 & _T_10801; // @[Switch.scala 30:36:@5093.4]
  assign _T_10804 = io_inAddr_21 == 5'h1f; // @[Switch.scala 30:53:@5095.4]
  assign valid_31_21 = io_inValid_21 & _T_10804; // @[Switch.scala 30:36:@5096.4]
  assign _T_10807 = io_inAddr_22 == 5'h1f; // @[Switch.scala 30:53:@5098.4]
  assign valid_31_22 = io_inValid_22 & _T_10807; // @[Switch.scala 30:36:@5099.4]
  assign _T_10810 = io_inAddr_23 == 5'h1f; // @[Switch.scala 30:53:@5101.4]
  assign valid_31_23 = io_inValid_23 & _T_10810; // @[Switch.scala 30:36:@5102.4]
  assign _T_10813 = io_inAddr_24 == 5'h1f; // @[Switch.scala 30:53:@5104.4]
  assign valid_31_24 = io_inValid_24 & _T_10813; // @[Switch.scala 30:36:@5105.4]
  assign _T_10816 = io_inAddr_25 == 5'h1f; // @[Switch.scala 30:53:@5107.4]
  assign valid_31_25 = io_inValid_25 & _T_10816; // @[Switch.scala 30:36:@5108.4]
  assign _T_10819 = io_inAddr_26 == 5'h1f; // @[Switch.scala 30:53:@5110.4]
  assign valid_31_26 = io_inValid_26 & _T_10819; // @[Switch.scala 30:36:@5111.4]
  assign _T_10822 = io_inAddr_27 == 5'h1f; // @[Switch.scala 30:53:@5113.4]
  assign valid_31_27 = io_inValid_27 & _T_10822; // @[Switch.scala 30:36:@5114.4]
  assign _T_10825 = io_inAddr_28 == 5'h1f; // @[Switch.scala 30:53:@5116.4]
  assign valid_31_28 = io_inValid_28 & _T_10825; // @[Switch.scala 30:36:@5117.4]
  assign _T_10828 = io_inAddr_29 == 5'h1f; // @[Switch.scala 30:53:@5119.4]
  assign valid_31_29 = io_inValid_29 & _T_10828; // @[Switch.scala 30:36:@5120.4]
  assign _T_10831 = io_inAddr_30 == 5'h1f; // @[Switch.scala 30:53:@5122.4]
  assign valid_31_30 = io_inValid_30 & _T_10831; // @[Switch.scala 30:36:@5123.4]
  assign _T_10834 = io_inAddr_31 == 5'h1f; // @[Switch.scala 30:53:@5125.4]
  assign valid_31_31 = io_inValid_31 & _T_10834; // @[Switch.scala 30:36:@5126.4]
  assign _T_10868 = valid_31_30 ? 5'h1e : 5'h1f; // @[Mux.scala 31:69:@5128.4]
  assign _T_10869 = valid_31_29 ? 5'h1d : _T_10868; // @[Mux.scala 31:69:@5129.4]
  assign _T_10870 = valid_31_28 ? 5'h1c : _T_10869; // @[Mux.scala 31:69:@5130.4]
  assign _T_10871 = valid_31_27 ? 5'h1b : _T_10870; // @[Mux.scala 31:69:@5131.4]
  assign _T_10872 = valid_31_26 ? 5'h1a : _T_10871; // @[Mux.scala 31:69:@5132.4]
  assign _T_10873 = valid_31_25 ? 5'h19 : _T_10872; // @[Mux.scala 31:69:@5133.4]
  assign _T_10874 = valid_31_24 ? 5'h18 : _T_10873; // @[Mux.scala 31:69:@5134.4]
  assign _T_10875 = valid_31_23 ? 5'h17 : _T_10874; // @[Mux.scala 31:69:@5135.4]
  assign _T_10876 = valid_31_22 ? 5'h16 : _T_10875; // @[Mux.scala 31:69:@5136.4]
  assign _T_10877 = valid_31_21 ? 5'h15 : _T_10876; // @[Mux.scala 31:69:@5137.4]
  assign _T_10878 = valid_31_20 ? 5'h14 : _T_10877; // @[Mux.scala 31:69:@5138.4]
  assign _T_10879 = valid_31_19 ? 5'h13 : _T_10878; // @[Mux.scala 31:69:@5139.4]
  assign _T_10880 = valid_31_18 ? 5'h12 : _T_10879; // @[Mux.scala 31:69:@5140.4]
  assign _T_10881 = valid_31_17 ? 5'h11 : _T_10880; // @[Mux.scala 31:69:@5141.4]
  assign _T_10882 = valid_31_16 ? 5'h10 : _T_10881; // @[Mux.scala 31:69:@5142.4]
  assign _T_10883 = valid_31_15 ? 5'hf : _T_10882; // @[Mux.scala 31:69:@5143.4]
  assign _T_10884 = valid_31_14 ? 5'he : _T_10883; // @[Mux.scala 31:69:@5144.4]
  assign _T_10885 = valid_31_13 ? 5'hd : _T_10884; // @[Mux.scala 31:69:@5145.4]
  assign _T_10886 = valid_31_12 ? 5'hc : _T_10885; // @[Mux.scala 31:69:@5146.4]
  assign _T_10887 = valid_31_11 ? 5'hb : _T_10886; // @[Mux.scala 31:69:@5147.4]
  assign _T_10888 = valid_31_10 ? 5'ha : _T_10887; // @[Mux.scala 31:69:@5148.4]
  assign _T_10889 = valid_31_9 ? 5'h9 : _T_10888; // @[Mux.scala 31:69:@5149.4]
  assign _T_10890 = valid_31_8 ? 5'h8 : _T_10889; // @[Mux.scala 31:69:@5150.4]
  assign _T_10891 = valid_31_7 ? 5'h7 : _T_10890; // @[Mux.scala 31:69:@5151.4]
  assign _T_10892 = valid_31_6 ? 5'h6 : _T_10891; // @[Mux.scala 31:69:@5152.4]
  assign _T_10893 = valid_31_5 ? 5'h5 : _T_10892; // @[Mux.scala 31:69:@5153.4]
  assign _T_10894 = valid_31_4 ? 5'h4 : _T_10893; // @[Mux.scala 31:69:@5154.4]
  assign _T_10895 = valid_31_3 ? 5'h3 : _T_10894; // @[Mux.scala 31:69:@5155.4]
  assign _T_10896 = valid_31_2 ? 5'h2 : _T_10895; // @[Mux.scala 31:69:@5156.4]
  assign _T_10897 = valid_31_1 ? 5'h1 : _T_10896; // @[Mux.scala 31:69:@5157.4]
  assign select_31 = valid_31_0 ? 5'h0 : _T_10897; // @[Mux.scala 31:69:@5158.4]
  assign _GEN_993 = 5'h1 == select_31 ? io_inData_1 : io_inData_0; // @[Switch.scala 33:19:@5160.4]
  assign _GEN_994 = 5'h2 == select_31 ? io_inData_2 : _GEN_993; // @[Switch.scala 33:19:@5160.4]
  assign _GEN_995 = 5'h3 == select_31 ? io_inData_3 : _GEN_994; // @[Switch.scala 33:19:@5160.4]
  assign _GEN_996 = 5'h4 == select_31 ? io_inData_4 : _GEN_995; // @[Switch.scala 33:19:@5160.4]
  assign _GEN_997 = 5'h5 == select_31 ? io_inData_5 : _GEN_996; // @[Switch.scala 33:19:@5160.4]
  assign _GEN_998 = 5'h6 == select_31 ? io_inData_6 : _GEN_997; // @[Switch.scala 33:19:@5160.4]
  assign _GEN_999 = 5'h7 == select_31 ? io_inData_7 : _GEN_998; // @[Switch.scala 33:19:@5160.4]
  assign _GEN_1000 = 5'h8 == select_31 ? io_inData_8 : _GEN_999; // @[Switch.scala 33:19:@5160.4]
  assign _GEN_1001 = 5'h9 == select_31 ? io_inData_9 : _GEN_1000; // @[Switch.scala 33:19:@5160.4]
  assign _GEN_1002 = 5'ha == select_31 ? io_inData_10 : _GEN_1001; // @[Switch.scala 33:19:@5160.4]
  assign _GEN_1003 = 5'hb == select_31 ? io_inData_11 : _GEN_1002; // @[Switch.scala 33:19:@5160.4]
  assign _GEN_1004 = 5'hc == select_31 ? io_inData_12 : _GEN_1003; // @[Switch.scala 33:19:@5160.4]
  assign _GEN_1005 = 5'hd == select_31 ? io_inData_13 : _GEN_1004; // @[Switch.scala 33:19:@5160.4]
  assign _GEN_1006 = 5'he == select_31 ? io_inData_14 : _GEN_1005; // @[Switch.scala 33:19:@5160.4]
  assign _GEN_1007 = 5'hf == select_31 ? io_inData_15 : _GEN_1006; // @[Switch.scala 33:19:@5160.4]
  assign _GEN_1008 = 5'h10 == select_31 ? io_inData_16 : _GEN_1007; // @[Switch.scala 33:19:@5160.4]
  assign _GEN_1009 = 5'h11 == select_31 ? io_inData_17 : _GEN_1008; // @[Switch.scala 33:19:@5160.4]
  assign _GEN_1010 = 5'h12 == select_31 ? io_inData_18 : _GEN_1009; // @[Switch.scala 33:19:@5160.4]
  assign _GEN_1011 = 5'h13 == select_31 ? io_inData_19 : _GEN_1010; // @[Switch.scala 33:19:@5160.4]
  assign _GEN_1012 = 5'h14 == select_31 ? io_inData_20 : _GEN_1011; // @[Switch.scala 33:19:@5160.4]
  assign _GEN_1013 = 5'h15 == select_31 ? io_inData_21 : _GEN_1012; // @[Switch.scala 33:19:@5160.4]
  assign _GEN_1014 = 5'h16 == select_31 ? io_inData_22 : _GEN_1013; // @[Switch.scala 33:19:@5160.4]
  assign _GEN_1015 = 5'h17 == select_31 ? io_inData_23 : _GEN_1014; // @[Switch.scala 33:19:@5160.4]
  assign _GEN_1016 = 5'h18 == select_31 ? io_inData_24 : _GEN_1015; // @[Switch.scala 33:19:@5160.4]
  assign _GEN_1017 = 5'h19 == select_31 ? io_inData_25 : _GEN_1016; // @[Switch.scala 33:19:@5160.4]
  assign _GEN_1018 = 5'h1a == select_31 ? io_inData_26 : _GEN_1017; // @[Switch.scala 33:19:@5160.4]
  assign _GEN_1019 = 5'h1b == select_31 ? io_inData_27 : _GEN_1018; // @[Switch.scala 33:19:@5160.4]
  assign _GEN_1020 = 5'h1c == select_31 ? io_inData_28 : _GEN_1019; // @[Switch.scala 33:19:@5160.4]
  assign _GEN_1021 = 5'h1d == select_31 ? io_inData_29 : _GEN_1020; // @[Switch.scala 33:19:@5160.4]
  assign _GEN_1022 = 5'h1e == select_31 ? io_inData_30 : _GEN_1021; // @[Switch.scala 33:19:@5160.4]
  assign _T_10906 = {valid_31_7,valid_31_6,valid_31_5,valid_31_4,valid_31_3,valid_31_2,valid_31_1,valid_31_0}; // @[Switch.scala 34:32:@5167.4]
  assign _T_10914 = {valid_31_15,valid_31_14,valid_31_13,valid_31_12,valid_31_11,valid_31_10,valid_31_9,valid_31_8,_T_10906}; // @[Switch.scala 34:32:@5175.4]
  assign _T_10921 = {valid_31_23,valid_31_22,valid_31_21,valid_31_20,valid_31_19,valid_31_18,valid_31_17,valid_31_16}; // @[Switch.scala 34:32:@5182.4]
  assign _T_10930 = {valid_31_31,valid_31_30,valid_31_29,valid_31_28,valid_31_27,valid_31_26,valid_31_25,valid_31_24,_T_10921,_T_10914}; // @[Switch.scala 34:32:@5191.4]
  assign _T_15428 = select_0 == 5'h0; // @[Switch.scala 41:52:@5195.4]
  assign output_0_0 = io_outValid_0 & _T_15428; // @[Switch.scala 41:38:@5196.4]
  assign _T_15431 = select_1 == 5'h0; // @[Switch.scala 41:52:@5198.4]
  assign output_0_1 = io_outValid_1 & _T_15431; // @[Switch.scala 41:38:@5199.4]
  assign _T_15434 = select_2 == 5'h0; // @[Switch.scala 41:52:@5201.4]
  assign output_0_2 = io_outValid_2 & _T_15434; // @[Switch.scala 41:38:@5202.4]
  assign _T_15437 = select_3 == 5'h0; // @[Switch.scala 41:52:@5204.4]
  assign output_0_3 = io_outValid_3 & _T_15437; // @[Switch.scala 41:38:@5205.4]
  assign _T_15440 = select_4 == 5'h0; // @[Switch.scala 41:52:@5207.4]
  assign output_0_4 = io_outValid_4 & _T_15440; // @[Switch.scala 41:38:@5208.4]
  assign _T_15443 = select_5 == 5'h0; // @[Switch.scala 41:52:@5210.4]
  assign output_0_5 = io_outValid_5 & _T_15443; // @[Switch.scala 41:38:@5211.4]
  assign _T_15446 = select_6 == 5'h0; // @[Switch.scala 41:52:@5213.4]
  assign output_0_6 = io_outValid_6 & _T_15446; // @[Switch.scala 41:38:@5214.4]
  assign _T_15449 = select_7 == 5'h0; // @[Switch.scala 41:52:@5216.4]
  assign output_0_7 = io_outValid_7 & _T_15449; // @[Switch.scala 41:38:@5217.4]
  assign _T_15452 = select_8 == 5'h0; // @[Switch.scala 41:52:@5219.4]
  assign output_0_8 = io_outValid_8 & _T_15452; // @[Switch.scala 41:38:@5220.4]
  assign _T_15455 = select_9 == 5'h0; // @[Switch.scala 41:52:@5222.4]
  assign output_0_9 = io_outValid_9 & _T_15455; // @[Switch.scala 41:38:@5223.4]
  assign _T_15458 = select_10 == 5'h0; // @[Switch.scala 41:52:@5225.4]
  assign output_0_10 = io_outValid_10 & _T_15458; // @[Switch.scala 41:38:@5226.4]
  assign _T_15461 = select_11 == 5'h0; // @[Switch.scala 41:52:@5228.4]
  assign output_0_11 = io_outValid_11 & _T_15461; // @[Switch.scala 41:38:@5229.4]
  assign _T_15464 = select_12 == 5'h0; // @[Switch.scala 41:52:@5231.4]
  assign output_0_12 = io_outValid_12 & _T_15464; // @[Switch.scala 41:38:@5232.4]
  assign _T_15467 = select_13 == 5'h0; // @[Switch.scala 41:52:@5234.4]
  assign output_0_13 = io_outValid_13 & _T_15467; // @[Switch.scala 41:38:@5235.4]
  assign _T_15470 = select_14 == 5'h0; // @[Switch.scala 41:52:@5237.4]
  assign output_0_14 = io_outValid_14 & _T_15470; // @[Switch.scala 41:38:@5238.4]
  assign _T_15473 = select_15 == 5'h0; // @[Switch.scala 41:52:@5240.4]
  assign output_0_15 = io_outValid_15 & _T_15473; // @[Switch.scala 41:38:@5241.4]
  assign _T_15476 = select_16 == 5'h0; // @[Switch.scala 41:52:@5243.4]
  assign output_0_16 = io_outValid_16 & _T_15476; // @[Switch.scala 41:38:@5244.4]
  assign _T_15479 = select_17 == 5'h0; // @[Switch.scala 41:52:@5246.4]
  assign output_0_17 = io_outValid_17 & _T_15479; // @[Switch.scala 41:38:@5247.4]
  assign _T_15482 = select_18 == 5'h0; // @[Switch.scala 41:52:@5249.4]
  assign output_0_18 = io_outValid_18 & _T_15482; // @[Switch.scala 41:38:@5250.4]
  assign _T_15485 = select_19 == 5'h0; // @[Switch.scala 41:52:@5252.4]
  assign output_0_19 = io_outValid_19 & _T_15485; // @[Switch.scala 41:38:@5253.4]
  assign _T_15488 = select_20 == 5'h0; // @[Switch.scala 41:52:@5255.4]
  assign output_0_20 = io_outValid_20 & _T_15488; // @[Switch.scala 41:38:@5256.4]
  assign _T_15491 = select_21 == 5'h0; // @[Switch.scala 41:52:@5258.4]
  assign output_0_21 = io_outValid_21 & _T_15491; // @[Switch.scala 41:38:@5259.4]
  assign _T_15494 = select_22 == 5'h0; // @[Switch.scala 41:52:@5261.4]
  assign output_0_22 = io_outValid_22 & _T_15494; // @[Switch.scala 41:38:@5262.4]
  assign _T_15497 = select_23 == 5'h0; // @[Switch.scala 41:52:@5264.4]
  assign output_0_23 = io_outValid_23 & _T_15497; // @[Switch.scala 41:38:@5265.4]
  assign _T_15500 = select_24 == 5'h0; // @[Switch.scala 41:52:@5267.4]
  assign output_0_24 = io_outValid_24 & _T_15500; // @[Switch.scala 41:38:@5268.4]
  assign _T_15503 = select_25 == 5'h0; // @[Switch.scala 41:52:@5270.4]
  assign output_0_25 = io_outValid_25 & _T_15503; // @[Switch.scala 41:38:@5271.4]
  assign _T_15506 = select_26 == 5'h0; // @[Switch.scala 41:52:@5273.4]
  assign output_0_26 = io_outValid_26 & _T_15506; // @[Switch.scala 41:38:@5274.4]
  assign _T_15509 = select_27 == 5'h0; // @[Switch.scala 41:52:@5276.4]
  assign output_0_27 = io_outValid_27 & _T_15509; // @[Switch.scala 41:38:@5277.4]
  assign _T_15512 = select_28 == 5'h0; // @[Switch.scala 41:52:@5279.4]
  assign output_0_28 = io_outValid_28 & _T_15512; // @[Switch.scala 41:38:@5280.4]
  assign _T_15515 = select_29 == 5'h0; // @[Switch.scala 41:52:@5282.4]
  assign output_0_29 = io_outValid_29 & _T_15515; // @[Switch.scala 41:38:@5283.4]
  assign _T_15518 = select_30 == 5'h0; // @[Switch.scala 41:52:@5285.4]
  assign output_0_30 = io_outValid_30 & _T_15518; // @[Switch.scala 41:38:@5286.4]
  assign _T_15521 = select_31 == 5'h0; // @[Switch.scala 41:52:@5288.4]
  assign output_0_31 = io_outValid_31 & _T_15521; // @[Switch.scala 41:38:@5289.4]
  assign _T_15529 = {output_0_7,output_0_6,output_0_5,output_0_4,output_0_3,output_0_2,output_0_1,output_0_0}; // @[Switch.scala 43:31:@5297.4]
  assign _T_15537 = {output_0_15,output_0_14,output_0_13,output_0_12,output_0_11,output_0_10,output_0_9,output_0_8,_T_15529}; // @[Switch.scala 43:31:@5305.4]
  assign _T_15544 = {output_0_23,output_0_22,output_0_21,output_0_20,output_0_19,output_0_18,output_0_17,output_0_16}; // @[Switch.scala 43:31:@5312.4]
  assign _T_15553 = {output_0_31,output_0_30,output_0_29,output_0_28,output_0_27,output_0_26,output_0_25,output_0_24,_T_15544,_T_15537}; // @[Switch.scala 43:31:@5321.4]
  assign _T_15557 = select_0 == 5'h1; // @[Switch.scala 41:52:@5324.4]
  assign output_1_0 = io_outValid_0 & _T_15557; // @[Switch.scala 41:38:@5325.4]
  assign _T_15560 = select_1 == 5'h1; // @[Switch.scala 41:52:@5327.4]
  assign output_1_1 = io_outValid_1 & _T_15560; // @[Switch.scala 41:38:@5328.4]
  assign _T_15563 = select_2 == 5'h1; // @[Switch.scala 41:52:@5330.4]
  assign output_1_2 = io_outValid_2 & _T_15563; // @[Switch.scala 41:38:@5331.4]
  assign _T_15566 = select_3 == 5'h1; // @[Switch.scala 41:52:@5333.4]
  assign output_1_3 = io_outValid_3 & _T_15566; // @[Switch.scala 41:38:@5334.4]
  assign _T_15569 = select_4 == 5'h1; // @[Switch.scala 41:52:@5336.4]
  assign output_1_4 = io_outValid_4 & _T_15569; // @[Switch.scala 41:38:@5337.4]
  assign _T_15572 = select_5 == 5'h1; // @[Switch.scala 41:52:@5339.4]
  assign output_1_5 = io_outValid_5 & _T_15572; // @[Switch.scala 41:38:@5340.4]
  assign _T_15575 = select_6 == 5'h1; // @[Switch.scala 41:52:@5342.4]
  assign output_1_6 = io_outValid_6 & _T_15575; // @[Switch.scala 41:38:@5343.4]
  assign _T_15578 = select_7 == 5'h1; // @[Switch.scala 41:52:@5345.4]
  assign output_1_7 = io_outValid_7 & _T_15578; // @[Switch.scala 41:38:@5346.4]
  assign _T_15581 = select_8 == 5'h1; // @[Switch.scala 41:52:@5348.4]
  assign output_1_8 = io_outValid_8 & _T_15581; // @[Switch.scala 41:38:@5349.4]
  assign _T_15584 = select_9 == 5'h1; // @[Switch.scala 41:52:@5351.4]
  assign output_1_9 = io_outValid_9 & _T_15584; // @[Switch.scala 41:38:@5352.4]
  assign _T_15587 = select_10 == 5'h1; // @[Switch.scala 41:52:@5354.4]
  assign output_1_10 = io_outValid_10 & _T_15587; // @[Switch.scala 41:38:@5355.4]
  assign _T_15590 = select_11 == 5'h1; // @[Switch.scala 41:52:@5357.4]
  assign output_1_11 = io_outValid_11 & _T_15590; // @[Switch.scala 41:38:@5358.4]
  assign _T_15593 = select_12 == 5'h1; // @[Switch.scala 41:52:@5360.4]
  assign output_1_12 = io_outValid_12 & _T_15593; // @[Switch.scala 41:38:@5361.4]
  assign _T_15596 = select_13 == 5'h1; // @[Switch.scala 41:52:@5363.4]
  assign output_1_13 = io_outValid_13 & _T_15596; // @[Switch.scala 41:38:@5364.4]
  assign _T_15599 = select_14 == 5'h1; // @[Switch.scala 41:52:@5366.4]
  assign output_1_14 = io_outValid_14 & _T_15599; // @[Switch.scala 41:38:@5367.4]
  assign _T_15602 = select_15 == 5'h1; // @[Switch.scala 41:52:@5369.4]
  assign output_1_15 = io_outValid_15 & _T_15602; // @[Switch.scala 41:38:@5370.4]
  assign _T_15605 = select_16 == 5'h1; // @[Switch.scala 41:52:@5372.4]
  assign output_1_16 = io_outValid_16 & _T_15605; // @[Switch.scala 41:38:@5373.4]
  assign _T_15608 = select_17 == 5'h1; // @[Switch.scala 41:52:@5375.4]
  assign output_1_17 = io_outValid_17 & _T_15608; // @[Switch.scala 41:38:@5376.4]
  assign _T_15611 = select_18 == 5'h1; // @[Switch.scala 41:52:@5378.4]
  assign output_1_18 = io_outValid_18 & _T_15611; // @[Switch.scala 41:38:@5379.4]
  assign _T_15614 = select_19 == 5'h1; // @[Switch.scala 41:52:@5381.4]
  assign output_1_19 = io_outValid_19 & _T_15614; // @[Switch.scala 41:38:@5382.4]
  assign _T_15617 = select_20 == 5'h1; // @[Switch.scala 41:52:@5384.4]
  assign output_1_20 = io_outValid_20 & _T_15617; // @[Switch.scala 41:38:@5385.4]
  assign _T_15620 = select_21 == 5'h1; // @[Switch.scala 41:52:@5387.4]
  assign output_1_21 = io_outValid_21 & _T_15620; // @[Switch.scala 41:38:@5388.4]
  assign _T_15623 = select_22 == 5'h1; // @[Switch.scala 41:52:@5390.4]
  assign output_1_22 = io_outValid_22 & _T_15623; // @[Switch.scala 41:38:@5391.4]
  assign _T_15626 = select_23 == 5'h1; // @[Switch.scala 41:52:@5393.4]
  assign output_1_23 = io_outValid_23 & _T_15626; // @[Switch.scala 41:38:@5394.4]
  assign _T_15629 = select_24 == 5'h1; // @[Switch.scala 41:52:@5396.4]
  assign output_1_24 = io_outValid_24 & _T_15629; // @[Switch.scala 41:38:@5397.4]
  assign _T_15632 = select_25 == 5'h1; // @[Switch.scala 41:52:@5399.4]
  assign output_1_25 = io_outValid_25 & _T_15632; // @[Switch.scala 41:38:@5400.4]
  assign _T_15635 = select_26 == 5'h1; // @[Switch.scala 41:52:@5402.4]
  assign output_1_26 = io_outValid_26 & _T_15635; // @[Switch.scala 41:38:@5403.4]
  assign _T_15638 = select_27 == 5'h1; // @[Switch.scala 41:52:@5405.4]
  assign output_1_27 = io_outValid_27 & _T_15638; // @[Switch.scala 41:38:@5406.4]
  assign _T_15641 = select_28 == 5'h1; // @[Switch.scala 41:52:@5408.4]
  assign output_1_28 = io_outValid_28 & _T_15641; // @[Switch.scala 41:38:@5409.4]
  assign _T_15644 = select_29 == 5'h1; // @[Switch.scala 41:52:@5411.4]
  assign output_1_29 = io_outValid_29 & _T_15644; // @[Switch.scala 41:38:@5412.4]
  assign _T_15647 = select_30 == 5'h1; // @[Switch.scala 41:52:@5414.4]
  assign output_1_30 = io_outValid_30 & _T_15647; // @[Switch.scala 41:38:@5415.4]
  assign _T_15650 = select_31 == 5'h1; // @[Switch.scala 41:52:@5417.4]
  assign output_1_31 = io_outValid_31 & _T_15650; // @[Switch.scala 41:38:@5418.4]
  assign _T_15658 = {output_1_7,output_1_6,output_1_5,output_1_4,output_1_3,output_1_2,output_1_1,output_1_0}; // @[Switch.scala 43:31:@5426.4]
  assign _T_15666 = {output_1_15,output_1_14,output_1_13,output_1_12,output_1_11,output_1_10,output_1_9,output_1_8,_T_15658}; // @[Switch.scala 43:31:@5434.4]
  assign _T_15673 = {output_1_23,output_1_22,output_1_21,output_1_20,output_1_19,output_1_18,output_1_17,output_1_16}; // @[Switch.scala 43:31:@5441.4]
  assign _T_15682 = {output_1_31,output_1_30,output_1_29,output_1_28,output_1_27,output_1_26,output_1_25,output_1_24,_T_15673,_T_15666}; // @[Switch.scala 43:31:@5450.4]
  assign _T_15686 = select_0 == 5'h2; // @[Switch.scala 41:52:@5453.4]
  assign output_2_0 = io_outValid_0 & _T_15686; // @[Switch.scala 41:38:@5454.4]
  assign _T_15689 = select_1 == 5'h2; // @[Switch.scala 41:52:@5456.4]
  assign output_2_1 = io_outValid_1 & _T_15689; // @[Switch.scala 41:38:@5457.4]
  assign _T_15692 = select_2 == 5'h2; // @[Switch.scala 41:52:@5459.4]
  assign output_2_2 = io_outValid_2 & _T_15692; // @[Switch.scala 41:38:@5460.4]
  assign _T_15695 = select_3 == 5'h2; // @[Switch.scala 41:52:@5462.4]
  assign output_2_3 = io_outValid_3 & _T_15695; // @[Switch.scala 41:38:@5463.4]
  assign _T_15698 = select_4 == 5'h2; // @[Switch.scala 41:52:@5465.4]
  assign output_2_4 = io_outValid_4 & _T_15698; // @[Switch.scala 41:38:@5466.4]
  assign _T_15701 = select_5 == 5'h2; // @[Switch.scala 41:52:@5468.4]
  assign output_2_5 = io_outValid_5 & _T_15701; // @[Switch.scala 41:38:@5469.4]
  assign _T_15704 = select_6 == 5'h2; // @[Switch.scala 41:52:@5471.4]
  assign output_2_6 = io_outValid_6 & _T_15704; // @[Switch.scala 41:38:@5472.4]
  assign _T_15707 = select_7 == 5'h2; // @[Switch.scala 41:52:@5474.4]
  assign output_2_7 = io_outValid_7 & _T_15707; // @[Switch.scala 41:38:@5475.4]
  assign _T_15710 = select_8 == 5'h2; // @[Switch.scala 41:52:@5477.4]
  assign output_2_8 = io_outValid_8 & _T_15710; // @[Switch.scala 41:38:@5478.4]
  assign _T_15713 = select_9 == 5'h2; // @[Switch.scala 41:52:@5480.4]
  assign output_2_9 = io_outValid_9 & _T_15713; // @[Switch.scala 41:38:@5481.4]
  assign _T_15716 = select_10 == 5'h2; // @[Switch.scala 41:52:@5483.4]
  assign output_2_10 = io_outValid_10 & _T_15716; // @[Switch.scala 41:38:@5484.4]
  assign _T_15719 = select_11 == 5'h2; // @[Switch.scala 41:52:@5486.4]
  assign output_2_11 = io_outValid_11 & _T_15719; // @[Switch.scala 41:38:@5487.4]
  assign _T_15722 = select_12 == 5'h2; // @[Switch.scala 41:52:@5489.4]
  assign output_2_12 = io_outValid_12 & _T_15722; // @[Switch.scala 41:38:@5490.4]
  assign _T_15725 = select_13 == 5'h2; // @[Switch.scala 41:52:@5492.4]
  assign output_2_13 = io_outValid_13 & _T_15725; // @[Switch.scala 41:38:@5493.4]
  assign _T_15728 = select_14 == 5'h2; // @[Switch.scala 41:52:@5495.4]
  assign output_2_14 = io_outValid_14 & _T_15728; // @[Switch.scala 41:38:@5496.4]
  assign _T_15731 = select_15 == 5'h2; // @[Switch.scala 41:52:@5498.4]
  assign output_2_15 = io_outValid_15 & _T_15731; // @[Switch.scala 41:38:@5499.4]
  assign _T_15734 = select_16 == 5'h2; // @[Switch.scala 41:52:@5501.4]
  assign output_2_16 = io_outValid_16 & _T_15734; // @[Switch.scala 41:38:@5502.4]
  assign _T_15737 = select_17 == 5'h2; // @[Switch.scala 41:52:@5504.4]
  assign output_2_17 = io_outValid_17 & _T_15737; // @[Switch.scala 41:38:@5505.4]
  assign _T_15740 = select_18 == 5'h2; // @[Switch.scala 41:52:@5507.4]
  assign output_2_18 = io_outValid_18 & _T_15740; // @[Switch.scala 41:38:@5508.4]
  assign _T_15743 = select_19 == 5'h2; // @[Switch.scala 41:52:@5510.4]
  assign output_2_19 = io_outValid_19 & _T_15743; // @[Switch.scala 41:38:@5511.4]
  assign _T_15746 = select_20 == 5'h2; // @[Switch.scala 41:52:@5513.4]
  assign output_2_20 = io_outValid_20 & _T_15746; // @[Switch.scala 41:38:@5514.4]
  assign _T_15749 = select_21 == 5'h2; // @[Switch.scala 41:52:@5516.4]
  assign output_2_21 = io_outValid_21 & _T_15749; // @[Switch.scala 41:38:@5517.4]
  assign _T_15752 = select_22 == 5'h2; // @[Switch.scala 41:52:@5519.4]
  assign output_2_22 = io_outValid_22 & _T_15752; // @[Switch.scala 41:38:@5520.4]
  assign _T_15755 = select_23 == 5'h2; // @[Switch.scala 41:52:@5522.4]
  assign output_2_23 = io_outValid_23 & _T_15755; // @[Switch.scala 41:38:@5523.4]
  assign _T_15758 = select_24 == 5'h2; // @[Switch.scala 41:52:@5525.4]
  assign output_2_24 = io_outValid_24 & _T_15758; // @[Switch.scala 41:38:@5526.4]
  assign _T_15761 = select_25 == 5'h2; // @[Switch.scala 41:52:@5528.4]
  assign output_2_25 = io_outValid_25 & _T_15761; // @[Switch.scala 41:38:@5529.4]
  assign _T_15764 = select_26 == 5'h2; // @[Switch.scala 41:52:@5531.4]
  assign output_2_26 = io_outValid_26 & _T_15764; // @[Switch.scala 41:38:@5532.4]
  assign _T_15767 = select_27 == 5'h2; // @[Switch.scala 41:52:@5534.4]
  assign output_2_27 = io_outValid_27 & _T_15767; // @[Switch.scala 41:38:@5535.4]
  assign _T_15770 = select_28 == 5'h2; // @[Switch.scala 41:52:@5537.4]
  assign output_2_28 = io_outValid_28 & _T_15770; // @[Switch.scala 41:38:@5538.4]
  assign _T_15773 = select_29 == 5'h2; // @[Switch.scala 41:52:@5540.4]
  assign output_2_29 = io_outValid_29 & _T_15773; // @[Switch.scala 41:38:@5541.4]
  assign _T_15776 = select_30 == 5'h2; // @[Switch.scala 41:52:@5543.4]
  assign output_2_30 = io_outValid_30 & _T_15776; // @[Switch.scala 41:38:@5544.4]
  assign _T_15779 = select_31 == 5'h2; // @[Switch.scala 41:52:@5546.4]
  assign output_2_31 = io_outValid_31 & _T_15779; // @[Switch.scala 41:38:@5547.4]
  assign _T_15787 = {output_2_7,output_2_6,output_2_5,output_2_4,output_2_3,output_2_2,output_2_1,output_2_0}; // @[Switch.scala 43:31:@5555.4]
  assign _T_15795 = {output_2_15,output_2_14,output_2_13,output_2_12,output_2_11,output_2_10,output_2_9,output_2_8,_T_15787}; // @[Switch.scala 43:31:@5563.4]
  assign _T_15802 = {output_2_23,output_2_22,output_2_21,output_2_20,output_2_19,output_2_18,output_2_17,output_2_16}; // @[Switch.scala 43:31:@5570.4]
  assign _T_15811 = {output_2_31,output_2_30,output_2_29,output_2_28,output_2_27,output_2_26,output_2_25,output_2_24,_T_15802,_T_15795}; // @[Switch.scala 43:31:@5579.4]
  assign _T_15815 = select_0 == 5'h3; // @[Switch.scala 41:52:@5582.4]
  assign output_3_0 = io_outValid_0 & _T_15815; // @[Switch.scala 41:38:@5583.4]
  assign _T_15818 = select_1 == 5'h3; // @[Switch.scala 41:52:@5585.4]
  assign output_3_1 = io_outValid_1 & _T_15818; // @[Switch.scala 41:38:@5586.4]
  assign _T_15821 = select_2 == 5'h3; // @[Switch.scala 41:52:@5588.4]
  assign output_3_2 = io_outValid_2 & _T_15821; // @[Switch.scala 41:38:@5589.4]
  assign _T_15824 = select_3 == 5'h3; // @[Switch.scala 41:52:@5591.4]
  assign output_3_3 = io_outValid_3 & _T_15824; // @[Switch.scala 41:38:@5592.4]
  assign _T_15827 = select_4 == 5'h3; // @[Switch.scala 41:52:@5594.4]
  assign output_3_4 = io_outValid_4 & _T_15827; // @[Switch.scala 41:38:@5595.4]
  assign _T_15830 = select_5 == 5'h3; // @[Switch.scala 41:52:@5597.4]
  assign output_3_5 = io_outValid_5 & _T_15830; // @[Switch.scala 41:38:@5598.4]
  assign _T_15833 = select_6 == 5'h3; // @[Switch.scala 41:52:@5600.4]
  assign output_3_6 = io_outValid_6 & _T_15833; // @[Switch.scala 41:38:@5601.4]
  assign _T_15836 = select_7 == 5'h3; // @[Switch.scala 41:52:@5603.4]
  assign output_3_7 = io_outValid_7 & _T_15836; // @[Switch.scala 41:38:@5604.4]
  assign _T_15839 = select_8 == 5'h3; // @[Switch.scala 41:52:@5606.4]
  assign output_3_8 = io_outValid_8 & _T_15839; // @[Switch.scala 41:38:@5607.4]
  assign _T_15842 = select_9 == 5'h3; // @[Switch.scala 41:52:@5609.4]
  assign output_3_9 = io_outValid_9 & _T_15842; // @[Switch.scala 41:38:@5610.4]
  assign _T_15845 = select_10 == 5'h3; // @[Switch.scala 41:52:@5612.4]
  assign output_3_10 = io_outValid_10 & _T_15845; // @[Switch.scala 41:38:@5613.4]
  assign _T_15848 = select_11 == 5'h3; // @[Switch.scala 41:52:@5615.4]
  assign output_3_11 = io_outValid_11 & _T_15848; // @[Switch.scala 41:38:@5616.4]
  assign _T_15851 = select_12 == 5'h3; // @[Switch.scala 41:52:@5618.4]
  assign output_3_12 = io_outValid_12 & _T_15851; // @[Switch.scala 41:38:@5619.4]
  assign _T_15854 = select_13 == 5'h3; // @[Switch.scala 41:52:@5621.4]
  assign output_3_13 = io_outValid_13 & _T_15854; // @[Switch.scala 41:38:@5622.4]
  assign _T_15857 = select_14 == 5'h3; // @[Switch.scala 41:52:@5624.4]
  assign output_3_14 = io_outValid_14 & _T_15857; // @[Switch.scala 41:38:@5625.4]
  assign _T_15860 = select_15 == 5'h3; // @[Switch.scala 41:52:@5627.4]
  assign output_3_15 = io_outValid_15 & _T_15860; // @[Switch.scala 41:38:@5628.4]
  assign _T_15863 = select_16 == 5'h3; // @[Switch.scala 41:52:@5630.4]
  assign output_3_16 = io_outValid_16 & _T_15863; // @[Switch.scala 41:38:@5631.4]
  assign _T_15866 = select_17 == 5'h3; // @[Switch.scala 41:52:@5633.4]
  assign output_3_17 = io_outValid_17 & _T_15866; // @[Switch.scala 41:38:@5634.4]
  assign _T_15869 = select_18 == 5'h3; // @[Switch.scala 41:52:@5636.4]
  assign output_3_18 = io_outValid_18 & _T_15869; // @[Switch.scala 41:38:@5637.4]
  assign _T_15872 = select_19 == 5'h3; // @[Switch.scala 41:52:@5639.4]
  assign output_3_19 = io_outValid_19 & _T_15872; // @[Switch.scala 41:38:@5640.4]
  assign _T_15875 = select_20 == 5'h3; // @[Switch.scala 41:52:@5642.4]
  assign output_3_20 = io_outValid_20 & _T_15875; // @[Switch.scala 41:38:@5643.4]
  assign _T_15878 = select_21 == 5'h3; // @[Switch.scala 41:52:@5645.4]
  assign output_3_21 = io_outValid_21 & _T_15878; // @[Switch.scala 41:38:@5646.4]
  assign _T_15881 = select_22 == 5'h3; // @[Switch.scala 41:52:@5648.4]
  assign output_3_22 = io_outValid_22 & _T_15881; // @[Switch.scala 41:38:@5649.4]
  assign _T_15884 = select_23 == 5'h3; // @[Switch.scala 41:52:@5651.4]
  assign output_3_23 = io_outValid_23 & _T_15884; // @[Switch.scala 41:38:@5652.4]
  assign _T_15887 = select_24 == 5'h3; // @[Switch.scala 41:52:@5654.4]
  assign output_3_24 = io_outValid_24 & _T_15887; // @[Switch.scala 41:38:@5655.4]
  assign _T_15890 = select_25 == 5'h3; // @[Switch.scala 41:52:@5657.4]
  assign output_3_25 = io_outValid_25 & _T_15890; // @[Switch.scala 41:38:@5658.4]
  assign _T_15893 = select_26 == 5'h3; // @[Switch.scala 41:52:@5660.4]
  assign output_3_26 = io_outValid_26 & _T_15893; // @[Switch.scala 41:38:@5661.4]
  assign _T_15896 = select_27 == 5'h3; // @[Switch.scala 41:52:@5663.4]
  assign output_3_27 = io_outValid_27 & _T_15896; // @[Switch.scala 41:38:@5664.4]
  assign _T_15899 = select_28 == 5'h3; // @[Switch.scala 41:52:@5666.4]
  assign output_3_28 = io_outValid_28 & _T_15899; // @[Switch.scala 41:38:@5667.4]
  assign _T_15902 = select_29 == 5'h3; // @[Switch.scala 41:52:@5669.4]
  assign output_3_29 = io_outValid_29 & _T_15902; // @[Switch.scala 41:38:@5670.4]
  assign _T_15905 = select_30 == 5'h3; // @[Switch.scala 41:52:@5672.4]
  assign output_3_30 = io_outValid_30 & _T_15905; // @[Switch.scala 41:38:@5673.4]
  assign _T_15908 = select_31 == 5'h3; // @[Switch.scala 41:52:@5675.4]
  assign output_3_31 = io_outValid_31 & _T_15908; // @[Switch.scala 41:38:@5676.4]
  assign _T_15916 = {output_3_7,output_3_6,output_3_5,output_3_4,output_3_3,output_3_2,output_3_1,output_3_0}; // @[Switch.scala 43:31:@5684.4]
  assign _T_15924 = {output_3_15,output_3_14,output_3_13,output_3_12,output_3_11,output_3_10,output_3_9,output_3_8,_T_15916}; // @[Switch.scala 43:31:@5692.4]
  assign _T_15931 = {output_3_23,output_3_22,output_3_21,output_3_20,output_3_19,output_3_18,output_3_17,output_3_16}; // @[Switch.scala 43:31:@5699.4]
  assign _T_15940 = {output_3_31,output_3_30,output_3_29,output_3_28,output_3_27,output_3_26,output_3_25,output_3_24,_T_15931,_T_15924}; // @[Switch.scala 43:31:@5708.4]
  assign _T_15944 = select_0 == 5'h4; // @[Switch.scala 41:52:@5711.4]
  assign output_4_0 = io_outValid_0 & _T_15944; // @[Switch.scala 41:38:@5712.4]
  assign _T_15947 = select_1 == 5'h4; // @[Switch.scala 41:52:@5714.4]
  assign output_4_1 = io_outValid_1 & _T_15947; // @[Switch.scala 41:38:@5715.4]
  assign _T_15950 = select_2 == 5'h4; // @[Switch.scala 41:52:@5717.4]
  assign output_4_2 = io_outValid_2 & _T_15950; // @[Switch.scala 41:38:@5718.4]
  assign _T_15953 = select_3 == 5'h4; // @[Switch.scala 41:52:@5720.4]
  assign output_4_3 = io_outValid_3 & _T_15953; // @[Switch.scala 41:38:@5721.4]
  assign _T_15956 = select_4 == 5'h4; // @[Switch.scala 41:52:@5723.4]
  assign output_4_4 = io_outValid_4 & _T_15956; // @[Switch.scala 41:38:@5724.4]
  assign _T_15959 = select_5 == 5'h4; // @[Switch.scala 41:52:@5726.4]
  assign output_4_5 = io_outValid_5 & _T_15959; // @[Switch.scala 41:38:@5727.4]
  assign _T_15962 = select_6 == 5'h4; // @[Switch.scala 41:52:@5729.4]
  assign output_4_6 = io_outValid_6 & _T_15962; // @[Switch.scala 41:38:@5730.4]
  assign _T_15965 = select_7 == 5'h4; // @[Switch.scala 41:52:@5732.4]
  assign output_4_7 = io_outValid_7 & _T_15965; // @[Switch.scala 41:38:@5733.4]
  assign _T_15968 = select_8 == 5'h4; // @[Switch.scala 41:52:@5735.4]
  assign output_4_8 = io_outValid_8 & _T_15968; // @[Switch.scala 41:38:@5736.4]
  assign _T_15971 = select_9 == 5'h4; // @[Switch.scala 41:52:@5738.4]
  assign output_4_9 = io_outValid_9 & _T_15971; // @[Switch.scala 41:38:@5739.4]
  assign _T_15974 = select_10 == 5'h4; // @[Switch.scala 41:52:@5741.4]
  assign output_4_10 = io_outValid_10 & _T_15974; // @[Switch.scala 41:38:@5742.4]
  assign _T_15977 = select_11 == 5'h4; // @[Switch.scala 41:52:@5744.4]
  assign output_4_11 = io_outValid_11 & _T_15977; // @[Switch.scala 41:38:@5745.4]
  assign _T_15980 = select_12 == 5'h4; // @[Switch.scala 41:52:@5747.4]
  assign output_4_12 = io_outValid_12 & _T_15980; // @[Switch.scala 41:38:@5748.4]
  assign _T_15983 = select_13 == 5'h4; // @[Switch.scala 41:52:@5750.4]
  assign output_4_13 = io_outValid_13 & _T_15983; // @[Switch.scala 41:38:@5751.4]
  assign _T_15986 = select_14 == 5'h4; // @[Switch.scala 41:52:@5753.4]
  assign output_4_14 = io_outValid_14 & _T_15986; // @[Switch.scala 41:38:@5754.4]
  assign _T_15989 = select_15 == 5'h4; // @[Switch.scala 41:52:@5756.4]
  assign output_4_15 = io_outValid_15 & _T_15989; // @[Switch.scala 41:38:@5757.4]
  assign _T_15992 = select_16 == 5'h4; // @[Switch.scala 41:52:@5759.4]
  assign output_4_16 = io_outValid_16 & _T_15992; // @[Switch.scala 41:38:@5760.4]
  assign _T_15995 = select_17 == 5'h4; // @[Switch.scala 41:52:@5762.4]
  assign output_4_17 = io_outValid_17 & _T_15995; // @[Switch.scala 41:38:@5763.4]
  assign _T_15998 = select_18 == 5'h4; // @[Switch.scala 41:52:@5765.4]
  assign output_4_18 = io_outValid_18 & _T_15998; // @[Switch.scala 41:38:@5766.4]
  assign _T_16001 = select_19 == 5'h4; // @[Switch.scala 41:52:@5768.4]
  assign output_4_19 = io_outValid_19 & _T_16001; // @[Switch.scala 41:38:@5769.4]
  assign _T_16004 = select_20 == 5'h4; // @[Switch.scala 41:52:@5771.4]
  assign output_4_20 = io_outValid_20 & _T_16004; // @[Switch.scala 41:38:@5772.4]
  assign _T_16007 = select_21 == 5'h4; // @[Switch.scala 41:52:@5774.4]
  assign output_4_21 = io_outValid_21 & _T_16007; // @[Switch.scala 41:38:@5775.4]
  assign _T_16010 = select_22 == 5'h4; // @[Switch.scala 41:52:@5777.4]
  assign output_4_22 = io_outValid_22 & _T_16010; // @[Switch.scala 41:38:@5778.4]
  assign _T_16013 = select_23 == 5'h4; // @[Switch.scala 41:52:@5780.4]
  assign output_4_23 = io_outValid_23 & _T_16013; // @[Switch.scala 41:38:@5781.4]
  assign _T_16016 = select_24 == 5'h4; // @[Switch.scala 41:52:@5783.4]
  assign output_4_24 = io_outValid_24 & _T_16016; // @[Switch.scala 41:38:@5784.4]
  assign _T_16019 = select_25 == 5'h4; // @[Switch.scala 41:52:@5786.4]
  assign output_4_25 = io_outValid_25 & _T_16019; // @[Switch.scala 41:38:@5787.4]
  assign _T_16022 = select_26 == 5'h4; // @[Switch.scala 41:52:@5789.4]
  assign output_4_26 = io_outValid_26 & _T_16022; // @[Switch.scala 41:38:@5790.4]
  assign _T_16025 = select_27 == 5'h4; // @[Switch.scala 41:52:@5792.4]
  assign output_4_27 = io_outValid_27 & _T_16025; // @[Switch.scala 41:38:@5793.4]
  assign _T_16028 = select_28 == 5'h4; // @[Switch.scala 41:52:@5795.4]
  assign output_4_28 = io_outValid_28 & _T_16028; // @[Switch.scala 41:38:@5796.4]
  assign _T_16031 = select_29 == 5'h4; // @[Switch.scala 41:52:@5798.4]
  assign output_4_29 = io_outValid_29 & _T_16031; // @[Switch.scala 41:38:@5799.4]
  assign _T_16034 = select_30 == 5'h4; // @[Switch.scala 41:52:@5801.4]
  assign output_4_30 = io_outValid_30 & _T_16034; // @[Switch.scala 41:38:@5802.4]
  assign _T_16037 = select_31 == 5'h4; // @[Switch.scala 41:52:@5804.4]
  assign output_4_31 = io_outValid_31 & _T_16037; // @[Switch.scala 41:38:@5805.4]
  assign _T_16045 = {output_4_7,output_4_6,output_4_5,output_4_4,output_4_3,output_4_2,output_4_1,output_4_0}; // @[Switch.scala 43:31:@5813.4]
  assign _T_16053 = {output_4_15,output_4_14,output_4_13,output_4_12,output_4_11,output_4_10,output_4_9,output_4_8,_T_16045}; // @[Switch.scala 43:31:@5821.4]
  assign _T_16060 = {output_4_23,output_4_22,output_4_21,output_4_20,output_4_19,output_4_18,output_4_17,output_4_16}; // @[Switch.scala 43:31:@5828.4]
  assign _T_16069 = {output_4_31,output_4_30,output_4_29,output_4_28,output_4_27,output_4_26,output_4_25,output_4_24,_T_16060,_T_16053}; // @[Switch.scala 43:31:@5837.4]
  assign _T_16073 = select_0 == 5'h5; // @[Switch.scala 41:52:@5840.4]
  assign output_5_0 = io_outValid_0 & _T_16073; // @[Switch.scala 41:38:@5841.4]
  assign _T_16076 = select_1 == 5'h5; // @[Switch.scala 41:52:@5843.4]
  assign output_5_1 = io_outValid_1 & _T_16076; // @[Switch.scala 41:38:@5844.4]
  assign _T_16079 = select_2 == 5'h5; // @[Switch.scala 41:52:@5846.4]
  assign output_5_2 = io_outValid_2 & _T_16079; // @[Switch.scala 41:38:@5847.4]
  assign _T_16082 = select_3 == 5'h5; // @[Switch.scala 41:52:@5849.4]
  assign output_5_3 = io_outValid_3 & _T_16082; // @[Switch.scala 41:38:@5850.4]
  assign _T_16085 = select_4 == 5'h5; // @[Switch.scala 41:52:@5852.4]
  assign output_5_4 = io_outValid_4 & _T_16085; // @[Switch.scala 41:38:@5853.4]
  assign _T_16088 = select_5 == 5'h5; // @[Switch.scala 41:52:@5855.4]
  assign output_5_5 = io_outValid_5 & _T_16088; // @[Switch.scala 41:38:@5856.4]
  assign _T_16091 = select_6 == 5'h5; // @[Switch.scala 41:52:@5858.4]
  assign output_5_6 = io_outValid_6 & _T_16091; // @[Switch.scala 41:38:@5859.4]
  assign _T_16094 = select_7 == 5'h5; // @[Switch.scala 41:52:@5861.4]
  assign output_5_7 = io_outValid_7 & _T_16094; // @[Switch.scala 41:38:@5862.4]
  assign _T_16097 = select_8 == 5'h5; // @[Switch.scala 41:52:@5864.4]
  assign output_5_8 = io_outValid_8 & _T_16097; // @[Switch.scala 41:38:@5865.4]
  assign _T_16100 = select_9 == 5'h5; // @[Switch.scala 41:52:@5867.4]
  assign output_5_9 = io_outValid_9 & _T_16100; // @[Switch.scala 41:38:@5868.4]
  assign _T_16103 = select_10 == 5'h5; // @[Switch.scala 41:52:@5870.4]
  assign output_5_10 = io_outValid_10 & _T_16103; // @[Switch.scala 41:38:@5871.4]
  assign _T_16106 = select_11 == 5'h5; // @[Switch.scala 41:52:@5873.4]
  assign output_5_11 = io_outValid_11 & _T_16106; // @[Switch.scala 41:38:@5874.4]
  assign _T_16109 = select_12 == 5'h5; // @[Switch.scala 41:52:@5876.4]
  assign output_5_12 = io_outValid_12 & _T_16109; // @[Switch.scala 41:38:@5877.4]
  assign _T_16112 = select_13 == 5'h5; // @[Switch.scala 41:52:@5879.4]
  assign output_5_13 = io_outValid_13 & _T_16112; // @[Switch.scala 41:38:@5880.4]
  assign _T_16115 = select_14 == 5'h5; // @[Switch.scala 41:52:@5882.4]
  assign output_5_14 = io_outValid_14 & _T_16115; // @[Switch.scala 41:38:@5883.4]
  assign _T_16118 = select_15 == 5'h5; // @[Switch.scala 41:52:@5885.4]
  assign output_5_15 = io_outValid_15 & _T_16118; // @[Switch.scala 41:38:@5886.4]
  assign _T_16121 = select_16 == 5'h5; // @[Switch.scala 41:52:@5888.4]
  assign output_5_16 = io_outValid_16 & _T_16121; // @[Switch.scala 41:38:@5889.4]
  assign _T_16124 = select_17 == 5'h5; // @[Switch.scala 41:52:@5891.4]
  assign output_5_17 = io_outValid_17 & _T_16124; // @[Switch.scala 41:38:@5892.4]
  assign _T_16127 = select_18 == 5'h5; // @[Switch.scala 41:52:@5894.4]
  assign output_5_18 = io_outValid_18 & _T_16127; // @[Switch.scala 41:38:@5895.4]
  assign _T_16130 = select_19 == 5'h5; // @[Switch.scala 41:52:@5897.4]
  assign output_5_19 = io_outValid_19 & _T_16130; // @[Switch.scala 41:38:@5898.4]
  assign _T_16133 = select_20 == 5'h5; // @[Switch.scala 41:52:@5900.4]
  assign output_5_20 = io_outValid_20 & _T_16133; // @[Switch.scala 41:38:@5901.4]
  assign _T_16136 = select_21 == 5'h5; // @[Switch.scala 41:52:@5903.4]
  assign output_5_21 = io_outValid_21 & _T_16136; // @[Switch.scala 41:38:@5904.4]
  assign _T_16139 = select_22 == 5'h5; // @[Switch.scala 41:52:@5906.4]
  assign output_5_22 = io_outValid_22 & _T_16139; // @[Switch.scala 41:38:@5907.4]
  assign _T_16142 = select_23 == 5'h5; // @[Switch.scala 41:52:@5909.4]
  assign output_5_23 = io_outValid_23 & _T_16142; // @[Switch.scala 41:38:@5910.4]
  assign _T_16145 = select_24 == 5'h5; // @[Switch.scala 41:52:@5912.4]
  assign output_5_24 = io_outValid_24 & _T_16145; // @[Switch.scala 41:38:@5913.4]
  assign _T_16148 = select_25 == 5'h5; // @[Switch.scala 41:52:@5915.4]
  assign output_5_25 = io_outValid_25 & _T_16148; // @[Switch.scala 41:38:@5916.4]
  assign _T_16151 = select_26 == 5'h5; // @[Switch.scala 41:52:@5918.4]
  assign output_5_26 = io_outValid_26 & _T_16151; // @[Switch.scala 41:38:@5919.4]
  assign _T_16154 = select_27 == 5'h5; // @[Switch.scala 41:52:@5921.4]
  assign output_5_27 = io_outValid_27 & _T_16154; // @[Switch.scala 41:38:@5922.4]
  assign _T_16157 = select_28 == 5'h5; // @[Switch.scala 41:52:@5924.4]
  assign output_5_28 = io_outValid_28 & _T_16157; // @[Switch.scala 41:38:@5925.4]
  assign _T_16160 = select_29 == 5'h5; // @[Switch.scala 41:52:@5927.4]
  assign output_5_29 = io_outValid_29 & _T_16160; // @[Switch.scala 41:38:@5928.4]
  assign _T_16163 = select_30 == 5'h5; // @[Switch.scala 41:52:@5930.4]
  assign output_5_30 = io_outValid_30 & _T_16163; // @[Switch.scala 41:38:@5931.4]
  assign _T_16166 = select_31 == 5'h5; // @[Switch.scala 41:52:@5933.4]
  assign output_5_31 = io_outValid_31 & _T_16166; // @[Switch.scala 41:38:@5934.4]
  assign _T_16174 = {output_5_7,output_5_6,output_5_5,output_5_4,output_5_3,output_5_2,output_5_1,output_5_0}; // @[Switch.scala 43:31:@5942.4]
  assign _T_16182 = {output_5_15,output_5_14,output_5_13,output_5_12,output_5_11,output_5_10,output_5_9,output_5_8,_T_16174}; // @[Switch.scala 43:31:@5950.4]
  assign _T_16189 = {output_5_23,output_5_22,output_5_21,output_5_20,output_5_19,output_5_18,output_5_17,output_5_16}; // @[Switch.scala 43:31:@5957.4]
  assign _T_16198 = {output_5_31,output_5_30,output_5_29,output_5_28,output_5_27,output_5_26,output_5_25,output_5_24,_T_16189,_T_16182}; // @[Switch.scala 43:31:@5966.4]
  assign _T_16202 = select_0 == 5'h6; // @[Switch.scala 41:52:@5969.4]
  assign output_6_0 = io_outValid_0 & _T_16202; // @[Switch.scala 41:38:@5970.4]
  assign _T_16205 = select_1 == 5'h6; // @[Switch.scala 41:52:@5972.4]
  assign output_6_1 = io_outValid_1 & _T_16205; // @[Switch.scala 41:38:@5973.4]
  assign _T_16208 = select_2 == 5'h6; // @[Switch.scala 41:52:@5975.4]
  assign output_6_2 = io_outValid_2 & _T_16208; // @[Switch.scala 41:38:@5976.4]
  assign _T_16211 = select_3 == 5'h6; // @[Switch.scala 41:52:@5978.4]
  assign output_6_3 = io_outValid_3 & _T_16211; // @[Switch.scala 41:38:@5979.4]
  assign _T_16214 = select_4 == 5'h6; // @[Switch.scala 41:52:@5981.4]
  assign output_6_4 = io_outValid_4 & _T_16214; // @[Switch.scala 41:38:@5982.4]
  assign _T_16217 = select_5 == 5'h6; // @[Switch.scala 41:52:@5984.4]
  assign output_6_5 = io_outValid_5 & _T_16217; // @[Switch.scala 41:38:@5985.4]
  assign _T_16220 = select_6 == 5'h6; // @[Switch.scala 41:52:@5987.4]
  assign output_6_6 = io_outValid_6 & _T_16220; // @[Switch.scala 41:38:@5988.4]
  assign _T_16223 = select_7 == 5'h6; // @[Switch.scala 41:52:@5990.4]
  assign output_6_7 = io_outValid_7 & _T_16223; // @[Switch.scala 41:38:@5991.4]
  assign _T_16226 = select_8 == 5'h6; // @[Switch.scala 41:52:@5993.4]
  assign output_6_8 = io_outValid_8 & _T_16226; // @[Switch.scala 41:38:@5994.4]
  assign _T_16229 = select_9 == 5'h6; // @[Switch.scala 41:52:@5996.4]
  assign output_6_9 = io_outValid_9 & _T_16229; // @[Switch.scala 41:38:@5997.4]
  assign _T_16232 = select_10 == 5'h6; // @[Switch.scala 41:52:@5999.4]
  assign output_6_10 = io_outValid_10 & _T_16232; // @[Switch.scala 41:38:@6000.4]
  assign _T_16235 = select_11 == 5'h6; // @[Switch.scala 41:52:@6002.4]
  assign output_6_11 = io_outValid_11 & _T_16235; // @[Switch.scala 41:38:@6003.4]
  assign _T_16238 = select_12 == 5'h6; // @[Switch.scala 41:52:@6005.4]
  assign output_6_12 = io_outValid_12 & _T_16238; // @[Switch.scala 41:38:@6006.4]
  assign _T_16241 = select_13 == 5'h6; // @[Switch.scala 41:52:@6008.4]
  assign output_6_13 = io_outValid_13 & _T_16241; // @[Switch.scala 41:38:@6009.4]
  assign _T_16244 = select_14 == 5'h6; // @[Switch.scala 41:52:@6011.4]
  assign output_6_14 = io_outValid_14 & _T_16244; // @[Switch.scala 41:38:@6012.4]
  assign _T_16247 = select_15 == 5'h6; // @[Switch.scala 41:52:@6014.4]
  assign output_6_15 = io_outValid_15 & _T_16247; // @[Switch.scala 41:38:@6015.4]
  assign _T_16250 = select_16 == 5'h6; // @[Switch.scala 41:52:@6017.4]
  assign output_6_16 = io_outValid_16 & _T_16250; // @[Switch.scala 41:38:@6018.4]
  assign _T_16253 = select_17 == 5'h6; // @[Switch.scala 41:52:@6020.4]
  assign output_6_17 = io_outValid_17 & _T_16253; // @[Switch.scala 41:38:@6021.4]
  assign _T_16256 = select_18 == 5'h6; // @[Switch.scala 41:52:@6023.4]
  assign output_6_18 = io_outValid_18 & _T_16256; // @[Switch.scala 41:38:@6024.4]
  assign _T_16259 = select_19 == 5'h6; // @[Switch.scala 41:52:@6026.4]
  assign output_6_19 = io_outValid_19 & _T_16259; // @[Switch.scala 41:38:@6027.4]
  assign _T_16262 = select_20 == 5'h6; // @[Switch.scala 41:52:@6029.4]
  assign output_6_20 = io_outValid_20 & _T_16262; // @[Switch.scala 41:38:@6030.4]
  assign _T_16265 = select_21 == 5'h6; // @[Switch.scala 41:52:@6032.4]
  assign output_6_21 = io_outValid_21 & _T_16265; // @[Switch.scala 41:38:@6033.4]
  assign _T_16268 = select_22 == 5'h6; // @[Switch.scala 41:52:@6035.4]
  assign output_6_22 = io_outValid_22 & _T_16268; // @[Switch.scala 41:38:@6036.4]
  assign _T_16271 = select_23 == 5'h6; // @[Switch.scala 41:52:@6038.4]
  assign output_6_23 = io_outValid_23 & _T_16271; // @[Switch.scala 41:38:@6039.4]
  assign _T_16274 = select_24 == 5'h6; // @[Switch.scala 41:52:@6041.4]
  assign output_6_24 = io_outValid_24 & _T_16274; // @[Switch.scala 41:38:@6042.4]
  assign _T_16277 = select_25 == 5'h6; // @[Switch.scala 41:52:@6044.4]
  assign output_6_25 = io_outValid_25 & _T_16277; // @[Switch.scala 41:38:@6045.4]
  assign _T_16280 = select_26 == 5'h6; // @[Switch.scala 41:52:@6047.4]
  assign output_6_26 = io_outValid_26 & _T_16280; // @[Switch.scala 41:38:@6048.4]
  assign _T_16283 = select_27 == 5'h6; // @[Switch.scala 41:52:@6050.4]
  assign output_6_27 = io_outValid_27 & _T_16283; // @[Switch.scala 41:38:@6051.4]
  assign _T_16286 = select_28 == 5'h6; // @[Switch.scala 41:52:@6053.4]
  assign output_6_28 = io_outValid_28 & _T_16286; // @[Switch.scala 41:38:@6054.4]
  assign _T_16289 = select_29 == 5'h6; // @[Switch.scala 41:52:@6056.4]
  assign output_6_29 = io_outValid_29 & _T_16289; // @[Switch.scala 41:38:@6057.4]
  assign _T_16292 = select_30 == 5'h6; // @[Switch.scala 41:52:@6059.4]
  assign output_6_30 = io_outValid_30 & _T_16292; // @[Switch.scala 41:38:@6060.4]
  assign _T_16295 = select_31 == 5'h6; // @[Switch.scala 41:52:@6062.4]
  assign output_6_31 = io_outValid_31 & _T_16295; // @[Switch.scala 41:38:@6063.4]
  assign _T_16303 = {output_6_7,output_6_6,output_6_5,output_6_4,output_6_3,output_6_2,output_6_1,output_6_0}; // @[Switch.scala 43:31:@6071.4]
  assign _T_16311 = {output_6_15,output_6_14,output_6_13,output_6_12,output_6_11,output_6_10,output_6_9,output_6_8,_T_16303}; // @[Switch.scala 43:31:@6079.4]
  assign _T_16318 = {output_6_23,output_6_22,output_6_21,output_6_20,output_6_19,output_6_18,output_6_17,output_6_16}; // @[Switch.scala 43:31:@6086.4]
  assign _T_16327 = {output_6_31,output_6_30,output_6_29,output_6_28,output_6_27,output_6_26,output_6_25,output_6_24,_T_16318,_T_16311}; // @[Switch.scala 43:31:@6095.4]
  assign _T_16331 = select_0 == 5'h7; // @[Switch.scala 41:52:@6098.4]
  assign output_7_0 = io_outValid_0 & _T_16331; // @[Switch.scala 41:38:@6099.4]
  assign _T_16334 = select_1 == 5'h7; // @[Switch.scala 41:52:@6101.4]
  assign output_7_1 = io_outValid_1 & _T_16334; // @[Switch.scala 41:38:@6102.4]
  assign _T_16337 = select_2 == 5'h7; // @[Switch.scala 41:52:@6104.4]
  assign output_7_2 = io_outValid_2 & _T_16337; // @[Switch.scala 41:38:@6105.4]
  assign _T_16340 = select_3 == 5'h7; // @[Switch.scala 41:52:@6107.4]
  assign output_7_3 = io_outValid_3 & _T_16340; // @[Switch.scala 41:38:@6108.4]
  assign _T_16343 = select_4 == 5'h7; // @[Switch.scala 41:52:@6110.4]
  assign output_7_4 = io_outValid_4 & _T_16343; // @[Switch.scala 41:38:@6111.4]
  assign _T_16346 = select_5 == 5'h7; // @[Switch.scala 41:52:@6113.4]
  assign output_7_5 = io_outValid_5 & _T_16346; // @[Switch.scala 41:38:@6114.4]
  assign _T_16349 = select_6 == 5'h7; // @[Switch.scala 41:52:@6116.4]
  assign output_7_6 = io_outValid_6 & _T_16349; // @[Switch.scala 41:38:@6117.4]
  assign _T_16352 = select_7 == 5'h7; // @[Switch.scala 41:52:@6119.4]
  assign output_7_7 = io_outValid_7 & _T_16352; // @[Switch.scala 41:38:@6120.4]
  assign _T_16355 = select_8 == 5'h7; // @[Switch.scala 41:52:@6122.4]
  assign output_7_8 = io_outValid_8 & _T_16355; // @[Switch.scala 41:38:@6123.4]
  assign _T_16358 = select_9 == 5'h7; // @[Switch.scala 41:52:@6125.4]
  assign output_7_9 = io_outValid_9 & _T_16358; // @[Switch.scala 41:38:@6126.4]
  assign _T_16361 = select_10 == 5'h7; // @[Switch.scala 41:52:@6128.4]
  assign output_7_10 = io_outValid_10 & _T_16361; // @[Switch.scala 41:38:@6129.4]
  assign _T_16364 = select_11 == 5'h7; // @[Switch.scala 41:52:@6131.4]
  assign output_7_11 = io_outValid_11 & _T_16364; // @[Switch.scala 41:38:@6132.4]
  assign _T_16367 = select_12 == 5'h7; // @[Switch.scala 41:52:@6134.4]
  assign output_7_12 = io_outValid_12 & _T_16367; // @[Switch.scala 41:38:@6135.4]
  assign _T_16370 = select_13 == 5'h7; // @[Switch.scala 41:52:@6137.4]
  assign output_7_13 = io_outValid_13 & _T_16370; // @[Switch.scala 41:38:@6138.4]
  assign _T_16373 = select_14 == 5'h7; // @[Switch.scala 41:52:@6140.4]
  assign output_7_14 = io_outValid_14 & _T_16373; // @[Switch.scala 41:38:@6141.4]
  assign _T_16376 = select_15 == 5'h7; // @[Switch.scala 41:52:@6143.4]
  assign output_7_15 = io_outValid_15 & _T_16376; // @[Switch.scala 41:38:@6144.4]
  assign _T_16379 = select_16 == 5'h7; // @[Switch.scala 41:52:@6146.4]
  assign output_7_16 = io_outValid_16 & _T_16379; // @[Switch.scala 41:38:@6147.4]
  assign _T_16382 = select_17 == 5'h7; // @[Switch.scala 41:52:@6149.4]
  assign output_7_17 = io_outValid_17 & _T_16382; // @[Switch.scala 41:38:@6150.4]
  assign _T_16385 = select_18 == 5'h7; // @[Switch.scala 41:52:@6152.4]
  assign output_7_18 = io_outValid_18 & _T_16385; // @[Switch.scala 41:38:@6153.4]
  assign _T_16388 = select_19 == 5'h7; // @[Switch.scala 41:52:@6155.4]
  assign output_7_19 = io_outValid_19 & _T_16388; // @[Switch.scala 41:38:@6156.4]
  assign _T_16391 = select_20 == 5'h7; // @[Switch.scala 41:52:@6158.4]
  assign output_7_20 = io_outValid_20 & _T_16391; // @[Switch.scala 41:38:@6159.4]
  assign _T_16394 = select_21 == 5'h7; // @[Switch.scala 41:52:@6161.4]
  assign output_7_21 = io_outValid_21 & _T_16394; // @[Switch.scala 41:38:@6162.4]
  assign _T_16397 = select_22 == 5'h7; // @[Switch.scala 41:52:@6164.4]
  assign output_7_22 = io_outValid_22 & _T_16397; // @[Switch.scala 41:38:@6165.4]
  assign _T_16400 = select_23 == 5'h7; // @[Switch.scala 41:52:@6167.4]
  assign output_7_23 = io_outValid_23 & _T_16400; // @[Switch.scala 41:38:@6168.4]
  assign _T_16403 = select_24 == 5'h7; // @[Switch.scala 41:52:@6170.4]
  assign output_7_24 = io_outValid_24 & _T_16403; // @[Switch.scala 41:38:@6171.4]
  assign _T_16406 = select_25 == 5'h7; // @[Switch.scala 41:52:@6173.4]
  assign output_7_25 = io_outValid_25 & _T_16406; // @[Switch.scala 41:38:@6174.4]
  assign _T_16409 = select_26 == 5'h7; // @[Switch.scala 41:52:@6176.4]
  assign output_7_26 = io_outValid_26 & _T_16409; // @[Switch.scala 41:38:@6177.4]
  assign _T_16412 = select_27 == 5'h7; // @[Switch.scala 41:52:@6179.4]
  assign output_7_27 = io_outValid_27 & _T_16412; // @[Switch.scala 41:38:@6180.4]
  assign _T_16415 = select_28 == 5'h7; // @[Switch.scala 41:52:@6182.4]
  assign output_7_28 = io_outValid_28 & _T_16415; // @[Switch.scala 41:38:@6183.4]
  assign _T_16418 = select_29 == 5'h7; // @[Switch.scala 41:52:@6185.4]
  assign output_7_29 = io_outValid_29 & _T_16418; // @[Switch.scala 41:38:@6186.4]
  assign _T_16421 = select_30 == 5'h7; // @[Switch.scala 41:52:@6188.4]
  assign output_7_30 = io_outValid_30 & _T_16421; // @[Switch.scala 41:38:@6189.4]
  assign _T_16424 = select_31 == 5'h7; // @[Switch.scala 41:52:@6191.4]
  assign output_7_31 = io_outValid_31 & _T_16424; // @[Switch.scala 41:38:@6192.4]
  assign _T_16432 = {output_7_7,output_7_6,output_7_5,output_7_4,output_7_3,output_7_2,output_7_1,output_7_0}; // @[Switch.scala 43:31:@6200.4]
  assign _T_16440 = {output_7_15,output_7_14,output_7_13,output_7_12,output_7_11,output_7_10,output_7_9,output_7_8,_T_16432}; // @[Switch.scala 43:31:@6208.4]
  assign _T_16447 = {output_7_23,output_7_22,output_7_21,output_7_20,output_7_19,output_7_18,output_7_17,output_7_16}; // @[Switch.scala 43:31:@6215.4]
  assign _T_16456 = {output_7_31,output_7_30,output_7_29,output_7_28,output_7_27,output_7_26,output_7_25,output_7_24,_T_16447,_T_16440}; // @[Switch.scala 43:31:@6224.4]
  assign _T_16460 = select_0 == 5'h8; // @[Switch.scala 41:52:@6227.4]
  assign output_8_0 = io_outValid_0 & _T_16460; // @[Switch.scala 41:38:@6228.4]
  assign _T_16463 = select_1 == 5'h8; // @[Switch.scala 41:52:@6230.4]
  assign output_8_1 = io_outValid_1 & _T_16463; // @[Switch.scala 41:38:@6231.4]
  assign _T_16466 = select_2 == 5'h8; // @[Switch.scala 41:52:@6233.4]
  assign output_8_2 = io_outValid_2 & _T_16466; // @[Switch.scala 41:38:@6234.4]
  assign _T_16469 = select_3 == 5'h8; // @[Switch.scala 41:52:@6236.4]
  assign output_8_3 = io_outValid_3 & _T_16469; // @[Switch.scala 41:38:@6237.4]
  assign _T_16472 = select_4 == 5'h8; // @[Switch.scala 41:52:@6239.4]
  assign output_8_4 = io_outValid_4 & _T_16472; // @[Switch.scala 41:38:@6240.4]
  assign _T_16475 = select_5 == 5'h8; // @[Switch.scala 41:52:@6242.4]
  assign output_8_5 = io_outValid_5 & _T_16475; // @[Switch.scala 41:38:@6243.4]
  assign _T_16478 = select_6 == 5'h8; // @[Switch.scala 41:52:@6245.4]
  assign output_8_6 = io_outValid_6 & _T_16478; // @[Switch.scala 41:38:@6246.4]
  assign _T_16481 = select_7 == 5'h8; // @[Switch.scala 41:52:@6248.4]
  assign output_8_7 = io_outValid_7 & _T_16481; // @[Switch.scala 41:38:@6249.4]
  assign _T_16484 = select_8 == 5'h8; // @[Switch.scala 41:52:@6251.4]
  assign output_8_8 = io_outValid_8 & _T_16484; // @[Switch.scala 41:38:@6252.4]
  assign _T_16487 = select_9 == 5'h8; // @[Switch.scala 41:52:@6254.4]
  assign output_8_9 = io_outValid_9 & _T_16487; // @[Switch.scala 41:38:@6255.4]
  assign _T_16490 = select_10 == 5'h8; // @[Switch.scala 41:52:@6257.4]
  assign output_8_10 = io_outValid_10 & _T_16490; // @[Switch.scala 41:38:@6258.4]
  assign _T_16493 = select_11 == 5'h8; // @[Switch.scala 41:52:@6260.4]
  assign output_8_11 = io_outValid_11 & _T_16493; // @[Switch.scala 41:38:@6261.4]
  assign _T_16496 = select_12 == 5'h8; // @[Switch.scala 41:52:@6263.4]
  assign output_8_12 = io_outValid_12 & _T_16496; // @[Switch.scala 41:38:@6264.4]
  assign _T_16499 = select_13 == 5'h8; // @[Switch.scala 41:52:@6266.4]
  assign output_8_13 = io_outValid_13 & _T_16499; // @[Switch.scala 41:38:@6267.4]
  assign _T_16502 = select_14 == 5'h8; // @[Switch.scala 41:52:@6269.4]
  assign output_8_14 = io_outValid_14 & _T_16502; // @[Switch.scala 41:38:@6270.4]
  assign _T_16505 = select_15 == 5'h8; // @[Switch.scala 41:52:@6272.4]
  assign output_8_15 = io_outValid_15 & _T_16505; // @[Switch.scala 41:38:@6273.4]
  assign _T_16508 = select_16 == 5'h8; // @[Switch.scala 41:52:@6275.4]
  assign output_8_16 = io_outValid_16 & _T_16508; // @[Switch.scala 41:38:@6276.4]
  assign _T_16511 = select_17 == 5'h8; // @[Switch.scala 41:52:@6278.4]
  assign output_8_17 = io_outValid_17 & _T_16511; // @[Switch.scala 41:38:@6279.4]
  assign _T_16514 = select_18 == 5'h8; // @[Switch.scala 41:52:@6281.4]
  assign output_8_18 = io_outValid_18 & _T_16514; // @[Switch.scala 41:38:@6282.4]
  assign _T_16517 = select_19 == 5'h8; // @[Switch.scala 41:52:@6284.4]
  assign output_8_19 = io_outValid_19 & _T_16517; // @[Switch.scala 41:38:@6285.4]
  assign _T_16520 = select_20 == 5'h8; // @[Switch.scala 41:52:@6287.4]
  assign output_8_20 = io_outValid_20 & _T_16520; // @[Switch.scala 41:38:@6288.4]
  assign _T_16523 = select_21 == 5'h8; // @[Switch.scala 41:52:@6290.4]
  assign output_8_21 = io_outValid_21 & _T_16523; // @[Switch.scala 41:38:@6291.4]
  assign _T_16526 = select_22 == 5'h8; // @[Switch.scala 41:52:@6293.4]
  assign output_8_22 = io_outValid_22 & _T_16526; // @[Switch.scala 41:38:@6294.4]
  assign _T_16529 = select_23 == 5'h8; // @[Switch.scala 41:52:@6296.4]
  assign output_8_23 = io_outValid_23 & _T_16529; // @[Switch.scala 41:38:@6297.4]
  assign _T_16532 = select_24 == 5'h8; // @[Switch.scala 41:52:@6299.4]
  assign output_8_24 = io_outValid_24 & _T_16532; // @[Switch.scala 41:38:@6300.4]
  assign _T_16535 = select_25 == 5'h8; // @[Switch.scala 41:52:@6302.4]
  assign output_8_25 = io_outValid_25 & _T_16535; // @[Switch.scala 41:38:@6303.4]
  assign _T_16538 = select_26 == 5'h8; // @[Switch.scala 41:52:@6305.4]
  assign output_8_26 = io_outValid_26 & _T_16538; // @[Switch.scala 41:38:@6306.4]
  assign _T_16541 = select_27 == 5'h8; // @[Switch.scala 41:52:@6308.4]
  assign output_8_27 = io_outValid_27 & _T_16541; // @[Switch.scala 41:38:@6309.4]
  assign _T_16544 = select_28 == 5'h8; // @[Switch.scala 41:52:@6311.4]
  assign output_8_28 = io_outValid_28 & _T_16544; // @[Switch.scala 41:38:@6312.4]
  assign _T_16547 = select_29 == 5'h8; // @[Switch.scala 41:52:@6314.4]
  assign output_8_29 = io_outValid_29 & _T_16547; // @[Switch.scala 41:38:@6315.4]
  assign _T_16550 = select_30 == 5'h8; // @[Switch.scala 41:52:@6317.4]
  assign output_8_30 = io_outValid_30 & _T_16550; // @[Switch.scala 41:38:@6318.4]
  assign _T_16553 = select_31 == 5'h8; // @[Switch.scala 41:52:@6320.4]
  assign output_8_31 = io_outValid_31 & _T_16553; // @[Switch.scala 41:38:@6321.4]
  assign _T_16561 = {output_8_7,output_8_6,output_8_5,output_8_4,output_8_3,output_8_2,output_8_1,output_8_0}; // @[Switch.scala 43:31:@6329.4]
  assign _T_16569 = {output_8_15,output_8_14,output_8_13,output_8_12,output_8_11,output_8_10,output_8_9,output_8_8,_T_16561}; // @[Switch.scala 43:31:@6337.4]
  assign _T_16576 = {output_8_23,output_8_22,output_8_21,output_8_20,output_8_19,output_8_18,output_8_17,output_8_16}; // @[Switch.scala 43:31:@6344.4]
  assign _T_16585 = {output_8_31,output_8_30,output_8_29,output_8_28,output_8_27,output_8_26,output_8_25,output_8_24,_T_16576,_T_16569}; // @[Switch.scala 43:31:@6353.4]
  assign _T_16589 = select_0 == 5'h9; // @[Switch.scala 41:52:@6356.4]
  assign output_9_0 = io_outValid_0 & _T_16589; // @[Switch.scala 41:38:@6357.4]
  assign _T_16592 = select_1 == 5'h9; // @[Switch.scala 41:52:@6359.4]
  assign output_9_1 = io_outValid_1 & _T_16592; // @[Switch.scala 41:38:@6360.4]
  assign _T_16595 = select_2 == 5'h9; // @[Switch.scala 41:52:@6362.4]
  assign output_9_2 = io_outValid_2 & _T_16595; // @[Switch.scala 41:38:@6363.4]
  assign _T_16598 = select_3 == 5'h9; // @[Switch.scala 41:52:@6365.4]
  assign output_9_3 = io_outValid_3 & _T_16598; // @[Switch.scala 41:38:@6366.4]
  assign _T_16601 = select_4 == 5'h9; // @[Switch.scala 41:52:@6368.4]
  assign output_9_4 = io_outValid_4 & _T_16601; // @[Switch.scala 41:38:@6369.4]
  assign _T_16604 = select_5 == 5'h9; // @[Switch.scala 41:52:@6371.4]
  assign output_9_5 = io_outValid_5 & _T_16604; // @[Switch.scala 41:38:@6372.4]
  assign _T_16607 = select_6 == 5'h9; // @[Switch.scala 41:52:@6374.4]
  assign output_9_6 = io_outValid_6 & _T_16607; // @[Switch.scala 41:38:@6375.4]
  assign _T_16610 = select_7 == 5'h9; // @[Switch.scala 41:52:@6377.4]
  assign output_9_7 = io_outValid_7 & _T_16610; // @[Switch.scala 41:38:@6378.4]
  assign _T_16613 = select_8 == 5'h9; // @[Switch.scala 41:52:@6380.4]
  assign output_9_8 = io_outValid_8 & _T_16613; // @[Switch.scala 41:38:@6381.4]
  assign _T_16616 = select_9 == 5'h9; // @[Switch.scala 41:52:@6383.4]
  assign output_9_9 = io_outValid_9 & _T_16616; // @[Switch.scala 41:38:@6384.4]
  assign _T_16619 = select_10 == 5'h9; // @[Switch.scala 41:52:@6386.4]
  assign output_9_10 = io_outValid_10 & _T_16619; // @[Switch.scala 41:38:@6387.4]
  assign _T_16622 = select_11 == 5'h9; // @[Switch.scala 41:52:@6389.4]
  assign output_9_11 = io_outValid_11 & _T_16622; // @[Switch.scala 41:38:@6390.4]
  assign _T_16625 = select_12 == 5'h9; // @[Switch.scala 41:52:@6392.4]
  assign output_9_12 = io_outValid_12 & _T_16625; // @[Switch.scala 41:38:@6393.4]
  assign _T_16628 = select_13 == 5'h9; // @[Switch.scala 41:52:@6395.4]
  assign output_9_13 = io_outValid_13 & _T_16628; // @[Switch.scala 41:38:@6396.4]
  assign _T_16631 = select_14 == 5'h9; // @[Switch.scala 41:52:@6398.4]
  assign output_9_14 = io_outValid_14 & _T_16631; // @[Switch.scala 41:38:@6399.4]
  assign _T_16634 = select_15 == 5'h9; // @[Switch.scala 41:52:@6401.4]
  assign output_9_15 = io_outValid_15 & _T_16634; // @[Switch.scala 41:38:@6402.4]
  assign _T_16637 = select_16 == 5'h9; // @[Switch.scala 41:52:@6404.4]
  assign output_9_16 = io_outValid_16 & _T_16637; // @[Switch.scala 41:38:@6405.4]
  assign _T_16640 = select_17 == 5'h9; // @[Switch.scala 41:52:@6407.4]
  assign output_9_17 = io_outValid_17 & _T_16640; // @[Switch.scala 41:38:@6408.4]
  assign _T_16643 = select_18 == 5'h9; // @[Switch.scala 41:52:@6410.4]
  assign output_9_18 = io_outValid_18 & _T_16643; // @[Switch.scala 41:38:@6411.4]
  assign _T_16646 = select_19 == 5'h9; // @[Switch.scala 41:52:@6413.4]
  assign output_9_19 = io_outValid_19 & _T_16646; // @[Switch.scala 41:38:@6414.4]
  assign _T_16649 = select_20 == 5'h9; // @[Switch.scala 41:52:@6416.4]
  assign output_9_20 = io_outValid_20 & _T_16649; // @[Switch.scala 41:38:@6417.4]
  assign _T_16652 = select_21 == 5'h9; // @[Switch.scala 41:52:@6419.4]
  assign output_9_21 = io_outValid_21 & _T_16652; // @[Switch.scala 41:38:@6420.4]
  assign _T_16655 = select_22 == 5'h9; // @[Switch.scala 41:52:@6422.4]
  assign output_9_22 = io_outValid_22 & _T_16655; // @[Switch.scala 41:38:@6423.4]
  assign _T_16658 = select_23 == 5'h9; // @[Switch.scala 41:52:@6425.4]
  assign output_9_23 = io_outValid_23 & _T_16658; // @[Switch.scala 41:38:@6426.4]
  assign _T_16661 = select_24 == 5'h9; // @[Switch.scala 41:52:@6428.4]
  assign output_9_24 = io_outValid_24 & _T_16661; // @[Switch.scala 41:38:@6429.4]
  assign _T_16664 = select_25 == 5'h9; // @[Switch.scala 41:52:@6431.4]
  assign output_9_25 = io_outValid_25 & _T_16664; // @[Switch.scala 41:38:@6432.4]
  assign _T_16667 = select_26 == 5'h9; // @[Switch.scala 41:52:@6434.4]
  assign output_9_26 = io_outValid_26 & _T_16667; // @[Switch.scala 41:38:@6435.4]
  assign _T_16670 = select_27 == 5'h9; // @[Switch.scala 41:52:@6437.4]
  assign output_9_27 = io_outValid_27 & _T_16670; // @[Switch.scala 41:38:@6438.4]
  assign _T_16673 = select_28 == 5'h9; // @[Switch.scala 41:52:@6440.4]
  assign output_9_28 = io_outValid_28 & _T_16673; // @[Switch.scala 41:38:@6441.4]
  assign _T_16676 = select_29 == 5'h9; // @[Switch.scala 41:52:@6443.4]
  assign output_9_29 = io_outValid_29 & _T_16676; // @[Switch.scala 41:38:@6444.4]
  assign _T_16679 = select_30 == 5'h9; // @[Switch.scala 41:52:@6446.4]
  assign output_9_30 = io_outValid_30 & _T_16679; // @[Switch.scala 41:38:@6447.4]
  assign _T_16682 = select_31 == 5'h9; // @[Switch.scala 41:52:@6449.4]
  assign output_9_31 = io_outValid_31 & _T_16682; // @[Switch.scala 41:38:@6450.4]
  assign _T_16690 = {output_9_7,output_9_6,output_9_5,output_9_4,output_9_3,output_9_2,output_9_1,output_9_0}; // @[Switch.scala 43:31:@6458.4]
  assign _T_16698 = {output_9_15,output_9_14,output_9_13,output_9_12,output_9_11,output_9_10,output_9_9,output_9_8,_T_16690}; // @[Switch.scala 43:31:@6466.4]
  assign _T_16705 = {output_9_23,output_9_22,output_9_21,output_9_20,output_9_19,output_9_18,output_9_17,output_9_16}; // @[Switch.scala 43:31:@6473.4]
  assign _T_16714 = {output_9_31,output_9_30,output_9_29,output_9_28,output_9_27,output_9_26,output_9_25,output_9_24,_T_16705,_T_16698}; // @[Switch.scala 43:31:@6482.4]
  assign _T_16718 = select_0 == 5'ha; // @[Switch.scala 41:52:@6485.4]
  assign output_10_0 = io_outValid_0 & _T_16718; // @[Switch.scala 41:38:@6486.4]
  assign _T_16721 = select_1 == 5'ha; // @[Switch.scala 41:52:@6488.4]
  assign output_10_1 = io_outValid_1 & _T_16721; // @[Switch.scala 41:38:@6489.4]
  assign _T_16724 = select_2 == 5'ha; // @[Switch.scala 41:52:@6491.4]
  assign output_10_2 = io_outValid_2 & _T_16724; // @[Switch.scala 41:38:@6492.4]
  assign _T_16727 = select_3 == 5'ha; // @[Switch.scala 41:52:@6494.4]
  assign output_10_3 = io_outValid_3 & _T_16727; // @[Switch.scala 41:38:@6495.4]
  assign _T_16730 = select_4 == 5'ha; // @[Switch.scala 41:52:@6497.4]
  assign output_10_4 = io_outValid_4 & _T_16730; // @[Switch.scala 41:38:@6498.4]
  assign _T_16733 = select_5 == 5'ha; // @[Switch.scala 41:52:@6500.4]
  assign output_10_5 = io_outValid_5 & _T_16733; // @[Switch.scala 41:38:@6501.4]
  assign _T_16736 = select_6 == 5'ha; // @[Switch.scala 41:52:@6503.4]
  assign output_10_6 = io_outValid_6 & _T_16736; // @[Switch.scala 41:38:@6504.4]
  assign _T_16739 = select_7 == 5'ha; // @[Switch.scala 41:52:@6506.4]
  assign output_10_7 = io_outValid_7 & _T_16739; // @[Switch.scala 41:38:@6507.4]
  assign _T_16742 = select_8 == 5'ha; // @[Switch.scala 41:52:@6509.4]
  assign output_10_8 = io_outValid_8 & _T_16742; // @[Switch.scala 41:38:@6510.4]
  assign _T_16745 = select_9 == 5'ha; // @[Switch.scala 41:52:@6512.4]
  assign output_10_9 = io_outValid_9 & _T_16745; // @[Switch.scala 41:38:@6513.4]
  assign _T_16748 = select_10 == 5'ha; // @[Switch.scala 41:52:@6515.4]
  assign output_10_10 = io_outValid_10 & _T_16748; // @[Switch.scala 41:38:@6516.4]
  assign _T_16751 = select_11 == 5'ha; // @[Switch.scala 41:52:@6518.4]
  assign output_10_11 = io_outValid_11 & _T_16751; // @[Switch.scala 41:38:@6519.4]
  assign _T_16754 = select_12 == 5'ha; // @[Switch.scala 41:52:@6521.4]
  assign output_10_12 = io_outValid_12 & _T_16754; // @[Switch.scala 41:38:@6522.4]
  assign _T_16757 = select_13 == 5'ha; // @[Switch.scala 41:52:@6524.4]
  assign output_10_13 = io_outValid_13 & _T_16757; // @[Switch.scala 41:38:@6525.4]
  assign _T_16760 = select_14 == 5'ha; // @[Switch.scala 41:52:@6527.4]
  assign output_10_14 = io_outValid_14 & _T_16760; // @[Switch.scala 41:38:@6528.4]
  assign _T_16763 = select_15 == 5'ha; // @[Switch.scala 41:52:@6530.4]
  assign output_10_15 = io_outValid_15 & _T_16763; // @[Switch.scala 41:38:@6531.4]
  assign _T_16766 = select_16 == 5'ha; // @[Switch.scala 41:52:@6533.4]
  assign output_10_16 = io_outValid_16 & _T_16766; // @[Switch.scala 41:38:@6534.4]
  assign _T_16769 = select_17 == 5'ha; // @[Switch.scala 41:52:@6536.4]
  assign output_10_17 = io_outValid_17 & _T_16769; // @[Switch.scala 41:38:@6537.4]
  assign _T_16772 = select_18 == 5'ha; // @[Switch.scala 41:52:@6539.4]
  assign output_10_18 = io_outValid_18 & _T_16772; // @[Switch.scala 41:38:@6540.4]
  assign _T_16775 = select_19 == 5'ha; // @[Switch.scala 41:52:@6542.4]
  assign output_10_19 = io_outValid_19 & _T_16775; // @[Switch.scala 41:38:@6543.4]
  assign _T_16778 = select_20 == 5'ha; // @[Switch.scala 41:52:@6545.4]
  assign output_10_20 = io_outValid_20 & _T_16778; // @[Switch.scala 41:38:@6546.4]
  assign _T_16781 = select_21 == 5'ha; // @[Switch.scala 41:52:@6548.4]
  assign output_10_21 = io_outValid_21 & _T_16781; // @[Switch.scala 41:38:@6549.4]
  assign _T_16784 = select_22 == 5'ha; // @[Switch.scala 41:52:@6551.4]
  assign output_10_22 = io_outValid_22 & _T_16784; // @[Switch.scala 41:38:@6552.4]
  assign _T_16787 = select_23 == 5'ha; // @[Switch.scala 41:52:@6554.4]
  assign output_10_23 = io_outValid_23 & _T_16787; // @[Switch.scala 41:38:@6555.4]
  assign _T_16790 = select_24 == 5'ha; // @[Switch.scala 41:52:@6557.4]
  assign output_10_24 = io_outValid_24 & _T_16790; // @[Switch.scala 41:38:@6558.4]
  assign _T_16793 = select_25 == 5'ha; // @[Switch.scala 41:52:@6560.4]
  assign output_10_25 = io_outValid_25 & _T_16793; // @[Switch.scala 41:38:@6561.4]
  assign _T_16796 = select_26 == 5'ha; // @[Switch.scala 41:52:@6563.4]
  assign output_10_26 = io_outValid_26 & _T_16796; // @[Switch.scala 41:38:@6564.4]
  assign _T_16799 = select_27 == 5'ha; // @[Switch.scala 41:52:@6566.4]
  assign output_10_27 = io_outValid_27 & _T_16799; // @[Switch.scala 41:38:@6567.4]
  assign _T_16802 = select_28 == 5'ha; // @[Switch.scala 41:52:@6569.4]
  assign output_10_28 = io_outValid_28 & _T_16802; // @[Switch.scala 41:38:@6570.4]
  assign _T_16805 = select_29 == 5'ha; // @[Switch.scala 41:52:@6572.4]
  assign output_10_29 = io_outValid_29 & _T_16805; // @[Switch.scala 41:38:@6573.4]
  assign _T_16808 = select_30 == 5'ha; // @[Switch.scala 41:52:@6575.4]
  assign output_10_30 = io_outValid_30 & _T_16808; // @[Switch.scala 41:38:@6576.4]
  assign _T_16811 = select_31 == 5'ha; // @[Switch.scala 41:52:@6578.4]
  assign output_10_31 = io_outValid_31 & _T_16811; // @[Switch.scala 41:38:@6579.4]
  assign _T_16819 = {output_10_7,output_10_6,output_10_5,output_10_4,output_10_3,output_10_2,output_10_1,output_10_0}; // @[Switch.scala 43:31:@6587.4]
  assign _T_16827 = {output_10_15,output_10_14,output_10_13,output_10_12,output_10_11,output_10_10,output_10_9,output_10_8,_T_16819}; // @[Switch.scala 43:31:@6595.4]
  assign _T_16834 = {output_10_23,output_10_22,output_10_21,output_10_20,output_10_19,output_10_18,output_10_17,output_10_16}; // @[Switch.scala 43:31:@6602.4]
  assign _T_16843 = {output_10_31,output_10_30,output_10_29,output_10_28,output_10_27,output_10_26,output_10_25,output_10_24,_T_16834,_T_16827}; // @[Switch.scala 43:31:@6611.4]
  assign _T_16847 = select_0 == 5'hb; // @[Switch.scala 41:52:@6614.4]
  assign output_11_0 = io_outValid_0 & _T_16847; // @[Switch.scala 41:38:@6615.4]
  assign _T_16850 = select_1 == 5'hb; // @[Switch.scala 41:52:@6617.4]
  assign output_11_1 = io_outValid_1 & _T_16850; // @[Switch.scala 41:38:@6618.4]
  assign _T_16853 = select_2 == 5'hb; // @[Switch.scala 41:52:@6620.4]
  assign output_11_2 = io_outValid_2 & _T_16853; // @[Switch.scala 41:38:@6621.4]
  assign _T_16856 = select_3 == 5'hb; // @[Switch.scala 41:52:@6623.4]
  assign output_11_3 = io_outValid_3 & _T_16856; // @[Switch.scala 41:38:@6624.4]
  assign _T_16859 = select_4 == 5'hb; // @[Switch.scala 41:52:@6626.4]
  assign output_11_4 = io_outValid_4 & _T_16859; // @[Switch.scala 41:38:@6627.4]
  assign _T_16862 = select_5 == 5'hb; // @[Switch.scala 41:52:@6629.4]
  assign output_11_5 = io_outValid_5 & _T_16862; // @[Switch.scala 41:38:@6630.4]
  assign _T_16865 = select_6 == 5'hb; // @[Switch.scala 41:52:@6632.4]
  assign output_11_6 = io_outValid_6 & _T_16865; // @[Switch.scala 41:38:@6633.4]
  assign _T_16868 = select_7 == 5'hb; // @[Switch.scala 41:52:@6635.4]
  assign output_11_7 = io_outValid_7 & _T_16868; // @[Switch.scala 41:38:@6636.4]
  assign _T_16871 = select_8 == 5'hb; // @[Switch.scala 41:52:@6638.4]
  assign output_11_8 = io_outValid_8 & _T_16871; // @[Switch.scala 41:38:@6639.4]
  assign _T_16874 = select_9 == 5'hb; // @[Switch.scala 41:52:@6641.4]
  assign output_11_9 = io_outValid_9 & _T_16874; // @[Switch.scala 41:38:@6642.4]
  assign _T_16877 = select_10 == 5'hb; // @[Switch.scala 41:52:@6644.4]
  assign output_11_10 = io_outValid_10 & _T_16877; // @[Switch.scala 41:38:@6645.4]
  assign _T_16880 = select_11 == 5'hb; // @[Switch.scala 41:52:@6647.4]
  assign output_11_11 = io_outValid_11 & _T_16880; // @[Switch.scala 41:38:@6648.4]
  assign _T_16883 = select_12 == 5'hb; // @[Switch.scala 41:52:@6650.4]
  assign output_11_12 = io_outValid_12 & _T_16883; // @[Switch.scala 41:38:@6651.4]
  assign _T_16886 = select_13 == 5'hb; // @[Switch.scala 41:52:@6653.4]
  assign output_11_13 = io_outValid_13 & _T_16886; // @[Switch.scala 41:38:@6654.4]
  assign _T_16889 = select_14 == 5'hb; // @[Switch.scala 41:52:@6656.4]
  assign output_11_14 = io_outValid_14 & _T_16889; // @[Switch.scala 41:38:@6657.4]
  assign _T_16892 = select_15 == 5'hb; // @[Switch.scala 41:52:@6659.4]
  assign output_11_15 = io_outValid_15 & _T_16892; // @[Switch.scala 41:38:@6660.4]
  assign _T_16895 = select_16 == 5'hb; // @[Switch.scala 41:52:@6662.4]
  assign output_11_16 = io_outValid_16 & _T_16895; // @[Switch.scala 41:38:@6663.4]
  assign _T_16898 = select_17 == 5'hb; // @[Switch.scala 41:52:@6665.4]
  assign output_11_17 = io_outValid_17 & _T_16898; // @[Switch.scala 41:38:@6666.4]
  assign _T_16901 = select_18 == 5'hb; // @[Switch.scala 41:52:@6668.4]
  assign output_11_18 = io_outValid_18 & _T_16901; // @[Switch.scala 41:38:@6669.4]
  assign _T_16904 = select_19 == 5'hb; // @[Switch.scala 41:52:@6671.4]
  assign output_11_19 = io_outValid_19 & _T_16904; // @[Switch.scala 41:38:@6672.4]
  assign _T_16907 = select_20 == 5'hb; // @[Switch.scala 41:52:@6674.4]
  assign output_11_20 = io_outValid_20 & _T_16907; // @[Switch.scala 41:38:@6675.4]
  assign _T_16910 = select_21 == 5'hb; // @[Switch.scala 41:52:@6677.4]
  assign output_11_21 = io_outValid_21 & _T_16910; // @[Switch.scala 41:38:@6678.4]
  assign _T_16913 = select_22 == 5'hb; // @[Switch.scala 41:52:@6680.4]
  assign output_11_22 = io_outValid_22 & _T_16913; // @[Switch.scala 41:38:@6681.4]
  assign _T_16916 = select_23 == 5'hb; // @[Switch.scala 41:52:@6683.4]
  assign output_11_23 = io_outValid_23 & _T_16916; // @[Switch.scala 41:38:@6684.4]
  assign _T_16919 = select_24 == 5'hb; // @[Switch.scala 41:52:@6686.4]
  assign output_11_24 = io_outValid_24 & _T_16919; // @[Switch.scala 41:38:@6687.4]
  assign _T_16922 = select_25 == 5'hb; // @[Switch.scala 41:52:@6689.4]
  assign output_11_25 = io_outValid_25 & _T_16922; // @[Switch.scala 41:38:@6690.4]
  assign _T_16925 = select_26 == 5'hb; // @[Switch.scala 41:52:@6692.4]
  assign output_11_26 = io_outValid_26 & _T_16925; // @[Switch.scala 41:38:@6693.4]
  assign _T_16928 = select_27 == 5'hb; // @[Switch.scala 41:52:@6695.4]
  assign output_11_27 = io_outValid_27 & _T_16928; // @[Switch.scala 41:38:@6696.4]
  assign _T_16931 = select_28 == 5'hb; // @[Switch.scala 41:52:@6698.4]
  assign output_11_28 = io_outValid_28 & _T_16931; // @[Switch.scala 41:38:@6699.4]
  assign _T_16934 = select_29 == 5'hb; // @[Switch.scala 41:52:@6701.4]
  assign output_11_29 = io_outValid_29 & _T_16934; // @[Switch.scala 41:38:@6702.4]
  assign _T_16937 = select_30 == 5'hb; // @[Switch.scala 41:52:@6704.4]
  assign output_11_30 = io_outValid_30 & _T_16937; // @[Switch.scala 41:38:@6705.4]
  assign _T_16940 = select_31 == 5'hb; // @[Switch.scala 41:52:@6707.4]
  assign output_11_31 = io_outValid_31 & _T_16940; // @[Switch.scala 41:38:@6708.4]
  assign _T_16948 = {output_11_7,output_11_6,output_11_5,output_11_4,output_11_3,output_11_2,output_11_1,output_11_0}; // @[Switch.scala 43:31:@6716.4]
  assign _T_16956 = {output_11_15,output_11_14,output_11_13,output_11_12,output_11_11,output_11_10,output_11_9,output_11_8,_T_16948}; // @[Switch.scala 43:31:@6724.4]
  assign _T_16963 = {output_11_23,output_11_22,output_11_21,output_11_20,output_11_19,output_11_18,output_11_17,output_11_16}; // @[Switch.scala 43:31:@6731.4]
  assign _T_16972 = {output_11_31,output_11_30,output_11_29,output_11_28,output_11_27,output_11_26,output_11_25,output_11_24,_T_16963,_T_16956}; // @[Switch.scala 43:31:@6740.4]
  assign _T_16976 = select_0 == 5'hc; // @[Switch.scala 41:52:@6743.4]
  assign output_12_0 = io_outValid_0 & _T_16976; // @[Switch.scala 41:38:@6744.4]
  assign _T_16979 = select_1 == 5'hc; // @[Switch.scala 41:52:@6746.4]
  assign output_12_1 = io_outValid_1 & _T_16979; // @[Switch.scala 41:38:@6747.4]
  assign _T_16982 = select_2 == 5'hc; // @[Switch.scala 41:52:@6749.4]
  assign output_12_2 = io_outValid_2 & _T_16982; // @[Switch.scala 41:38:@6750.4]
  assign _T_16985 = select_3 == 5'hc; // @[Switch.scala 41:52:@6752.4]
  assign output_12_3 = io_outValid_3 & _T_16985; // @[Switch.scala 41:38:@6753.4]
  assign _T_16988 = select_4 == 5'hc; // @[Switch.scala 41:52:@6755.4]
  assign output_12_4 = io_outValid_4 & _T_16988; // @[Switch.scala 41:38:@6756.4]
  assign _T_16991 = select_5 == 5'hc; // @[Switch.scala 41:52:@6758.4]
  assign output_12_5 = io_outValid_5 & _T_16991; // @[Switch.scala 41:38:@6759.4]
  assign _T_16994 = select_6 == 5'hc; // @[Switch.scala 41:52:@6761.4]
  assign output_12_6 = io_outValid_6 & _T_16994; // @[Switch.scala 41:38:@6762.4]
  assign _T_16997 = select_7 == 5'hc; // @[Switch.scala 41:52:@6764.4]
  assign output_12_7 = io_outValid_7 & _T_16997; // @[Switch.scala 41:38:@6765.4]
  assign _T_17000 = select_8 == 5'hc; // @[Switch.scala 41:52:@6767.4]
  assign output_12_8 = io_outValid_8 & _T_17000; // @[Switch.scala 41:38:@6768.4]
  assign _T_17003 = select_9 == 5'hc; // @[Switch.scala 41:52:@6770.4]
  assign output_12_9 = io_outValid_9 & _T_17003; // @[Switch.scala 41:38:@6771.4]
  assign _T_17006 = select_10 == 5'hc; // @[Switch.scala 41:52:@6773.4]
  assign output_12_10 = io_outValid_10 & _T_17006; // @[Switch.scala 41:38:@6774.4]
  assign _T_17009 = select_11 == 5'hc; // @[Switch.scala 41:52:@6776.4]
  assign output_12_11 = io_outValid_11 & _T_17009; // @[Switch.scala 41:38:@6777.4]
  assign _T_17012 = select_12 == 5'hc; // @[Switch.scala 41:52:@6779.4]
  assign output_12_12 = io_outValid_12 & _T_17012; // @[Switch.scala 41:38:@6780.4]
  assign _T_17015 = select_13 == 5'hc; // @[Switch.scala 41:52:@6782.4]
  assign output_12_13 = io_outValid_13 & _T_17015; // @[Switch.scala 41:38:@6783.4]
  assign _T_17018 = select_14 == 5'hc; // @[Switch.scala 41:52:@6785.4]
  assign output_12_14 = io_outValid_14 & _T_17018; // @[Switch.scala 41:38:@6786.4]
  assign _T_17021 = select_15 == 5'hc; // @[Switch.scala 41:52:@6788.4]
  assign output_12_15 = io_outValid_15 & _T_17021; // @[Switch.scala 41:38:@6789.4]
  assign _T_17024 = select_16 == 5'hc; // @[Switch.scala 41:52:@6791.4]
  assign output_12_16 = io_outValid_16 & _T_17024; // @[Switch.scala 41:38:@6792.4]
  assign _T_17027 = select_17 == 5'hc; // @[Switch.scala 41:52:@6794.4]
  assign output_12_17 = io_outValid_17 & _T_17027; // @[Switch.scala 41:38:@6795.4]
  assign _T_17030 = select_18 == 5'hc; // @[Switch.scala 41:52:@6797.4]
  assign output_12_18 = io_outValid_18 & _T_17030; // @[Switch.scala 41:38:@6798.4]
  assign _T_17033 = select_19 == 5'hc; // @[Switch.scala 41:52:@6800.4]
  assign output_12_19 = io_outValid_19 & _T_17033; // @[Switch.scala 41:38:@6801.4]
  assign _T_17036 = select_20 == 5'hc; // @[Switch.scala 41:52:@6803.4]
  assign output_12_20 = io_outValid_20 & _T_17036; // @[Switch.scala 41:38:@6804.4]
  assign _T_17039 = select_21 == 5'hc; // @[Switch.scala 41:52:@6806.4]
  assign output_12_21 = io_outValid_21 & _T_17039; // @[Switch.scala 41:38:@6807.4]
  assign _T_17042 = select_22 == 5'hc; // @[Switch.scala 41:52:@6809.4]
  assign output_12_22 = io_outValid_22 & _T_17042; // @[Switch.scala 41:38:@6810.4]
  assign _T_17045 = select_23 == 5'hc; // @[Switch.scala 41:52:@6812.4]
  assign output_12_23 = io_outValid_23 & _T_17045; // @[Switch.scala 41:38:@6813.4]
  assign _T_17048 = select_24 == 5'hc; // @[Switch.scala 41:52:@6815.4]
  assign output_12_24 = io_outValid_24 & _T_17048; // @[Switch.scala 41:38:@6816.4]
  assign _T_17051 = select_25 == 5'hc; // @[Switch.scala 41:52:@6818.4]
  assign output_12_25 = io_outValid_25 & _T_17051; // @[Switch.scala 41:38:@6819.4]
  assign _T_17054 = select_26 == 5'hc; // @[Switch.scala 41:52:@6821.4]
  assign output_12_26 = io_outValid_26 & _T_17054; // @[Switch.scala 41:38:@6822.4]
  assign _T_17057 = select_27 == 5'hc; // @[Switch.scala 41:52:@6824.4]
  assign output_12_27 = io_outValid_27 & _T_17057; // @[Switch.scala 41:38:@6825.4]
  assign _T_17060 = select_28 == 5'hc; // @[Switch.scala 41:52:@6827.4]
  assign output_12_28 = io_outValid_28 & _T_17060; // @[Switch.scala 41:38:@6828.4]
  assign _T_17063 = select_29 == 5'hc; // @[Switch.scala 41:52:@6830.4]
  assign output_12_29 = io_outValid_29 & _T_17063; // @[Switch.scala 41:38:@6831.4]
  assign _T_17066 = select_30 == 5'hc; // @[Switch.scala 41:52:@6833.4]
  assign output_12_30 = io_outValid_30 & _T_17066; // @[Switch.scala 41:38:@6834.4]
  assign _T_17069 = select_31 == 5'hc; // @[Switch.scala 41:52:@6836.4]
  assign output_12_31 = io_outValid_31 & _T_17069; // @[Switch.scala 41:38:@6837.4]
  assign _T_17077 = {output_12_7,output_12_6,output_12_5,output_12_4,output_12_3,output_12_2,output_12_1,output_12_0}; // @[Switch.scala 43:31:@6845.4]
  assign _T_17085 = {output_12_15,output_12_14,output_12_13,output_12_12,output_12_11,output_12_10,output_12_9,output_12_8,_T_17077}; // @[Switch.scala 43:31:@6853.4]
  assign _T_17092 = {output_12_23,output_12_22,output_12_21,output_12_20,output_12_19,output_12_18,output_12_17,output_12_16}; // @[Switch.scala 43:31:@6860.4]
  assign _T_17101 = {output_12_31,output_12_30,output_12_29,output_12_28,output_12_27,output_12_26,output_12_25,output_12_24,_T_17092,_T_17085}; // @[Switch.scala 43:31:@6869.4]
  assign _T_17105 = select_0 == 5'hd; // @[Switch.scala 41:52:@6872.4]
  assign output_13_0 = io_outValid_0 & _T_17105; // @[Switch.scala 41:38:@6873.4]
  assign _T_17108 = select_1 == 5'hd; // @[Switch.scala 41:52:@6875.4]
  assign output_13_1 = io_outValid_1 & _T_17108; // @[Switch.scala 41:38:@6876.4]
  assign _T_17111 = select_2 == 5'hd; // @[Switch.scala 41:52:@6878.4]
  assign output_13_2 = io_outValid_2 & _T_17111; // @[Switch.scala 41:38:@6879.4]
  assign _T_17114 = select_3 == 5'hd; // @[Switch.scala 41:52:@6881.4]
  assign output_13_3 = io_outValid_3 & _T_17114; // @[Switch.scala 41:38:@6882.4]
  assign _T_17117 = select_4 == 5'hd; // @[Switch.scala 41:52:@6884.4]
  assign output_13_4 = io_outValid_4 & _T_17117; // @[Switch.scala 41:38:@6885.4]
  assign _T_17120 = select_5 == 5'hd; // @[Switch.scala 41:52:@6887.4]
  assign output_13_5 = io_outValid_5 & _T_17120; // @[Switch.scala 41:38:@6888.4]
  assign _T_17123 = select_6 == 5'hd; // @[Switch.scala 41:52:@6890.4]
  assign output_13_6 = io_outValid_6 & _T_17123; // @[Switch.scala 41:38:@6891.4]
  assign _T_17126 = select_7 == 5'hd; // @[Switch.scala 41:52:@6893.4]
  assign output_13_7 = io_outValid_7 & _T_17126; // @[Switch.scala 41:38:@6894.4]
  assign _T_17129 = select_8 == 5'hd; // @[Switch.scala 41:52:@6896.4]
  assign output_13_8 = io_outValid_8 & _T_17129; // @[Switch.scala 41:38:@6897.4]
  assign _T_17132 = select_9 == 5'hd; // @[Switch.scala 41:52:@6899.4]
  assign output_13_9 = io_outValid_9 & _T_17132; // @[Switch.scala 41:38:@6900.4]
  assign _T_17135 = select_10 == 5'hd; // @[Switch.scala 41:52:@6902.4]
  assign output_13_10 = io_outValid_10 & _T_17135; // @[Switch.scala 41:38:@6903.4]
  assign _T_17138 = select_11 == 5'hd; // @[Switch.scala 41:52:@6905.4]
  assign output_13_11 = io_outValid_11 & _T_17138; // @[Switch.scala 41:38:@6906.4]
  assign _T_17141 = select_12 == 5'hd; // @[Switch.scala 41:52:@6908.4]
  assign output_13_12 = io_outValid_12 & _T_17141; // @[Switch.scala 41:38:@6909.4]
  assign _T_17144 = select_13 == 5'hd; // @[Switch.scala 41:52:@6911.4]
  assign output_13_13 = io_outValid_13 & _T_17144; // @[Switch.scala 41:38:@6912.4]
  assign _T_17147 = select_14 == 5'hd; // @[Switch.scala 41:52:@6914.4]
  assign output_13_14 = io_outValid_14 & _T_17147; // @[Switch.scala 41:38:@6915.4]
  assign _T_17150 = select_15 == 5'hd; // @[Switch.scala 41:52:@6917.4]
  assign output_13_15 = io_outValid_15 & _T_17150; // @[Switch.scala 41:38:@6918.4]
  assign _T_17153 = select_16 == 5'hd; // @[Switch.scala 41:52:@6920.4]
  assign output_13_16 = io_outValid_16 & _T_17153; // @[Switch.scala 41:38:@6921.4]
  assign _T_17156 = select_17 == 5'hd; // @[Switch.scala 41:52:@6923.4]
  assign output_13_17 = io_outValid_17 & _T_17156; // @[Switch.scala 41:38:@6924.4]
  assign _T_17159 = select_18 == 5'hd; // @[Switch.scala 41:52:@6926.4]
  assign output_13_18 = io_outValid_18 & _T_17159; // @[Switch.scala 41:38:@6927.4]
  assign _T_17162 = select_19 == 5'hd; // @[Switch.scala 41:52:@6929.4]
  assign output_13_19 = io_outValid_19 & _T_17162; // @[Switch.scala 41:38:@6930.4]
  assign _T_17165 = select_20 == 5'hd; // @[Switch.scala 41:52:@6932.4]
  assign output_13_20 = io_outValid_20 & _T_17165; // @[Switch.scala 41:38:@6933.4]
  assign _T_17168 = select_21 == 5'hd; // @[Switch.scala 41:52:@6935.4]
  assign output_13_21 = io_outValid_21 & _T_17168; // @[Switch.scala 41:38:@6936.4]
  assign _T_17171 = select_22 == 5'hd; // @[Switch.scala 41:52:@6938.4]
  assign output_13_22 = io_outValid_22 & _T_17171; // @[Switch.scala 41:38:@6939.4]
  assign _T_17174 = select_23 == 5'hd; // @[Switch.scala 41:52:@6941.4]
  assign output_13_23 = io_outValid_23 & _T_17174; // @[Switch.scala 41:38:@6942.4]
  assign _T_17177 = select_24 == 5'hd; // @[Switch.scala 41:52:@6944.4]
  assign output_13_24 = io_outValid_24 & _T_17177; // @[Switch.scala 41:38:@6945.4]
  assign _T_17180 = select_25 == 5'hd; // @[Switch.scala 41:52:@6947.4]
  assign output_13_25 = io_outValid_25 & _T_17180; // @[Switch.scala 41:38:@6948.4]
  assign _T_17183 = select_26 == 5'hd; // @[Switch.scala 41:52:@6950.4]
  assign output_13_26 = io_outValid_26 & _T_17183; // @[Switch.scala 41:38:@6951.4]
  assign _T_17186 = select_27 == 5'hd; // @[Switch.scala 41:52:@6953.4]
  assign output_13_27 = io_outValid_27 & _T_17186; // @[Switch.scala 41:38:@6954.4]
  assign _T_17189 = select_28 == 5'hd; // @[Switch.scala 41:52:@6956.4]
  assign output_13_28 = io_outValid_28 & _T_17189; // @[Switch.scala 41:38:@6957.4]
  assign _T_17192 = select_29 == 5'hd; // @[Switch.scala 41:52:@6959.4]
  assign output_13_29 = io_outValid_29 & _T_17192; // @[Switch.scala 41:38:@6960.4]
  assign _T_17195 = select_30 == 5'hd; // @[Switch.scala 41:52:@6962.4]
  assign output_13_30 = io_outValid_30 & _T_17195; // @[Switch.scala 41:38:@6963.4]
  assign _T_17198 = select_31 == 5'hd; // @[Switch.scala 41:52:@6965.4]
  assign output_13_31 = io_outValid_31 & _T_17198; // @[Switch.scala 41:38:@6966.4]
  assign _T_17206 = {output_13_7,output_13_6,output_13_5,output_13_4,output_13_3,output_13_2,output_13_1,output_13_0}; // @[Switch.scala 43:31:@6974.4]
  assign _T_17214 = {output_13_15,output_13_14,output_13_13,output_13_12,output_13_11,output_13_10,output_13_9,output_13_8,_T_17206}; // @[Switch.scala 43:31:@6982.4]
  assign _T_17221 = {output_13_23,output_13_22,output_13_21,output_13_20,output_13_19,output_13_18,output_13_17,output_13_16}; // @[Switch.scala 43:31:@6989.4]
  assign _T_17230 = {output_13_31,output_13_30,output_13_29,output_13_28,output_13_27,output_13_26,output_13_25,output_13_24,_T_17221,_T_17214}; // @[Switch.scala 43:31:@6998.4]
  assign _T_17234 = select_0 == 5'he; // @[Switch.scala 41:52:@7001.4]
  assign output_14_0 = io_outValid_0 & _T_17234; // @[Switch.scala 41:38:@7002.4]
  assign _T_17237 = select_1 == 5'he; // @[Switch.scala 41:52:@7004.4]
  assign output_14_1 = io_outValid_1 & _T_17237; // @[Switch.scala 41:38:@7005.4]
  assign _T_17240 = select_2 == 5'he; // @[Switch.scala 41:52:@7007.4]
  assign output_14_2 = io_outValid_2 & _T_17240; // @[Switch.scala 41:38:@7008.4]
  assign _T_17243 = select_3 == 5'he; // @[Switch.scala 41:52:@7010.4]
  assign output_14_3 = io_outValid_3 & _T_17243; // @[Switch.scala 41:38:@7011.4]
  assign _T_17246 = select_4 == 5'he; // @[Switch.scala 41:52:@7013.4]
  assign output_14_4 = io_outValid_4 & _T_17246; // @[Switch.scala 41:38:@7014.4]
  assign _T_17249 = select_5 == 5'he; // @[Switch.scala 41:52:@7016.4]
  assign output_14_5 = io_outValid_5 & _T_17249; // @[Switch.scala 41:38:@7017.4]
  assign _T_17252 = select_6 == 5'he; // @[Switch.scala 41:52:@7019.4]
  assign output_14_6 = io_outValid_6 & _T_17252; // @[Switch.scala 41:38:@7020.4]
  assign _T_17255 = select_7 == 5'he; // @[Switch.scala 41:52:@7022.4]
  assign output_14_7 = io_outValid_7 & _T_17255; // @[Switch.scala 41:38:@7023.4]
  assign _T_17258 = select_8 == 5'he; // @[Switch.scala 41:52:@7025.4]
  assign output_14_8 = io_outValid_8 & _T_17258; // @[Switch.scala 41:38:@7026.4]
  assign _T_17261 = select_9 == 5'he; // @[Switch.scala 41:52:@7028.4]
  assign output_14_9 = io_outValid_9 & _T_17261; // @[Switch.scala 41:38:@7029.4]
  assign _T_17264 = select_10 == 5'he; // @[Switch.scala 41:52:@7031.4]
  assign output_14_10 = io_outValid_10 & _T_17264; // @[Switch.scala 41:38:@7032.4]
  assign _T_17267 = select_11 == 5'he; // @[Switch.scala 41:52:@7034.4]
  assign output_14_11 = io_outValid_11 & _T_17267; // @[Switch.scala 41:38:@7035.4]
  assign _T_17270 = select_12 == 5'he; // @[Switch.scala 41:52:@7037.4]
  assign output_14_12 = io_outValid_12 & _T_17270; // @[Switch.scala 41:38:@7038.4]
  assign _T_17273 = select_13 == 5'he; // @[Switch.scala 41:52:@7040.4]
  assign output_14_13 = io_outValid_13 & _T_17273; // @[Switch.scala 41:38:@7041.4]
  assign _T_17276 = select_14 == 5'he; // @[Switch.scala 41:52:@7043.4]
  assign output_14_14 = io_outValid_14 & _T_17276; // @[Switch.scala 41:38:@7044.4]
  assign _T_17279 = select_15 == 5'he; // @[Switch.scala 41:52:@7046.4]
  assign output_14_15 = io_outValid_15 & _T_17279; // @[Switch.scala 41:38:@7047.4]
  assign _T_17282 = select_16 == 5'he; // @[Switch.scala 41:52:@7049.4]
  assign output_14_16 = io_outValid_16 & _T_17282; // @[Switch.scala 41:38:@7050.4]
  assign _T_17285 = select_17 == 5'he; // @[Switch.scala 41:52:@7052.4]
  assign output_14_17 = io_outValid_17 & _T_17285; // @[Switch.scala 41:38:@7053.4]
  assign _T_17288 = select_18 == 5'he; // @[Switch.scala 41:52:@7055.4]
  assign output_14_18 = io_outValid_18 & _T_17288; // @[Switch.scala 41:38:@7056.4]
  assign _T_17291 = select_19 == 5'he; // @[Switch.scala 41:52:@7058.4]
  assign output_14_19 = io_outValid_19 & _T_17291; // @[Switch.scala 41:38:@7059.4]
  assign _T_17294 = select_20 == 5'he; // @[Switch.scala 41:52:@7061.4]
  assign output_14_20 = io_outValid_20 & _T_17294; // @[Switch.scala 41:38:@7062.4]
  assign _T_17297 = select_21 == 5'he; // @[Switch.scala 41:52:@7064.4]
  assign output_14_21 = io_outValid_21 & _T_17297; // @[Switch.scala 41:38:@7065.4]
  assign _T_17300 = select_22 == 5'he; // @[Switch.scala 41:52:@7067.4]
  assign output_14_22 = io_outValid_22 & _T_17300; // @[Switch.scala 41:38:@7068.4]
  assign _T_17303 = select_23 == 5'he; // @[Switch.scala 41:52:@7070.4]
  assign output_14_23 = io_outValid_23 & _T_17303; // @[Switch.scala 41:38:@7071.4]
  assign _T_17306 = select_24 == 5'he; // @[Switch.scala 41:52:@7073.4]
  assign output_14_24 = io_outValid_24 & _T_17306; // @[Switch.scala 41:38:@7074.4]
  assign _T_17309 = select_25 == 5'he; // @[Switch.scala 41:52:@7076.4]
  assign output_14_25 = io_outValid_25 & _T_17309; // @[Switch.scala 41:38:@7077.4]
  assign _T_17312 = select_26 == 5'he; // @[Switch.scala 41:52:@7079.4]
  assign output_14_26 = io_outValid_26 & _T_17312; // @[Switch.scala 41:38:@7080.4]
  assign _T_17315 = select_27 == 5'he; // @[Switch.scala 41:52:@7082.4]
  assign output_14_27 = io_outValid_27 & _T_17315; // @[Switch.scala 41:38:@7083.4]
  assign _T_17318 = select_28 == 5'he; // @[Switch.scala 41:52:@7085.4]
  assign output_14_28 = io_outValid_28 & _T_17318; // @[Switch.scala 41:38:@7086.4]
  assign _T_17321 = select_29 == 5'he; // @[Switch.scala 41:52:@7088.4]
  assign output_14_29 = io_outValid_29 & _T_17321; // @[Switch.scala 41:38:@7089.4]
  assign _T_17324 = select_30 == 5'he; // @[Switch.scala 41:52:@7091.4]
  assign output_14_30 = io_outValid_30 & _T_17324; // @[Switch.scala 41:38:@7092.4]
  assign _T_17327 = select_31 == 5'he; // @[Switch.scala 41:52:@7094.4]
  assign output_14_31 = io_outValid_31 & _T_17327; // @[Switch.scala 41:38:@7095.4]
  assign _T_17335 = {output_14_7,output_14_6,output_14_5,output_14_4,output_14_3,output_14_2,output_14_1,output_14_0}; // @[Switch.scala 43:31:@7103.4]
  assign _T_17343 = {output_14_15,output_14_14,output_14_13,output_14_12,output_14_11,output_14_10,output_14_9,output_14_8,_T_17335}; // @[Switch.scala 43:31:@7111.4]
  assign _T_17350 = {output_14_23,output_14_22,output_14_21,output_14_20,output_14_19,output_14_18,output_14_17,output_14_16}; // @[Switch.scala 43:31:@7118.4]
  assign _T_17359 = {output_14_31,output_14_30,output_14_29,output_14_28,output_14_27,output_14_26,output_14_25,output_14_24,_T_17350,_T_17343}; // @[Switch.scala 43:31:@7127.4]
  assign _T_17363 = select_0 == 5'hf; // @[Switch.scala 41:52:@7130.4]
  assign output_15_0 = io_outValid_0 & _T_17363; // @[Switch.scala 41:38:@7131.4]
  assign _T_17366 = select_1 == 5'hf; // @[Switch.scala 41:52:@7133.4]
  assign output_15_1 = io_outValid_1 & _T_17366; // @[Switch.scala 41:38:@7134.4]
  assign _T_17369 = select_2 == 5'hf; // @[Switch.scala 41:52:@7136.4]
  assign output_15_2 = io_outValid_2 & _T_17369; // @[Switch.scala 41:38:@7137.4]
  assign _T_17372 = select_3 == 5'hf; // @[Switch.scala 41:52:@7139.4]
  assign output_15_3 = io_outValid_3 & _T_17372; // @[Switch.scala 41:38:@7140.4]
  assign _T_17375 = select_4 == 5'hf; // @[Switch.scala 41:52:@7142.4]
  assign output_15_4 = io_outValid_4 & _T_17375; // @[Switch.scala 41:38:@7143.4]
  assign _T_17378 = select_5 == 5'hf; // @[Switch.scala 41:52:@7145.4]
  assign output_15_5 = io_outValid_5 & _T_17378; // @[Switch.scala 41:38:@7146.4]
  assign _T_17381 = select_6 == 5'hf; // @[Switch.scala 41:52:@7148.4]
  assign output_15_6 = io_outValid_6 & _T_17381; // @[Switch.scala 41:38:@7149.4]
  assign _T_17384 = select_7 == 5'hf; // @[Switch.scala 41:52:@7151.4]
  assign output_15_7 = io_outValid_7 & _T_17384; // @[Switch.scala 41:38:@7152.4]
  assign _T_17387 = select_8 == 5'hf; // @[Switch.scala 41:52:@7154.4]
  assign output_15_8 = io_outValid_8 & _T_17387; // @[Switch.scala 41:38:@7155.4]
  assign _T_17390 = select_9 == 5'hf; // @[Switch.scala 41:52:@7157.4]
  assign output_15_9 = io_outValid_9 & _T_17390; // @[Switch.scala 41:38:@7158.4]
  assign _T_17393 = select_10 == 5'hf; // @[Switch.scala 41:52:@7160.4]
  assign output_15_10 = io_outValid_10 & _T_17393; // @[Switch.scala 41:38:@7161.4]
  assign _T_17396 = select_11 == 5'hf; // @[Switch.scala 41:52:@7163.4]
  assign output_15_11 = io_outValid_11 & _T_17396; // @[Switch.scala 41:38:@7164.4]
  assign _T_17399 = select_12 == 5'hf; // @[Switch.scala 41:52:@7166.4]
  assign output_15_12 = io_outValid_12 & _T_17399; // @[Switch.scala 41:38:@7167.4]
  assign _T_17402 = select_13 == 5'hf; // @[Switch.scala 41:52:@7169.4]
  assign output_15_13 = io_outValid_13 & _T_17402; // @[Switch.scala 41:38:@7170.4]
  assign _T_17405 = select_14 == 5'hf; // @[Switch.scala 41:52:@7172.4]
  assign output_15_14 = io_outValid_14 & _T_17405; // @[Switch.scala 41:38:@7173.4]
  assign _T_17408 = select_15 == 5'hf; // @[Switch.scala 41:52:@7175.4]
  assign output_15_15 = io_outValid_15 & _T_17408; // @[Switch.scala 41:38:@7176.4]
  assign _T_17411 = select_16 == 5'hf; // @[Switch.scala 41:52:@7178.4]
  assign output_15_16 = io_outValid_16 & _T_17411; // @[Switch.scala 41:38:@7179.4]
  assign _T_17414 = select_17 == 5'hf; // @[Switch.scala 41:52:@7181.4]
  assign output_15_17 = io_outValid_17 & _T_17414; // @[Switch.scala 41:38:@7182.4]
  assign _T_17417 = select_18 == 5'hf; // @[Switch.scala 41:52:@7184.4]
  assign output_15_18 = io_outValid_18 & _T_17417; // @[Switch.scala 41:38:@7185.4]
  assign _T_17420 = select_19 == 5'hf; // @[Switch.scala 41:52:@7187.4]
  assign output_15_19 = io_outValid_19 & _T_17420; // @[Switch.scala 41:38:@7188.4]
  assign _T_17423 = select_20 == 5'hf; // @[Switch.scala 41:52:@7190.4]
  assign output_15_20 = io_outValid_20 & _T_17423; // @[Switch.scala 41:38:@7191.4]
  assign _T_17426 = select_21 == 5'hf; // @[Switch.scala 41:52:@7193.4]
  assign output_15_21 = io_outValid_21 & _T_17426; // @[Switch.scala 41:38:@7194.4]
  assign _T_17429 = select_22 == 5'hf; // @[Switch.scala 41:52:@7196.4]
  assign output_15_22 = io_outValid_22 & _T_17429; // @[Switch.scala 41:38:@7197.4]
  assign _T_17432 = select_23 == 5'hf; // @[Switch.scala 41:52:@7199.4]
  assign output_15_23 = io_outValid_23 & _T_17432; // @[Switch.scala 41:38:@7200.4]
  assign _T_17435 = select_24 == 5'hf; // @[Switch.scala 41:52:@7202.4]
  assign output_15_24 = io_outValid_24 & _T_17435; // @[Switch.scala 41:38:@7203.4]
  assign _T_17438 = select_25 == 5'hf; // @[Switch.scala 41:52:@7205.4]
  assign output_15_25 = io_outValid_25 & _T_17438; // @[Switch.scala 41:38:@7206.4]
  assign _T_17441 = select_26 == 5'hf; // @[Switch.scala 41:52:@7208.4]
  assign output_15_26 = io_outValid_26 & _T_17441; // @[Switch.scala 41:38:@7209.4]
  assign _T_17444 = select_27 == 5'hf; // @[Switch.scala 41:52:@7211.4]
  assign output_15_27 = io_outValid_27 & _T_17444; // @[Switch.scala 41:38:@7212.4]
  assign _T_17447 = select_28 == 5'hf; // @[Switch.scala 41:52:@7214.4]
  assign output_15_28 = io_outValid_28 & _T_17447; // @[Switch.scala 41:38:@7215.4]
  assign _T_17450 = select_29 == 5'hf; // @[Switch.scala 41:52:@7217.4]
  assign output_15_29 = io_outValid_29 & _T_17450; // @[Switch.scala 41:38:@7218.4]
  assign _T_17453 = select_30 == 5'hf; // @[Switch.scala 41:52:@7220.4]
  assign output_15_30 = io_outValid_30 & _T_17453; // @[Switch.scala 41:38:@7221.4]
  assign _T_17456 = select_31 == 5'hf; // @[Switch.scala 41:52:@7223.4]
  assign output_15_31 = io_outValid_31 & _T_17456; // @[Switch.scala 41:38:@7224.4]
  assign _T_17464 = {output_15_7,output_15_6,output_15_5,output_15_4,output_15_3,output_15_2,output_15_1,output_15_0}; // @[Switch.scala 43:31:@7232.4]
  assign _T_17472 = {output_15_15,output_15_14,output_15_13,output_15_12,output_15_11,output_15_10,output_15_9,output_15_8,_T_17464}; // @[Switch.scala 43:31:@7240.4]
  assign _T_17479 = {output_15_23,output_15_22,output_15_21,output_15_20,output_15_19,output_15_18,output_15_17,output_15_16}; // @[Switch.scala 43:31:@7247.4]
  assign _T_17488 = {output_15_31,output_15_30,output_15_29,output_15_28,output_15_27,output_15_26,output_15_25,output_15_24,_T_17479,_T_17472}; // @[Switch.scala 43:31:@7256.4]
  assign _T_17492 = select_0 == 5'h10; // @[Switch.scala 41:52:@7259.4]
  assign output_16_0 = io_outValid_0 & _T_17492; // @[Switch.scala 41:38:@7260.4]
  assign _T_17495 = select_1 == 5'h10; // @[Switch.scala 41:52:@7262.4]
  assign output_16_1 = io_outValid_1 & _T_17495; // @[Switch.scala 41:38:@7263.4]
  assign _T_17498 = select_2 == 5'h10; // @[Switch.scala 41:52:@7265.4]
  assign output_16_2 = io_outValid_2 & _T_17498; // @[Switch.scala 41:38:@7266.4]
  assign _T_17501 = select_3 == 5'h10; // @[Switch.scala 41:52:@7268.4]
  assign output_16_3 = io_outValid_3 & _T_17501; // @[Switch.scala 41:38:@7269.4]
  assign _T_17504 = select_4 == 5'h10; // @[Switch.scala 41:52:@7271.4]
  assign output_16_4 = io_outValid_4 & _T_17504; // @[Switch.scala 41:38:@7272.4]
  assign _T_17507 = select_5 == 5'h10; // @[Switch.scala 41:52:@7274.4]
  assign output_16_5 = io_outValid_5 & _T_17507; // @[Switch.scala 41:38:@7275.4]
  assign _T_17510 = select_6 == 5'h10; // @[Switch.scala 41:52:@7277.4]
  assign output_16_6 = io_outValid_6 & _T_17510; // @[Switch.scala 41:38:@7278.4]
  assign _T_17513 = select_7 == 5'h10; // @[Switch.scala 41:52:@7280.4]
  assign output_16_7 = io_outValid_7 & _T_17513; // @[Switch.scala 41:38:@7281.4]
  assign _T_17516 = select_8 == 5'h10; // @[Switch.scala 41:52:@7283.4]
  assign output_16_8 = io_outValid_8 & _T_17516; // @[Switch.scala 41:38:@7284.4]
  assign _T_17519 = select_9 == 5'h10; // @[Switch.scala 41:52:@7286.4]
  assign output_16_9 = io_outValid_9 & _T_17519; // @[Switch.scala 41:38:@7287.4]
  assign _T_17522 = select_10 == 5'h10; // @[Switch.scala 41:52:@7289.4]
  assign output_16_10 = io_outValid_10 & _T_17522; // @[Switch.scala 41:38:@7290.4]
  assign _T_17525 = select_11 == 5'h10; // @[Switch.scala 41:52:@7292.4]
  assign output_16_11 = io_outValid_11 & _T_17525; // @[Switch.scala 41:38:@7293.4]
  assign _T_17528 = select_12 == 5'h10; // @[Switch.scala 41:52:@7295.4]
  assign output_16_12 = io_outValid_12 & _T_17528; // @[Switch.scala 41:38:@7296.4]
  assign _T_17531 = select_13 == 5'h10; // @[Switch.scala 41:52:@7298.4]
  assign output_16_13 = io_outValid_13 & _T_17531; // @[Switch.scala 41:38:@7299.4]
  assign _T_17534 = select_14 == 5'h10; // @[Switch.scala 41:52:@7301.4]
  assign output_16_14 = io_outValid_14 & _T_17534; // @[Switch.scala 41:38:@7302.4]
  assign _T_17537 = select_15 == 5'h10; // @[Switch.scala 41:52:@7304.4]
  assign output_16_15 = io_outValid_15 & _T_17537; // @[Switch.scala 41:38:@7305.4]
  assign _T_17540 = select_16 == 5'h10; // @[Switch.scala 41:52:@7307.4]
  assign output_16_16 = io_outValid_16 & _T_17540; // @[Switch.scala 41:38:@7308.4]
  assign _T_17543 = select_17 == 5'h10; // @[Switch.scala 41:52:@7310.4]
  assign output_16_17 = io_outValid_17 & _T_17543; // @[Switch.scala 41:38:@7311.4]
  assign _T_17546 = select_18 == 5'h10; // @[Switch.scala 41:52:@7313.4]
  assign output_16_18 = io_outValid_18 & _T_17546; // @[Switch.scala 41:38:@7314.4]
  assign _T_17549 = select_19 == 5'h10; // @[Switch.scala 41:52:@7316.4]
  assign output_16_19 = io_outValid_19 & _T_17549; // @[Switch.scala 41:38:@7317.4]
  assign _T_17552 = select_20 == 5'h10; // @[Switch.scala 41:52:@7319.4]
  assign output_16_20 = io_outValid_20 & _T_17552; // @[Switch.scala 41:38:@7320.4]
  assign _T_17555 = select_21 == 5'h10; // @[Switch.scala 41:52:@7322.4]
  assign output_16_21 = io_outValid_21 & _T_17555; // @[Switch.scala 41:38:@7323.4]
  assign _T_17558 = select_22 == 5'h10; // @[Switch.scala 41:52:@7325.4]
  assign output_16_22 = io_outValid_22 & _T_17558; // @[Switch.scala 41:38:@7326.4]
  assign _T_17561 = select_23 == 5'h10; // @[Switch.scala 41:52:@7328.4]
  assign output_16_23 = io_outValid_23 & _T_17561; // @[Switch.scala 41:38:@7329.4]
  assign _T_17564 = select_24 == 5'h10; // @[Switch.scala 41:52:@7331.4]
  assign output_16_24 = io_outValid_24 & _T_17564; // @[Switch.scala 41:38:@7332.4]
  assign _T_17567 = select_25 == 5'h10; // @[Switch.scala 41:52:@7334.4]
  assign output_16_25 = io_outValid_25 & _T_17567; // @[Switch.scala 41:38:@7335.4]
  assign _T_17570 = select_26 == 5'h10; // @[Switch.scala 41:52:@7337.4]
  assign output_16_26 = io_outValid_26 & _T_17570; // @[Switch.scala 41:38:@7338.4]
  assign _T_17573 = select_27 == 5'h10; // @[Switch.scala 41:52:@7340.4]
  assign output_16_27 = io_outValid_27 & _T_17573; // @[Switch.scala 41:38:@7341.4]
  assign _T_17576 = select_28 == 5'h10; // @[Switch.scala 41:52:@7343.4]
  assign output_16_28 = io_outValid_28 & _T_17576; // @[Switch.scala 41:38:@7344.4]
  assign _T_17579 = select_29 == 5'h10; // @[Switch.scala 41:52:@7346.4]
  assign output_16_29 = io_outValid_29 & _T_17579; // @[Switch.scala 41:38:@7347.4]
  assign _T_17582 = select_30 == 5'h10; // @[Switch.scala 41:52:@7349.4]
  assign output_16_30 = io_outValid_30 & _T_17582; // @[Switch.scala 41:38:@7350.4]
  assign _T_17585 = select_31 == 5'h10; // @[Switch.scala 41:52:@7352.4]
  assign output_16_31 = io_outValid_31 & _T_17585; // @[Switch.scala 41:38:@7353.4]
  assign _T_17593 = {output_16_7,output_16_6,output_16_5,output_16_4,output_16_3,output_16_2,output_16_1,output_16_0}; // @[Switch.scala 43:31:@7361.4]
  assign _T_17601 = {output_16_15,output_16_14,output_16_13,output_16_12,output_16_11,output_16_10,output_16_9,output_16_8,_T_17593}; // @[Switch.scala 43:31:@7369.4]
  assign _T_17608 = {output_16_23,output_16_22,output_16_21,output_16_20,output_16_19,output_16_18,output_16_17,output_16_16}; // @[Switch.scala 43:31:@7376.4]
  assign _T_17617 = {output_16_31,output_16_30,output_16_29,output_16_28,output_16_27,output_16_26,output_16_25,output_16_24,_T_17608,_T_17601}; // @[Switch.scala 43:31:@7385.4]
  assign _T_17621 = select_0 == 5'h11; // @[Switch.scala 41:52:@7388.4]
  assign output_17_0 = io_outValid_0 & _T_17621; // @[Switch.scala 41:38:@7389.4]
  assign _T_17624 = select_1 == 5'h11; // @[Switch.scala 41:52:@7391.4]
  assign output_17_1 = io_outValid_1 & _T_17624; // @[Switch.scala 41:38:@7392.4]
  assign _T_17627 = select_2 == 5'h11; // @[Switch.scala 41:52:@7394.4]
  assign output_17_2 = io_outValid_2 & _T_17627; // @[Switch.scala 41:38:@7395.4]
  assign _T_17630 = select_3 == 5'h11; // @[Switch.scala 41:52:@7397.4]
  assign output_17_3 = io_outValid_3 & _T_17630; // @[Switch.scala 41:38:@7398.4]
  assign _T_17633 = select_4 == 5'h11; // @[Switch.scala 41:52:@7400.4]
  assign output_17_4 = io_outValid_4 & _T_17633; // @[Switch.scala 41:38:@7401.4]
  assign _T_17636 = select_5 == 5'h11; // @[Switch.scala 41:52:@7403.4]
  assign output_17_5 = io_outValid_5 & _T_17636; // @[Switch.scala 41:38:@7404.4]
  assign _T_17639 = select_6 == 5'h11; // @[Switch.scala 41:52:@7406.4]
  assign output_17_6 = io_outValid_6 & _T_17639; // @[Switch.scala 41:38:@7407.4]
  assign _T_17642 = select_7 == 5'h11; // @[Switch.scala 41:52:@7409.4]
  assign output_17_7 = io_outValid_7 & _T_17642; // @[Switch.scala 41:38:@7410.4]
  assign _T_17645 = select_8 == 5'h11; // @[Switch.scala 41:52:@7412.4]
  assign output_17_8 = io_outValid_8 & _T_17645; // @[Switch.scala 41:38:@7413.4]
  assign _T_17648 = select_9 == 5'h11; // @[Switch.scala 41:52:@7415.4]
  assign output_17_9 = io_outValid_9 & _T_17648; // @[Switch.scala 41:38:@7416.4]
  assign _T_17651 = select_10 == 5'h11; // @[Switch.scala 41:52:@7418.4]
  assign output_17_10 = io_outValid_10 & _T_17651; // @[Switch.scala 41:38:@7419.4]
  assign _T_17654 = select_11 == 5'h11; // @[Switch.scala 41:52:@7421.4]
  assign output_17_11 = io_outValid_11 & _T_17654; // @[Switch.scala 41:38:@7422.4]
  assign _T_17657 = select_12 == 5'h11; // @[Switch.scala 41:52:@7424.4]
  assign output_17_12 = io_outValid_12 & _T_17657; // @[Switch.scala 41:38:@7425.4]
  assign _T_17660 = select_13 == 5'h11; // @[Switch.scala 41:52:@7427.4]
  assign output_17_13 = io_outValid_13 & _T_17660; // @[Switch.scala 41:38:@7428.4]
  assign _T_17663 = select_14 == 5'h11; // @[Switch.scala 41:52:@7430.4]
  assign output_17_14 = io_outValid_14 & _T_17663; // @[Switch.scala 41:38:@7431.4]
  assign _T_17666 = select_15 == 5'h11; // @[Switch.scala 41:52:@7433.4]
  assign output_17_15 = io_outValid_15 & _T_17666; // @[Switch.scala 41:38:@7434.4]
  assign _T_17669 = select_16 == 5'h11; // @[Switch.scala 41:52:@7436.4]
  assign output_17_16 = io_outValid_16 & _T_17669; // @[Switch.scala 41:38:@7437.4]
  assign _T_17672 = select_17 == 5'h11; // @[Switch.scala 41:52:@7439.4]
  assign output_17_17 = io_outValid_17 & _T_17672; // @[Switch.scala 41:38:@7440.4]
  assign _T_17675 = select_18 == 5'h11; // @[Switch.scala 41:52:@7442.4]
  assign output_17_18 = io_outValid_18 & _T_17675; // @[Switch.scala 41:38:@7443.4]
  assign _T_17678 = select_19 == 5'h11; // @[Switch.scala 41:52:@7445.4]
  assign output_17_19 = io_outValid_19 & _T_17678; // @[Switch.scala 41:38:@7446.4]
  assign _T_17681 = select_20 == 5'h11; // @[Switch.scala 41:52:@7448.4]
  assign output_17_20 = io_outValid_20 & _T_17681; // @[Switch.scala 41:38:@7449.4]
  assign _T_17684 = select_21 == 5'h11; // @[Switch.scala 41:52:@7451.4]
  assign output_17_21 = io_outValid_21 & _T_17684; // @[Switch.scala 41:38:@7452.4]
  assign _T_17687 = select_22 == 5'h11; // @[Switch.scala 41:52:@7454.4]
  assign output_17_22 = io_outValid_22 & _T_17687; // @[Switch.scala 41:38:@7455.4]
  assign _T_17690 = select_23 == 5'h11; // @[Switch.scala 41:52:@7457.4]
  assign output_17_23 = io_outValid_23 & _T_17690; // @[Switch.scala 41:38:@7458.4]
  assign _T_17693 = select_24 == 5'h11; // @[Switch.scala 41:52:@7460.4]
  assign output_17_24 = io_outValid_24 & _T_17693; // @[Switch.scala 41:38:@7461.4]
  assign _T_17696 = select_25 == 5'h11; // @[Switch.scala 41:52:@7463.4]
  assign output_17_25 = io_outValid_25 & _T_17696; // @[Switch.scala 41:38:@7464.4]
  assign _T_17699 = select_26 == 5'h11; // @[Switch.scala 41:52:@7466.4]
  assign output_17_26 = io_outValid_26 & _T_17699; // @[Switch.scala 41:38:@7467.4]
  assign _T_17702 = select_27 == 5'h11; // @[Switch.scala 41:52:@7469.4]
  assign output_17_27 = io_outValid_27 & _T_17702; // @[Switch.scala 41:38:@7470.4]
  assign _T_17705 = select_28 == 5'h11; // @[Switch.scala 41:52:@7472.4]
  assign output_17_28 = io_outValid_28 & _T_17705; // @[Switch.scala 41:38:@7473.4]
  assign _T_17708 = select_29 == 5'h11; // @[Switch.scala 41:52:@7475.4]
  assign output_17_29 = io_outValid_29 & _T_17708; // @[Switch.scala 41:38:@7476.4]
  assign _T_17711 = select_30 == 5'h11; // @[Switch.scala 41:52:@7478.4]
  assign output_17_30 = io_outValid_30 & _T_17711; // @[Switch.scala 41:38:@7479.4]
  assign _T_17714 = select_31 == 5'h11; // @[Switch.scala 41:52:@7481.4]
  assign output_17_31 = io_outValid_31 & _T_17714; // @[Switch.scala 41:38:@7482.4]
  assign _T_17722 = {output_17_7,output_17_6,output_17_5,output_17_4,output_17_3,output_17_2,output_17_1,output_17_0}; // @[Switch.scala 43:31:@7490.4]
  assign _T_17730 = {output_17_15,output_17_14,output_17_13,output_17_12,output_17_11,output_17_10,output_17_9,output_17_8,_T_17722}; // @[Switch.scala 43:31:@7498.4]
  assign _T_17737 = {output_17_23,output_17_22,output_17_21,output_17_20,output_17_19,output_17_18,output_17_17,output_17_16}; // @[Switch.scala 43:31:@7505.4]
  assign _T_17746 = {output_17_31,output_17_30,output_17_29,output_17_28,output_17_27,output_17_26,output_17_25,output_17_24,_T_17737,_T_17730}; // @[Switch.scala 43:31:@7514.4]
  assign _T_17750 = select_0 == 5'h12; // @[Switch.scala 41:52:@7517.4]
  assign output_18_0 = io_outValid_0 & _T_17750; // @[Switch.scala 41:38:@7518.4]
  assign _T_17753 = select_1 == 5'h12; // @[Switch.scala 41:52:@7520.4]
  assign output_18_1 = io_outValid_1 & _T_17753; // @[Switch.scala 41:38:@7521.4]
  assign _T_17756 = select_2 == 5'h12; // @[Switch.scala 41:52:@7523.4]
  assign output_18_2 = io_outValid_2 & _T_17756; // @[Switch.scala 41:38:@7524.4]
  assign _T_17759 = select_3 == 5'h12; // @[Switch.scala 41:52:@7526.4]
  assign output_18_3 = io_outValid_3 & _T_17759; // @[Switch.scala 41:38:@7527.4]
  assign _T_17762 = select_4 == 5'h12; // @[Switch.scala 41:52:@7529.4]
  assign output_18_4 = io_outValid_4 & _T_17762; // @[Switch.scala 41:38:@7530.4]
  assign _T_17765 = select_5 == 5'h12; // @[Switch.scala 41:52:@7532.4]
  assign output_18_5 = io_outValid_5 & _T_17765; // @[Switch.scala 41:38:@7533.4]
  assign _T_17768 = select_6 == 5'h12; // @[Switch.scala 41:52:@7535.4]
  assign output_18_6 = io_outValid_6 & _T_17768; // @[Switch.scala 41:38:@7536.4]
  assign _T_17771 = select_7 == 5'h12; // @[Switch.scala 41:52:@7538.4]
  assign output_18_7 = io_outValid_7 & _T_17771; // @[Switch.scala 41:38:@7539.4]
  assign _T_17774 = select_8 == 5'h12; // @[Switch.scala 41:52:@7541.4]
  assign output_18_8 = io_outValid_8 & _T_17774; // @[Switch.scala 41:38:@7542.4]
  assign _T_17777 = select_9 == 5'h12; // @[Switch.scala 41:52:@7544.4]
  assign output_18_9 = io_outValid_9 & _T_17777; // @[Switch.scala 41:38:@7545.4]
  assign _T_17780 = select_10 == 5'h12; // @[Switch.scala 41:52:@7547.4]
  assign output_18_10 = io_outValid_10 & _T_17780; // @[Switch.scala 41:38:@7548.4]
  assign _T_17783 = select_11 == 5'h12; // @[Switch.scala 41:52:@7550.4]
  assign output_18_11 = io_outValid_11 & _T_17783; // @[Switch.scala 41:38:@7551.4]
  assign _T_17786 = select_12 == 5'h12; // @[Switch.scala 41:52:@7553.4]
  assign output_18_12 = io_outValid_12 & _T_17786; // @[Switch.scala 41:38:@7554.4]
  assign _T_17789 = select_13 == 5'h12; // @[Switch.scala 41:52:@7556.4]
  assign output_18_13 = io_outValid_13 & _T_17789; // @[Switch.scala 41:38:@7557.4]
  assign _T_17792 = select_14 == 5'h12; // @[Switch.scala 41:52:@7559.4]
  assign output_18_14 = io_outValid_14 & _T_17792; // @[Switch.scala 41:38:@7560.4]
  assign _T_17795 = select_15 == 5'h12; // @[Switch.scala 41:52:@7562.4]
  assign output_18_15 = io_outValid_15 & _T_17795; // @[Switch.scala 41:38:@7563.4]
  assign _T_17798 = select_16 == 5'h12; // @[Switch.scala 41:52:@7565.4]
  assign output_18_16 = io_outValid_16 & _T_17798; // @[Switch.scala 41:38:@7566.4]
  assign _T_17801 = select_17 == 5'h12; // @[Switch.scala 41:52:@7568.4]
  assign output_18_17 = io_outValid_17 & _T_17801; // @[Switch.scala 41:38:@7569.4]
  assign _T_17804 = select_18 == 5'h12; // @[Switch.scala 41:52:@7571.4]
  assign output_18_18 = io_outValid_18 & _T_17804; // @[Switch.scala 41:38:@7572.4]
  assign _T_17807 = select_19 == 5'h12; // @[Switch.scala 41:52:@7574.4]
  assign output_18_19 = io_outValid_19 & _T_17807; // @[Switch.scala 41:38:@7575.4]
  assign _T_17810 = select_20 == 5'h12; // @[Switch.scala 41:52:@7577.4]
  assign output_18_20 = io_outValid_20 & _T_17810; // @[Switch.scala 41:38:@7578.4]
  assign _T_17813 = select_21 == 5'h12; // @[Switch.scala 41:52:@7580.4]
  assign output_18_21 = io_outValid_21 & _T_17813; // @[Switch.scala 41:38:@7581.4]
  assign _T_17816 = select_22 == 5'h12; // @[Switch.scala 41:52:@7583.4]
  assign output_18_22 = io_outValid_22 & _T_17816; // @[Switch.scala 41:38:@7584.4]
  assign _T_17819 = select_23 == 5'h12; // @[Switch.scala 41:52:@7586.4]
  assign output_18_23 = io_outValid_23 & _T_17819; // @[Switch.scala 41:38:@7587.4]
  assign _T_17822 = select_24 == 5'h12; // @[Switch.scala 41:52:@7589.4]
  assign output_18_24 = io_outValid_24 & _T_17822; // @[Switch.scala 41:38:@7590.4]
  assign _T_17825 = select_25 == 5'h12; // @[Switch.scala 41:52:@7592.4]
  assign output_18_25 = io_outValid_25 & _T_17825; // @[Switch.scala 41:38:@7593.4]
  assign _T_17828 = select_26 == 5'h12; // @[Switch.scala 41:52:@7595.4]
  assign output_18_26 = io_outValid_26 & _T_17828; // @[Switch.scala 41:38:@7596.4]
  assign _T_17831 = select_27 == 5'h12; // @[Switch.scala 41:52:@7598.4]
  assign output_18_27 = io_outValid_27 & _T_17831; // @[Switch.scala 41:38:@7599.4]
  assign _T_17834 = select_28 == 5'h12; // @[Switch.scala 41:52:@7601.4]
  assign output_18_28 = io_outValid_28 & _T_17834; // @[Switch.scala 41:38:@7602.4]
  assign _T_17837 = select_29 == 5'h12; // @[Switch.scala 41:52:@7604.4]
  assign output_18_29 = io_outValid_29 & _T_17837; // @[Switch.scala 41:38:@7605.4]
  assign _T_17840 = select_30 == 5'h12; // @[Switch.scala 41:52:@7607.4]
  assign output_18_30 = io_outValid_30 & _T_17840; // @[Switch.scala 41:38:@7608.4]
  assign _T_17843 = select_31 == 5'h12; // @[Switch.scala 41:52:@7610.4]
  assign output_18_31 = io_outValid_31 & _T_17843; // @[Switch.scala 41:38:@7611.4]
  assign _T_17851 = {output_18_7,output_18_6,output_18_5,output_18_4,output_18_3,output_18_2,output_18_1,output_18_0}; // @[Switch.scala 43:31:@7619.4]
  assign _T_17859 = {output_18_15,output_18_14,output_18_13,output_18_12,output_18_11,output_18_10,output_18_9,output_18_8,_T_17851}; // @[Switch.scala 43:31:@7627.4]
  assign _T_17866 = {output_18_23,output_18_22,output_18_21,output_18_20,output_18_19,output_18_18,output_18_17,output_18_16}; // @[Switch.scala 43:31:@7634.4]
  assign _T_17875 = {output_18_31,output_18_30,output_18_29,output_18_28,output_18_27,output_18_26,output_18_25,output_18_24,_T_17866,_T_17859}; // @[Switch.scala 43:31:@7643.4]
  assign _T_17879 = select_0 == 5'h13; // @[Switch.scala 41:52:@7646.4]
  assign output_19_0 = io_outValid_0 & _T_17879; // @[Switch.scala 41:38:@7647.4]
  assign _T_17882 = select_1 == 5'h13; // @[Switch.scala 41:52:@7649.4]
  assign output_19_1 = io_outValid_1 & _T_17882; // @[Switch.scala 41:38:@7650.4]
  assign _T_17885 = select_2 == 5'h13; // @[Switch.scala 41:52:@7652.4]
  assign output_19_2 = io_outValid_2 & _T_17885; // @[Switch.scala 41:38:@7653.4]
  assign _T_17888 = select_3 == 5'h13; // @[Switch.scala 41:52:@7655.4]
  assign output_19_3 = io_outValid_3 & _T_17888; // @[Switch.scala 41:38:@7656.4]
  assign _T_17891 = select_4 == 5'h13; // @[Switch.scala 41:52:@7658.4]
  assign output_19_4 = io_outValid_4 & _T_17891; // @[Switch.scala 41:38:@7659.4]
  assign _T_17894 = select_5 == 5'h13; // @[Switch.scala 41:52:@7661.4]
  assign output_19_5 = io_outValid_5 & _T_17894; // @[Switch.scala 41:38:@7662.4]
  assign _T_17897 = select_6 == 5'h13; // @[Switch.scala 41:52:@7664.4]
  assign output_19_6 = io_outValid_6 & _T_17897; // @[Switch.scala 41:38:@7665.4]
  assign _T_17900 = select_7 == 5'h13; // @[Switch.scala 41:52:@7667.4]
  assign output_19_7 = io_outValid_7 & _T_17900; // @[Switch.scala 41:38:@7668.4]
  assign _T_17903 = select_8 == 5'h13; // @[Switch.scala 41:52:@7670.4]
  assign output_19_8 = io_outValid_8 & _T_17903; // @[Switch.scala 41:38:@7671.4]
  assign _T_17906 = select_9 == 5'h13; // @[Switch.scala 41:52:@7673.4]
  assign output_19_9 = io_outValid_9 & _T_17906; // @[Switch.scala 41:38:@7674.4]
  assign _T_17909 = select_10 == 5'h13; // @[Switch.scala 41:52:@7676.4]
  assign output_19_10 = io_outValid_10 & _T_17909; // @[Switch.scala 41:38:@7677.4]
  assign _T_17912 = select_11 == 5'h13; // @[Switch.scala 41:52:@7679.4]
  assign output_19_11 = io_outValid_11 & _T_17912; // @[Switch.scala 41:38:@7680.4]
  assign _T_17915 = select_12 == 5'h13; // @[Switch.scala 41:52:@7682.4]
  assign output_19_12 = io_outValid_12 & _T_17915; // @[Switch.scala 41:38:@7683.4]
  assign _T_17918 = select_13 == 5'h13; // @[Switch.scala 41:52:@7685.4]
  assign output_19_13 = io_outValid_13 & _T_17918; // @[Switch.scala 41:38:@7686.4]
  assign _T_17921 = select_14 == 5'h13; // @[Switch.scala 41:52:@7688.4]
  assign output_19_14 = io_outValid_14 & _T_17921; // @[Switch.scala 41:38:@7689.4]
  assign _T_17924 = select_15 == 5'h13; // @[Switch.scala 41:52:@7691.4]
  assign output_19_15 = io_outValid_15 & _T_17924; // @[Switch.scala 41:38:@7692.4]
  assign _T_17927 = select_16 == 5'h13; // @[Switch.scala 41:52:@7694.4]
  assign output_19_16 = io_outValid_16 & _T_17927; // @[Switch.scala 41:38:@7695.4]
  assign _T_17930 = select_17 == 5'h13; // @[Switch.scala 41:52:@7697.4]
  assign output_19_17 = io_outValid_17 & _T_17930; // @[Switch.scala 41:38:@7698.4]
  assign _T_17933 = select_18 == 5'h13; // @[Switch.scala 41:52:@7700.4]
  assign output_19_18 = io_outValid_18 & _T_17933; // @[Switch.scala 41:38:@7701.4]
  assign _T_17936 = select_19 == 5'h13; // @[Switch.scala 41:52:@7703.4]
  assign output_19_19 = io_outValid_19 & _T_17936; // @[Switch.scala 41:38:@7704.4]
  assign _T_17939 = select_20 == 5'h13; // @[Switch.scala 41:52:@7706.4]
  assign output_19_20 = io_outValid_20 & _T_17939; // @[Switch.scala 41:38:@7707.4]
  assign _T_17942 = select_21 == 5'h13; // @[Switch.scala 41:52:@7709.4]
  assign output_19_21 = io_outValid_21 & _T_17942; // @[Switch.scala 41:38:@7710.4]
  assign _T_17945 = select_22 == 5'h13; // @[Switch.scala 41:52:@7712.4]
  assign output_19_22 = io_outValid_22 & _T_17945; // @[Switch.scala 41:38:@7713.4]
  assign _T_17948 = select_23 == 5'h13; // @[Switch.scala 41:52:@7715.4]
  assign output_19_23 = io_outValid_23 & _T_17948; // @[Switch.scala 41:38:@7716.4]
  assign _T_17951 = select_24 == 5'h13; // @[Switch.scala 41:52:@7718.4]
  assign output_19_24 = io_outValid_24 & _T_17951; // @[Switch.scala 41:38:@7719.4]
  assign _T_17954 = select_25 == 5'h13; // @[Switch.scala 41:52:@7721.4]
  assign output_19_25 = io_outValid_25 & _T_17954; // @[Switch.scala 41:38:@7722.4]
  assign _T_17957 = select_26 == 5'h13; // @[Switch.scala 41:52:@7724.4]
  assign output_19_26 = io_outValid_26 & _T_17957; // @[Switch.scala 41:38:@7725.4]
  assign _T_17960 = select_27 == 5'h13; // @[Switch.scala 41:52:@7727.4]
  assign output_19_27 = io_outValid_27 & _T_17960; // @[Switch.scala 41:38:@7728.4]
  assign _T_17963 = select_28 == 5'h13; // @[Switch.scala 41:52:@7730.4]
  assign output_19_28 = io_outValid_28 & _T_17963; // @[Switch.scala 41:38:@7731.4]
  assign _T_17966 = select_29 == 5'h13; // @[Switch.scala 41:52:@7733.4]
  assign output_19_29 = io_outValid_29 & _T_17966; // @[Switch.scala 41:38:@7734.4]
  assign _T_17969 = select_30 == 5'h13; // @[Switch.scala 41:52:@7736.4]
  assign output_19_30 = io_outValid_30 & _T_17969; // @[Switch.scala 41:38:@7737.4]
  assign _T_17972 = select_31 == 5'h13; // @[Switch.scala 41:52:@7739.4]
  assign output_19_31 = io_outValid_31 & _T_17972; // @[Switch.scala 41:38:@7740.4]
  assign _T_17980 = {output_19_7,output_19_6,output_19_5,output_19_4,output_19_3,output_19_2,output_19_1,output_19_0}; // @[Switch.scala 43:31:@7748.4]
  assign _T_17988 = {output_19_15,output_19_14,output_19_13,output_19_12,output_19_11,output_19_10,output_19_9,output_19_8,_T_17980}; // @[Switch.scala 43:31:@7756.4]
  assign _T_17995 = {output_19_23,output_19_22,output_19_21,output_19_20,output_19_19,output_19_18,output_19_17,output_19_16}; // @[Switch.scala 43:31:@7763.4]
  assign _T_18004 = {output_19_31,output_19_30,output_19_29,output_19_28,output_19_27,output_19_26,output_19_25,output_19_24,_T_17995,_T_17988}; // @[Switch.scala 43:31:@7772.4]
  assign _T_18008 = select_0 == 5'h14; // @[Switch.scala 41:52:@7775.4]
  assign output_20_0 = io_outValid_0 & _T_18008; // @[Switch.scala 41:38:@7776.4]
  assign _T_18011 = select_1 == 5'h14; // @[Switch.scala 41:52:@7778.4]
  assign output_20_1 = io_outValid_1 & _T_18011; // @[Switch.scala 41:38:@7779.4]
  assign _T_18014 = select_2 == 5'h14; // @[Switch.scala 41:52:@7781.4]
  assign output_20_2 = io_outValid_2 & _T_18014; // @[Switch.scala 41:38:@7782.4]
  assign _T_18017 = select_3 == 5'h14; // @[Switch.scala 41:52:@7784.4]
  assign output_20_3 = io_outValid_3 & _T_18017; // @[Switch.scala 41:38:@7785.4]
  assign _T_18020 = select_4 == 5'h14; // @[Switch.scala 41:52:@7787.4]
  assign output_20_4 = io_outValid_4 & _T_18020; // @[Switch.scala 41:38:@7788.4]
  assign _T_18023 = select_5 == 5'h14; // @[Switch.scala 41:52:@7790.4]
  assign output_20_5 = io_outValid_5 & _T_18023; // @[Switch.scala 41:38:@7791.4]
  assign _T_18026 = select_6 == 5'h14; // @[Switch.scala 41:52:@7793.4]
  assign output_20_6 = io_outValid_6 & _T_18026; // @[Switch.scala 41:38:@7794.4]
  assign _T_18029 = select_7 == 5'h14; // @[Switch.scala 41:52:@7796.4]
  assign output_20_7 = io_outValid_7 & _T_18029; // @[Switch.scala 41:38:@7797.4]
  assign _T_18032 = select_8 == 5'h14; // @[Switch.scala 41:52:@7799.4]
  assign output_20_8 = io_outValid_8 & _T_18032; // @[Switch.scala 41:38:@7800.4]
  assign _T_18035 = select_9 == 5'h14; // @[Switch.scala 41:52:@7802.4]
  assign output_20_9 = io_outValid_9 & _T_18035; // @[Switch.scala 41:38:@7803.4]
  assign _T_18038 = select_10 == 5'h14; // @[Switch.scala 41:52:@7805.4]
  assign output_20_10 = io_outValid_10 & _T_18038; // @[Switch.scala 41:38:@7806.4]
  assign _T_18041 = select_11 == 5'h14; // @[Switch.scala 41:52:@7808.4]
  assign output_20_11 = io_outValid_11 & _T_18041; // @[Switch.scala 41:38:@7809.4]
  assign _T_18044 = select_12 == 5'h14; // @[Switch.scala 41:52:@7811.4]
  assign output_20_12 = io_outValid_12 & _T_18044; // @[Switch.scala 41:38:@7812.4]
  assign _T_18047 = select_13 == 5'h14; // @[Switch.scala 41:52:@7814.4]
  assign output_20_13 = io_outValid_13 & _T_18047; // @[Switch.scala 41:38:@7815.4]
  assign _T_18050 = select_14 == 5'h14; // @[Switch.scala 41:52:@7817.4]
  assign output_20_14 = io_outValid_14 & _T_18050; // @[Switch.scala 41:38:@7818.4]
  assign _T_18053 = select_15 == 5'h14; // @[Switch.scala 41:52:@7820.4]
  assign output_20_15 = io_outValid_15 & _T_18053; // @[Switch.scala 41:38:@7821.4]
  assign _T_18056 = select_16 == 5'h14; // @[Switch.scala 41:52:@7823.4]
  assign output_20_16 = io_outValid_16 & _T_18056; // @[Switch.scala 41:38:@7824.4]
  assign _T_18059 = select_17 == 5'h14; // @[Switch.scala 41:52:@7826.4]
  assign output_20_17 = io_outValid_17 & _T_18059; // @[Switch.scala 41:38:@7827.4]
  assign _T_18062 = select_18 == 5'h14; // @[Switch.scala 41:52:@7829.4]
  assign output_20_18 = io_outValid_18 & _T_18062; // @[Switch.scala 41:38:@7830.4]
  assign _T_18065 = select_19 == 5'h14; // @[Switch.scala 41:52:@7832.4]
  assign output_20_19 = io_outValid_19 & _T_18065; // @[Switch.scala 41:38:@7833.4]
  assign _T_18068 = select_20 == 5'h14; // @[Switch.scala 41:52:@7835.4]
  assign output_20_20 = io_outValid_20 & _T_18068; // @[Switch.scala 41:38:@7836.4]
  assign _T_18071 = select_21 == 5'h14; // @[Switch.scala 41:52:@7838.4]
  assign output_20_21 = io_outValid_21 & _T_18071; // @[Switch.scala 41:38:@7839.4]
  assign _T_18074 = select_22 == 5'h14; // @[Switch.scala 41:52:@7841.4]
  assign output_20_22 = io_outValid_22 & _T_18074; // @[Switch.scala 41:38:@7842.4]
  assign _T_18077 = select_23 == 5'h14; // @[Switch.scala 41:52:@7844.4]
  assign output_20_23 = io_outValid_23 & _T_18077; // @[Switch.scala 41:38:@7845.4]
  assign _T_18080 = select_24 == 5'h14; // @[Switch.scala 41:52:@7847.4]
  assign output_20_24 = io_outValid_24 & _T_18080; // @[Switch.scala 41:38:@7848.4]
  assign _T_18083 = select_25 == 5'h14; // @[Switch.scala 41:52:@7850.4]
  assign output_20_25 = io_outValid_25 & _T_18083; // @[Switch.scala 41:38:@7851.4]
  assign _T_18086 = select_26 == 5'h14; // @[Switch.scala 41:52:@7853.4]
  assign output_20_26 = io_outValid_26 & _T_18086; // @[Switch.scala 41:38:@7854.4]
  assign _T_18089 = select_27 == 5'h14; // @[Switch.scala 41:52:@7856.4]
  assign output_20_27 = io_outValid_27 & _T_18089; // @[Switch.scala 41:38:@7857.4]
  assign _T_18092 = select_28 == 5'h14; // @[Switch.scala 41:52:@7859.4]
  assign output_20_28 = io_outValid_28 & _T_18092; // @[Switch.scala 41:38:@7860.4]
  assign _T_18095 = select_29 == 5'h14; // @[Switch.scala 41:52:@7862.4]
  assign output_20_29 = io_outValid_29 & _T_18095; // @[Switch.scala 41:38:@7863.4]
  assign _T_18098 = select_30 == 5'h14; // @[Switch.scala 41:52:@7865.4]
  assign output_20_30 = io_outValid_30 & _T_18098; // @[Switch.scala 41:38:@7866.4]
  assign _T_18101 = select_31 == 5'h14; // @[Switch.scala 41:52:@7868.4]
  assign output_20_31 = io_outValid_31 & _T_18101; // @[Switch.scala 41:38:@7869.4]
  assign _T_18109 = {output_20_7,output_20_6,output_20_5,output_20_4,output_20_3,output_20_2,output_20_1,output_20_0}; // @[Switch.scala 43:31:@7877.4]
  assign _T_18117 = {output_20_15,output_20_14,output_20_13,output_20_12,output_20_11,output_20_10,output_20_9,output_20_8,_T_18109}; // @[Switch.scala 43:31:@7885.4]
  assign _T_18124 = {output_20_23,output_20_22,output_20_21,output_20_20,output_20_19,output_20_18,output_20_17,output_20_16}; // @[Switch.scala 43:31:@7892.4]
  assign _T_18133 = {output_20_31,output_20_30,output_20_29,output_20_28,output_20_27,output_20_26,output_20_25,output_20_24,_T_18124,_T_18117}; // @[Switch.scala 43:31:@7901.4]
  assign _T_18137 = select_0 == 5'h15; // @[Switch.scala 41:52:@7904.4]
  assign output_21_0 = io_outValid_0 & _T_18137; // @[Switch.scala 41:38:@7905.4]
  assign _T_18140 = select_1 == 5'h15; // @[Switch.scala 41:52:@7907.4]
  assign output_21_1 = io_outValid_1 & _T_18140; // @[Switch.scala 41:38:@7908.4]
  assign _T_18143 = select_2 == 5'h15; // @[Switch.scala 41:52:@7910.4]
  assign output_21_2 = io_outValid_2 & _T_18143; // @[Switch.scala 41:38:@7911.4]
  assign _T_18146 = select_3 == 5'h15; // @[Switch.scala 41:52:@7913.4]
  assign output_21_3 = io_outValid_3 & _T_18146; // @[Switch.scala 41:38:@7914.4]
  assign _T_18149 = select_4 == 5'h15; // @[Switch.scala 41:52:@7916.4]
  assign output_21_4 = io_outValid_4 & _T_18149; // @[Switch.scala 41:38:@7917.4]
  assign _T_18152 = select_5 == 5'h15; // @[Switch.scala 41:52:@7919.4]
  assign output_21_5 = io_outValid_5 & _T_18152; // @[Switch.scala 41:38:@7920.4]
  assign _T_18155 = select_6 == 5'h15; // @[Switch.scala 41:52:@7922.4]
  assign output_21_6 = io_outValid_6 & _T_18155; // @[Switch.scala 41:38:@7923.4]
  assign _T_18158 = select_7 == 5'h15; // @[Switch.scala 41:52:@7925.4]
  assign output_21_7 = io_outValid_7 & _T_18158; // @[Switch.scala 41:38:@7926.4]
  assign _T_18161 = select_8 == 5'h15; // @[Switch.scala 41:52:@7928.4]
  assign output_21_8 = io_outValid_8 & _T_18161; // @[Switch.scala 41:38:@7929.4]
  assign _T_18164 = select_9 == 5'h15; // @[Switch.scala 41:52:@7931.4]
  assign output_21_9 = io_outValid_9 & _T_18164; // @[Switch.scala 41:38:@7932.4]
  assign _T_18167 = select_10 == 5'h15; // @[Switch.scala 41:52:@7934.4]
  assign output_21_10 = io_outValid_10 & _T_18167; // @[Switch.scala 41:38:@7935.4]
  assign _T_18170 = select_11 == 5'h15; // @[Switch.scala 41:52:@7937.4]
  assign output_21_11 = io_outValid_11 & _T_18170; // @[Switch.scala 41:38:@7938.4]
  assign _T_18173 = select_12 == 5'h15; // @[Switch.scala 41:52:@7940.4]
  assign output_21_12 = io_outValid_12 & _T_18173; // @[Switch.scala 41:38:@7941.4]
  assign _T_18176 = select_13 == 5'h15; // @[Switch.scala 41:52:@7943.4]
  assign output_21_13 = io_outValid_13 & _T_18176; // @[Switch.scala 41:38:@7944.4]
  assign _T_18179 = select_14 == 5'h15; // @[Switch.scala 41:52:@7946.4]
  assign output_21_14 = io_outValid_14 & _T_18179; // @[Switch.scala 41:38:@7947.4]
  assign _T_18182 = select_15 == 5'h15; // @[Switch.scala 41:52:@7949.4]
  assign output_21_15 = io_outValid_15 & _T_18182; // @[Switch.scala 41:38:@7950.4]
  assign _T_18185 = select_16 == 5'h15; // @[Switch.scala 41:52:@7952.4]
  assign output_21_16 = io_outValid_16 & _T_18185; // @[Switch.scala 41:38:@7953.4]
  assign _T_18188 = select_17 == 5'h15; // @[Switch.scala 41:52:@7955.4]
  assign output_21_17 = io_outValid_17 & _T_18188; // @[Switch.scala 41:38:@7956.4]
  assign _T_18191 = select_18 == 5'h15; // @[Switch.scala 41:52:@7958.4]
  assign output_21_18 = io_outValid_18 & _T_18191; // @[Switch.scala 41:38:@7959.4]
  assign _T_18194 = select_19 == 5'h15; // @[Switch.scala 41:52:@7961.4]
  assign output_21_19 = io_outValid_19 & _T_18194; // @[Switch.scala 41:38:@7962.4]
  assign _T_18197 = select_20 == 5'h15; // @[Switch.scala 41:52:@7964.4]
  assign output_21_20 = io_outValid_20 & _T_18197; // @[Switch.scala 41:38:@7965.4]
  assign _T_18200 = select_21 == 5'h15; // @[Switch.scala 41:52:@7967.4]
  assign output_21_21 = io_outValid_21 & _T_18200; // @[Switch.scala 41:38:@7968.4]
  assign _T_18203 = select_22 == 5'h15; // @[Switch.scala 41:52:@7970.4]
  assign output_21_22 = io_outValid_22 & _T_18203; // @[Switch.scala 41:38:@7971.4]
  assign _T_18206 = select_23 == 5'h15; // @[Switch.scala 41:52:@7973.4]
  assign output_21_23 = io_outValid_23 & _T_18206; // @[Switch.scala 41:38:@7974.4]
  assign _T_18209 = select_24 == 5'h15; // @[Switch.scala 41:52:@7976.4]
  assign output_21_24 = io_outValid_24 & _T_18209; // @[Switch.scala 41:38:@7977.4]
  assign _T_18212 = select_25 == 5'h15; // @[Switch.scala 41:52:@7979.4]
  assign output_21_25 = io_outValid_25 & _T_18212; // @[Switch.scala 41:38:@7980.4]
  assign _T_18215 = select_26 == 5'h15; // @[Switch.scala 41:52:@7982.4]
  assign output_21_26 = io_outValid_26 & _T_18215; // @[Switch.scala 41:38:@7983.4]
  assign _T_18218 = select_27 == 5'h15; // @[Switch.scala 41:52:@7985.4]
  assign output_21_27 = io_outValid_27 & _T_18218; // @[Switch.scala 41:38:@7986.4]
  assign _T_18221 = select_28 == 5'h15; // @[Switch.scala 41:52:@7988.4]
  assign output_21_28 = io_outValid_28 & _T_18221; // @[Switch.scala 41:38:@7989.4]
  assign _T_18224 = select_29 == 5'h15; // @[Switch.scala 41:52:@7991.4]
  assign output_21_29 = io_outValid_29 & _T_18224; // @[Switch.scala 41:38:@7992.4]
  assign _T_18227 = select_30 == 5'h15; // @[Switch.scala 41:52:@7994.4]
  assign output_21_30 = io_outValid_30 & _T_18227; // @[Switch.scala 41:38:@7995.4]
  assign _T_18230 = select_31 == 5'h15; // @[Switch.scala 41:52:@7997.4]
  assign output_21_31 = io_outValid_31 & _T_18230; // @[Switch.scala 41:38:@7998.4]
  assign _T_18238 = {output_21_7,output_21_6,output_21_5,output_21_4,output_21_3,output_21_2,output_21_1,output_21_0}; // @[Switch.scala 43:31:@8006.4]
  assign _T_18246 = {output_21_15,output_21_14,output_21_13,output_21_12,output_21_11,output_21_10,output_21_9,output_21_8,_T_18238}; // @[Switch.scala 43:31:@8014.4]
  assign _T_18253 = {output_21_23,output_21_22,output_21_21,output_21_20,output_21_19,output_21_18,output_21_17,output_21_16}; // @[Switch.scala 43:31:@8021.4]
  assign _T_18262 = {output_21_31,output_21_30,output_21_29,output_21_28,output_21_27,output_21_26,output_21_25,output_21_24,_T_18253,_T_18246}; // @[Switch.scala 43:31:@8030.4]
  assign _T_18266 = select_0 == 5'h16; // @[Switch.scala 41:52:@8033.4]
  assign output_22_0 = io_outValid_0 & _T_18266; // @[Switch.scala 41:38:@8034.4]
  assign _T_18269 = select_1 == 5'h16; // @[Switch.scala 41:52:@8036.4]
  assign output_22_1 = io_outValid_1 & _T_18269; // @[Switch.scala 41:38:@8037.4]
  assign _T_18272 = select_2 == 5'h16; // @[Switch.scala 41:52:@8039.4]
  assign output_22_2 = io_outValid_2 & _T_18272; // @[Switch.scala 41:38:@8040.4]
  assign _T_18275 = select_3 == 5'h16; // @[Switch.scala 41:52:@8042.4]
  assign output_22_3 = io_outValid_3 & _T_18275; // @[Switch.scala 41:38:@8043.4]
  assign _T_18278 = select_4 == 5'h16; // @[Switch.scala 41:52:@8045.4]
  assign output_22_4 = io_outValid_4 & _T_18278; // @[Switch.scala 41:38:@8046.4]
  assign _T_18281 = select_5 == 5'h16; // @[Switch.scala 41:52:@8048.4]
  assign output_22_5 = io_outValid_5 & _T_18281; // @[Switch.scala 41:38:@8049.4]
  assign _T_18284 = select_6 == 5'h16; // @[Switch.scala 41:52:@8051.4]
  assign output_22_6 = io_outValid_6 & _T_18284; // @[Switch.scala 41:38:@8052.4]
  assign _T_18287 = select_7 == 5'h16; // @[Switch.scala 41:52:@8054.4]
  assign output_22_7 = io_outValid_7 & _T_18287; // @[Switch.scala 41:38:@8055.4]
  assign _T_18290 = select_8 == 5'h16; // @[Switch.scala 41:52:@8057.4]
  assign output_22_8 = io_outValid_8 & _T_18290; // @[Switch.scala 41:38:@8058.4]
  assign _T_18293 = select_9 == 5'h16; // @[Switch.scala 41:52:@8060.4]
  assign output_22_9 = io_outValid_9 & _T_18293; // @[Switch.scala 41:38:@8061.4]
  assign _T_18296 = select_10 == 5'h16; // @[Switch.scala 41:52:@8063.4]
  assign output_22_10 = io_outValid_10 & _T_18296; // @[Switch.scala 41:38:@8064.4]
  assign _T_18299 = select_11 == 5'h16; // @[Switch.scala 41:52:@8066.4]
  assign output_22_11 = io_outValid_11 & _T_18299; // @[Switch.scala 41:38:@8067.4]
  assign _T_18302 = select_12 == 5'h16; // @[Switch.scala 41:52:@8069.4]
  assign output_22_12 = io_outValid_12 & _T_18302; // @[Switch.scala 41:38:@8070.4]
  assign _T_18305 = select_13 == 5'h16; // @[Switch.scala 41:52:@8072.4]
  assign output_22_13 = io_outValid_13 & _T_18305; // @[Switch.scala 41:38:@8073.4]
  assign _T_18308 = select_14 == 5'h16; // @[Switch.scala 41:52:@8075.4]
  assign output_22_14 = io_outValid_14 & _T_18308; // @[Switch.scala 41:38:@8076.4]
  assign _T_18311 = select_15 == 5'h16; // @[Switch.scala 41:52:@8078.4]
  assign output_22_15 = io_outValid_15 & _T_18311; // @[Switch.scala 41:38:@8079.4]
  assign _T_18314 = select_16 == 5'h16; // @[Switch.scala 41:52:@8081.4]
  assign output_22_16 = io_outValid_16 & _T_18314; // @[Switch.scala 41:38:@8082.4]
  assign _T_18317 = select_17 == 5'h16; // @[Switch.scala 41:52:@8084.4]
  assign output_22_17 = io_outValid_17 & _T_18317; // @[Switch.scala 41:38:@8085.4]
  assign _T_18320 = select_18 == 5'h16; // @[Switch.scala 41:52:@8087.4]
  assign output_22_18 = io_outValid_18 & _T_18320; // @[Switch.scala 41:38:@8088.4]
  assign _T_18323 = select_19 == 5'h16; // @[Switch.scala 41:52:@8090.4]
  assign output_22_19 = io_outValid_19 & _T_18323; // @[Switch.scala 41:38:@8091.4]
  assign _T_18326 = select_20 == 5'h16; // @[Switch.scala 41:52:@8093.4]
  assign output_22_20 = io_outValid_20 & _T_18326; // @[Switch.scala 41:38:@8094.4]
  assign _T_18329 = select_21 == 5'h16; // @[Switch.scala 41:52:@8096.4]
  assign output_22_21 = io_outValid_21 & _T_18329; // @[Switch.scala 41:38:@8097.4]
  assign _T_18332 = select_22 == 5'h16; // @[Switch.scala 41:52:@8099.4]
  assign output_22_22 = io_outValid_22 & _T_18332; // @[Switch.scala 41:38:@8100.4]
  assign _T_18335 = select_23 == 5'h16; // @[Switch.scala 41:52:@8102.4]
  assign output_22_23 = io_outValid_23 & _T_18335; // @[Switch.scala 41:38:@8103.4]
  assign _T_18338 = select_24 == 5'h16; // @[Switch.scala 41:52:@8105.4]
  assign output_22_24 = io_outValid_24 & _T_18338; // @[Switch.scala 41:38:@8106.4]
  assign _T_18341 = select_25 == 5'h16; // @[Switch.scala 41:52:@8108.4]
  assign output_22_25 = io_outValid_25 & _T_18341; // @[Switch.scala 41:38:@8109.4]
  assign _T_18344 = select_26 == 5'h16; // @[Switch.scala 41:52:@8111.4]
  assign output_22_26 = io_outValid_26 & _T_18344; // @[Switch.scala 41:38:@8112.4]
  assign _T_18347 = select_27 == 5'h16; // @[Switch.scala 41:52:@8114.4]
  assign output_22_27 = io_outValid_27 & _T_18347; // @[Switch.scala 41:38:@8115.4]
  assign _T_18350 = select_28 == 5'h16; // @[Switch.scala 41:52:@8117.4]
  assign output_22_28 = io_outValid_28 & _T_18350; // @[Switch.scala 41:38:@8118.4]
  assign _T_18353 = select_29 == 5'h16; // @[Switch.scala 41:52:@8120.4]
  assign output_22_29 = io_outValid_29 & _T_18353; // @[Switch.scala 41:38:@8121.4]
  assign _T_18356 = select_30 == 5'h16; // @[Switch.scala 41:52:@8123.4]
  assign output_22_30 = io_outValid_30 & _T_18356; // @[Switch.scala 41:38:@8124.4]
  assign _T_18359 = select_31 == 5'h16; // @[Switch.scala 41:52:@8126.4]
  assign output_22_31 = io_outValid_31 & _T_18359; // @[Switch.scala 41:38:@8127.4]
  assign _T_18367 = {output_22_7,output_22_6,output_22_5,output_22_4,output_22_3,output_22_2,output_22_1,output_22_0}; // @[Switch.scala 43:31:@8135.4]
  assign _T_18375 = {output_22_15,output_22_14,output_22_13,output_22_12,output_22_11,output_22_10,output_22_9,output_22_8,_T_18367}; // @[Switch.scala 43:31:@8143.4]
  assign _T_18382 = {output_22_23,output_22_22,output_22_21,output_22_20,output_22_19,output_22_18,output_22_17,output_22_16}; // @[Switch.scala 43:31:@8150.4]
  assign _T_18391 = {output_22_31,output_22_30,output_22_29,output_22_28,output_22_27,output_22_26,output_22_25,output_22_24,_T_18382,_T_18375}; // @[Switch.scala 43:31:@8159.4]
  assign _T_18395 = select_0 == 5'h17; // @[Switch.scala 41:52:@8162.4]
  assign output_23_0 = io_outValid_0 & _T_18395; // @[Switch.scala 41:38:@8163.4]
  assign _T_18398 = select_1 == 5'h17; // @[Switch.scala 41:52:@8165.4]
  assign output_23_1 = io_outValid_1 & _T_18398; // @[Switch.scala 41:38:@8166.4]
  assign _T_18401 = select_2 == 5'h17; // @[Switch.scala 41:52:@8168.4]
  assign output_23_2 = io_outValid_2 & _T_18401; // @[Switch.scala 41:38:@8169.4]
  assign _T_18404 = select_3 == 5'h17; // @[Switch.scala 41:52:@8171.4]
  assign output_23_3 = io_outValid_3 & _T_18404; // @[Switch.scala 41:38:@8172.4]
  assign _T_18407 = select_4 == 5'h17; // @[Switch.scala 41:52:@8174.4]
  assign output_23_4 = io_outValid_4 & _T_18407; // @[Switch.scala 41:38:@8175.4]
  assign _T_18410 = select_5 == 5'h17; // @[Switch.scala 41:52:@8177.4]
  assign output_23_5 = io_outValid_5 & _T_18410; // @[Switch.scala 41:38:@8178.4]
  assign _T_18413 = select_6 == 5'h17; // @[Switch.scala 41:52:@8180.4]
  assign output_23_6 = io_outValid_6 & _T_18413; // @[Switch.scala 41:38:@8181.4]
  assign _T_18416 = select_7 == 5'h17; // @[Switch.scala 41:52:@8183.4]
  assign output_23_7 = io_outValid_7 & _T_18416; // @[Switch.scala 41:38:@8184.4]
  assign _T_18419 = select_8 == 5'h17; // @[Switch.scala 41:52:@8186.4]
  assign output_23_8 = io_outValid_8 & _T_18419; // @[Switch.scala 41:38:@8187.4]
  assign _T_18422 = select_9 == 5'h17; // @[Switch.scala 41:52:@8189.4]
  assign output_23_9 = io_outValid_9 & _T_18422; // @[Switch.scala 41:38:@8190.4]
  assign _T_18425 = select_10 == 5'h17; // @[Switch.scala 41:52:@8192.4]
  assign output_23_10 = io_outValid_10 & _T_18425; // @[Switch.scala 41:38:@8193.4]
  assign _T_18428 = select_11 == 5'h17; // @[Switch.scala 41:52:@8195.4]
  assign output_23_11 = io_outValid_11 & _T_18428; // @[Switch.scala 41:38:@8196.4]
  assign _T_18431 = select_12 == 5'h17; // @[Switch.scala 41:52:@8198.4]
  assign output_23_12 = io_outValid_12 & _T_18431; // @[Switch.scala 41:38:@8199.4]
  assign _T_18434 = select_13 == 5'h17; // @[Switch.scala 41:52:@8201.4]
  assign output_23_13 = io_outValid_13 & _T_18434; // @[Switch.scala 41:38:@8202.4]
  assign _T_18437 = select_14 == 5'h17; // @[Switch.scala 41:52:@8204.4]
  assign output_23_14 = io_outValid_14 & _T_18437; // @[Switch.scala 41:38:@8205.4]
  assign _T_18440 = select_15 == 5'h17; // @[Switch.scala 41:52:@8207.4]
  assign output_23_15 = io_outValid_15 & _T_18440; // @[Switch.scala 41:38:@8208.4]
  assign _T_18443 = select_16 == 5'h17; // @[Switch.scala 41:52:@8210.4]
  assign output_23_16 = io_outValid_16 & _T_18443; // @[Switch.scala 41:38:@8211.4]
  assign _T_18446 = select_17 == 5'h17; // @[Switch.scala 41:52:@8213.4]
  assign output_23_17 = io_outValid_17 & _T_18446; // @[Switch.scala 41:38:@8214.4]
  assign _T_18449 = select_18 == 5'h17; // @[Switch.scala 41:52:@8216.4]
  assign output_23_18 = io_outValid_18 & _T_18449; // @[Switch.scala 41:38:@8217.4]
  assign _T_18452 = select_19 == 5'h17; // @[Switch.scala 41:52:@8219.4]
  assign output_23_19 = io_outValid_19 & _T_18452; // @[Switch.scala 41:38:@8220.4]
  assign _T_18455 = select_20 == 5'h17; // @[Switch.scala 41:52:@8222.4]
  assign output_23_20 = io_outValid_20 & _T_18455; // @[Switch.scala 41:38:@8223.4]
  assign _T_18458 = select_21 == 5'h17; // @[Switch.scala 41:52:@8225.4]
  assign output_23_21 = io_outValid_21 & _T_18458; // @[Switch.scala 41:38:@8226.4]
  assign _T_18461 = select_22 == 5'h17; // @[Switch.scala 41:52:@8228.4]
  assign output_23_22 = io_outValid_22 & _T_18461; // @[Switch.scala 41:38:@8229.4]
  assign _T_18464 = select_23 == 5'h17; // @[Switch.scala 41:52:@8231.4]
  assign output_23_23 = io_outValid_23 & _T_18464; // @[Switch.scala 41:38:@8232.4]
  assign _T_18467 = select_24 == 5'h17; // @[Switch.scala 41:52:@8234.4]
  assign output_23_24 = io_outValid_24 & _T_18467; // @[Switch.scala 41:38:@8235.4]
  assign _T_18470 = select_25 == 5'h17; // @[Switch.scala 41:52:@8237.4]
  assign output_23_25 = io_outValid_25 & _T_18470; // @[Switch.scala 41:38:@8238.4]
  assign _T_18473 = select_26 == 5'h17; // @[Switch.scala 41:52:@8240.4]
  assign output_23_26 = io_outValid_26 & _T_18473; // @[Switch.scala 41:38:@8241.4]
  assign _T_18476 = select_27 == 5'h17; // @[Switch.scala 41:52:@8243.4]
  assign output_23_27 = io_outValid_27 & _T_18476; // @[Switch.scala 41:38:@8244.4]
  assign _T_18479 = select_28 == 5'h17; // @[Switch.scala 41:52:@8246.4]
  assign output_23_28 = io_outValid_28 & _T_18479; // @[Switch.scala 41:38:@8247.4]
  assign _T_18482 = select_29 == 5'h17; // @[Switch.scala 41:52:@8249.4]
  assign output_23_29 = io_outValid_29 & _T_18482; // @[Switch.scala 41:38:@8250.4]
  assign _T_18485 = select_30 == 5'h17; // @[Switch.scala 41:52:@8252.4]
  assign output_23_30 = io_outValid_30 & _T_18485; // @[Switch.scala 41:38:@8253.4]
  assign _T_18488 = select_31 == 5'h17; // @[Switch.scala 41:52:@8255.4]
  assign output_23_31 = io_outValid_31 & _T_18488; // @[Switch.scala 41:38:@8256.4]
  assign _T_18496 = {output_23_7,output_23_6,output_23_5,output_23_4,output_23_3,output_23_2,output_23_1,output_23_0}; // @[Switch.scala 43:31:@8264.4]
  assign _T_18504 = {output_23_15,output_23_14,output_23_13,output_23_12,output_23_11,output_23_10,output_23_9,output_23_8,_T_18496}; // @[Switch.scala 43:31:@8272.4]
  assign _T_18511 = {output_23_23,output_23_22,output_23_21,output_23_20,output_23_19,output_23_18,output_23_17,output_23_16}; // @[Switch.scala 43:31:@8279.4]
  assign _T_18520 = {output_23_31,output_23_30,output_23_29,output_23_28,output_23_27,output_23_26,output_23_25,output_23_24,_T_18511,_T_18504}; // @[Switch.scala 43:31:@8288.4]
  assign _T_18524 = select_0 == 5'h18; // @[Switch.scala 41:52:@8291.4]
  assign output_24_0 = io_outValid_0 & _T_18524; // @[Switch.scala 41:38:@8292.4]
  assign _T_18527 = select_1 == 5'h18; // @[Switch.scala 41:52:@8294.4]
  assign output_24_1 = io_outValid_1 & _T_18527; // @[Switch.scala 41:38:@8295.4]
  assign _T_18530 = select_2 == 5'h18; // @[Switch.scala 41:52:@8297.4]
  assign output_24_2 = io_outValid_2 & _T_18530; // @[Switch.scala 41:38:@8298.4]
  assign _T_18533 = select_3 == 5'h18; // @[Switch.scala 41:52:@8300.4]
  assign output_24_3 = io_outValid_3 & _T_18533; // @[Switch.scala 41:38:@8301.4]
  assign _T_18536 = select_4 == 5'h18; // @[Switch.scala 41:52:@8303.4]
  assign output_24_4 = io_outValid_4 & _T_18536; // @[Switch.scala 41:38:@8304.4]
  assign _T_18539 = select_5 == 5'h18; // @[Switch.scala 41:52:@8306.4]
  assign output_24_5 = io_outValid_5 & _T_18539; // @[Switch.scala 41:38:@8307.4]
  assign _T_18542 = select_6 == 5'h18; // @[Switch.scala 41:52:@8309.4]
  assign output_24_6 = io_outValid_6 & _T_18542; // @[Switch.scala 41:38:@8310.4]
  assign _T_18545 = select_7 == 5'h18; // @[Switch.scala 41:52:@8312.4]
  assign output_24_7 = io_outValid_7 & _T_18545; // @[Switch.scala 41:38:@8313.4]
  assign _T_18548 = select_8 == 5'h18; // @[Switch.scala 41:52:@8315.4]
  assign output_24_8 = io_outValid_8 & _T_18548; // @[Switch.scala 41:38:@8316.4]
  assign _T_18551 = select_9 == 5'h18; // @[Switch.scala 41:52:@8318.4]
  assign output_24_9 = io_outValid_9 & _T_18551; // @[Switch.scala 41:38:@8319.4]
  assign _T_18554 = select_10 == 5'h18; // @[Switch.scala 41:52:@8321.4]
  assign output_24_10 = io_outValid_10 & _T_18554; // @[Switch.scala 41:38:@8322.4]
  assign _T_18557 = select_11 == 5'h18; // @[Switch.scala 41:52:@8324.4]
  assign output_24_11 = io_outValid_11 & _T_18557; // @[Switch.scala 41:38:@8325.4]
  assign _T_18560 = select_12 == 5'h18; // @[Switch.scala 41:52:@8327.4]
  assign output_24_12 = io_outValid_12 & _T_18560; // @[Switch.scala 41:38:@8328.4]
  assign _T_18563 = select_13 == 5'h18; // @[Switch.scala 41:52:@8330.4]
  assign output_24_13 = io_outValid_13 & _T_18563; // @[Switch.scala 41:38:@8331.4]
  assign _T_18566 = select_14 == 5'h18; // @[Switch.scala 41:52:@8333.4]
  assign output_24_14 = io_outValid_14 & _T_18566; // @[Switch.scala 41:38:@8334.4]
  assign _T_18569 = select_15 == 5'h18; // @[Switch.scala 41:52:@8336.4]
  assign output_24_15 = io_outValid_15 & _T_18569; // @[Switch.scala 41:38:@8337.4]
  assign _T_18572 = select_16 == 5'h18; // @[Switch.scala 41:52:@8339.4]
  assign output_24_16 = io_outValid_16 & _T_18572; // @[Switch.scala 41:38:@8340.4]
  assign _T_18575 = select_17 == 5'h18; // @[Switch.scala 41:52:@8342.4]
  assign output_24_17 = io_outValid_17 & _T_18575; // @[Switch.scala 41:38:@8343.4]
  assign _T_18578 = select_18 == 5'h18; // @[Switch.scala 41:52:@8345.4]
  assign output_24_18 = io_outValid_18 & _T_18578; // @[Switch.scala 41:38:@8346.4]
  assign _T_18581 = select_19 == 5'h18; // @[Switch.scala 41:52:@8348.4]
  assign output_24_19 = io_outValid_19 & _T_18581; // @[Switch.scala 41:38:@8349.4]
  assign _T_18584 = select_20 == 5'h18; // @[Switch.scala 41:52:@8351.4]
  assign output_24_20 = io_outValid_20 & _T_18584; // @[Switch.scala 41:38:@8352.4]
  assign _T_18587 = select_21 == 5'h18; // @[Switch.scala 41:52:@8354.4]
  assign output_24_21 = io_outValid_21 & _T_18587; // @[Switch.scala 41:38:@8355.4]
  assign _T_18590 = select_22 == 5'h18; // @[Switch.scala 41:52:@8357.4]
  assign output_24_22 = io_outValid_22 & _T_18590; // @[Switch.scala 41:38:@8358.4]
  assign _T_18593 = select_23 == 5'h18; // @[Switch.scala 41:52:@8360.4]
  assign output_24_23 = io_outValid_23 & _T_18593; // @[Switch.scala 41:38:@8361.4]
  assign _T_18596 = select_24 == 5'h18; // @[Switch.scala 41:52:@8363.4]
  assign output_24_24 = io_outValid_24 & _T_18596; // @[Switch.scala 41:38:@8364.4]
  assign _T_18599 = select_25 == 5'h18; // @[Switch.scala 41:52:@8366.4]
  assign output_24_25 = io_outValid_25 & _T_18599; // @[Switch.scala 41:38:@8367.4]
  assign _T_18602 = select_26 == 5'h18; // @[Switch.scala 41:52:@8369.4]
  assign output_24_26 = io_outValid_26 & _T_18602; // @[Switch.scala 41:38:@8370.4]
  assign _T_18605 = select_27 == 5'h18; // @[Switch.scala 41:52:@8372.4]
  assign output_24_27 = io_outValid_27 & _T_18605; // @[Switch.scala 41:38:@8373.4]
  assign _T_18608 = select_28 == 5'h18; // @[Switch.scala 41:52:@8375.4]
  assign output_24_28 = io_outValid_28 & _T_18608; // @[Switch.scala 41:38:@8376.4]
  assign _T_18611 = select_29 == 5'h18; // @[Switch.scala 41:52:@8378.4]
  assign output_24_29 = io_outValid_29 & _T_18611; // @[Switch.scala 41:38:@8379.4]
  assign _T_18614 = select_30 == 5'h18; // @[Switch.scala 41:52:@8381.4]
  assign output_24_30 = io_outValid_30 & _T_18614; // @[Switch.scala 41:38:@8382.4]
  assign _T_18617 = select_31 == 5'h18; // @[Switch.scala 41:52:@8384.4]
  assign output_24_31 = io_outValid_31 & _T_18617; // @[Switch.scala 41:38:@8385.4]
  assign _T_18625 = {output_24_7,output_24_6,output_24_5,output_24_4,output_24_3,output_24_2,output_24_1,output_24_0}; // @[Switch.scala 43:31:@8393.4]
  assign _T_18633 = {output_24_15,output_24_14,output_24_13,output_24_12,output_24_11,output_24_10,output_24_9,output_24_8,_T_18625}; // @[Switch.scala 43:31:@8401.4]
  assign _T_18640 = {output_24_23,output_24_22,output_24_21,output_24_20,output_24_19,output_24_18,output_24_17,output_24_16}; // @[Switch.scala 43:31:@8408.4]
  assign _T_18649 = {output_24_31,output_24_30,output_24_29,output_24_28,output_24_27,output_24_26,output_24_25,output_24_24,_T_18640,_T_18633}; // @[Switch.scala 43:31:@8417.4]
  assign _T_18653 = select_0 == 5'h19; // @[Switch.scala 41:52:@8420.4]
  assign output_25_0 = io_outValid_0 & _T_18653; // @[Switch.scala 41:38:@8421.4]
  assign _T_18656 = select_1 == 5'h19; // @[Switch.scala 41:52:@8423.4]
  assign output_25_1 = io_outValid_1 & _T_18656; // @[Switch.scala 41:38:@8424.4]
  assign _T_18659 = select_2 == 5'h19; // @[Switch.scala 41:52:@8426.4]
  assign output_25_2 = io_outValid_2 & _T_18659; // @[Switch.scala 41:38:@8427.4]
  assign _T_18662 = select_3 == 5'h19; // @[Switch.scala 41:52:@8429.4]
  assign output_25_3 = io_outValid_3 & _T_18662; // @[Switch.scala 41:38:@8430.4]
  assign _T_18665 = select_4 == 5'h19; // @[Switch.scala 41:52:@8432.4]
  assign output_25_4 = io_outValid_4 & _T_18665; // @[Switch.scala 41:38:@8433.4]
  assign _T_18668 = select_5 == 5'h19; // @[Switch.scala 41:52:@8435.4]
  assign output_25_5 = io_outValid_5 & _T_18668; // @[Switch.scala 41:38:@8436.4]
  assign _T_18671 = select_6 == 5'h19; // @[Switch.scala 41:52:@8438.4]
  assign output_25_6 = io_outValid_6 & _T_18671; // @[Switch.scala 41:38:@8439.4]
  assign _T_18674 = select_7 == 5'h19; // @[Switch.scala 41:52:@8441.4]
  assign output_25_7 = io_outValid_7 & _T_18674; // @[Switch.scala 41:38:@8442.4]
  assign _T_18677 = select_8 == 5'h19; // @[Switch.scala 41:52:@8444.4]
  assign output_25_8 = io_outValid_8 & _T_18677; // @[Switch.scala 41:38:@8445.4]
  assign _T_18680 = select_9 == 5'h19; // @[Switch.scala 41:52:@8447.4]
  assign output_25_9 = io_outValid_9 & _T_18680; // @[Switch.scala 41:38:@8448.4]
  assign _T_18683 = select_10 == 5'h19; // @[Switch.scala 41:52:@8450.4]
  assign output_25_10 = io_outValid_10 & _T_18683; // @[Switch.scala 41:38:@8451.4]
  assign _T_18686 = select_11 == 5'h19; // @[Switch.scala 41:52:@8453.4]
  assign output_25_11 = io_outValid_11 & _T_18686; // @[Switch.scala 41:38:@8454.4]
  assign _T_18689 = select_12 == 5'h19; // @[Switch.scala 41:52:@8456.4]
  assign output_25_12 = io_outValid_12 & _T_18689; // @[Switch.scala 41:38:@8457.4]
  assign _T_18692 = select_13 == 5'h19; // @[Switch.scala 41:52:@8459.4]
  assign output_25_13 = io_outValid_13 & _T_18692; // @[Switch.scala 41:38:@8460.4]
  assign _T_18695 = select_14 == 5'h19; // @[Switch.scala 41:52:@8462.4]
  assign output_25_14 = io_outValid_14 & _T_18695; // @[Switch.scala 41:38:@8463.4]
  assign _T_18698 = select_15 == 5'h19; // @[Switch.scala 41:52:@8465.4]
  assign output_25_15 = io_outValid_15 & _T_18698; // @[Switch.scala 41:38:@8466.4]
  assign _T_18701 = select_16 == 5'h19; // @[Switch.scala 41:52:@8468.4]
  assign output_25_16 = io_outValid_16 & _T_18701; // @[Switch.scala 41:38:@8469.4]
  assign _T_18704 = select_17 == 5'h19; // @[Switch.scala 41:52:@8471.4]
  assign output_25_17 = io_outValid_17 & _T_18704; // @[Switch.scala 41:38:@8472.4]
  assign _T_18707 = select_18 == 5'h19; // @[Switch.scala 41:52:@8474.4]
  assign output_25_18 = io_outValid_18 & _T_18707; // @[Switch.scala 41:38:@8475.4]
  assign _T_18710 = select_19 == 5'h19; // @[Switch.scala 41:52:@8477.4]
  assign output_25_19 = io_outValid_19 & _T_18710; // @[Switch.scala 41:38:@8478.4]
  assign _T_18713 = select_20 == 5'h19; // @[Switch.scala 41:52:@8480.4]
  assign output_25_20 = io_outValid_20 & _T_18713; // @[Switch.scala 41:38:@8481.4]
  assign _T_18716 = select_21 == 5'h19; // @[Switch.scala 41:52:@8483.4]
  assign output_25_21 = io_outValid_21 & _T_18716; // @[Switch.scala 41:38:@8484.4]
  assign _T_18719 = select_22 == 5'h19; // @[Switch.scala 41:52:@8486.4]
  assign output_25_22 = io_outValid_22 & _T_18719; // @[Switch.scala 41:38:@8487.4]
  assign _T_18722 = select_23 == 5'h19; // @[Switch.scala 41:52:@8489.4]
  assign output_25_23 = io_outValid_23 & _T_18722; // @[Switch.scala 41:38:@8490.4]
  assign _T_18725 = select_24 == 5'h19; // @[Switch.scala 41:52:@8492.4]
  assign output_25_24 = io_outValid_24 & _T_18725; // @[Switch.scala 41:38:@8493.4]
  assign _T_18728 = select_25 == 5'h19; // @[Switch.scala 41:52:@8495.4]
  assign output_25_25 = io_outValid_25 & _T_18728; // @[Switch.scala 41:38:@8496.4]
  assign _T_18731 = select_26 == 5'h19; // @[Switch.scala 41:52:@8498.4]
  assign output_25_26 = io_outValid_26 & _T_18731; // @[Switch.scala 41:38:@8499.4]
  assign _T_18734 = select_27 == 5'h19; // @[Switch.scala 41:52:@8501.4]
  assign output_25_27 = io_outValid_27 & _T_18734; // @[Switch.scala 41:38:@8502.4]
  assign _T_18737 = select_28 == 5'h19; // @[Switch.scala 41:52:@8504.4]
  assign output_25_28 = io_outValid_28 & _T_18737; // @[Switch.scala 41:38:@8505.4]
  assign _T_18740 = select_29 == 5'h19; // @[Switch.scala 41:52:@8507.4]
  assign output_25_29 = io_outValid_29 & _T_18740; // @[Switch.scala 41:38:@8508.4]
  assign _T_18743 = select_30 == 5'h19; // @[Switch.scala 41:52:@8510.4]
  assign output_25_30 = io_outValid_30 & _T_18743; // @[Switch.scala 41:38:@8511.4]
  assign _T_18746 = select_31 == 5'h19; // @[Switch.scala 41:52:@8513.4]
  assign output_25_31 = io_outValid_31 & _T_18746; // @[Switch.scala 41:38:@8514.4]
  assign _T_18754 = {output_25_7,output_25_6,output_25_5,output_25_4,output_25_3,output_25_2,output_25_1,output_25_0}; // @[Switch.scala 43:31:@8522.4]
  assign _T_18762 = {output_25_15,output_25_14,output_25_13,output_25_12,output_25_11,output_25_10,output_25_9,output_25_8,_T_18754}; // @[Switch.scala 43:31:@8530.4]
  assign _T_18769 = {output_25_23,output_25_22,output_25_21,output_25_20,output_25_19,output_25_18,output_25_17,output_25_16}; // @[Switch.scala 43:31:@8537.4]
  assign _T_18778 = {output_25_31,output_25_30,output_25_29,output_25_28,output_25_27,output_25_26,output_25_25,output_25_24,_T_18769,_T_18762}; // @[Switch.scala 43:31:@8546.4]
  assign _T_18782 = select_0 == 5'h1a; // @[Switch.scala 41:52:@8549.4]
  assign output_26_0 = io_outValid_0 & _T_18782; // @[Switch.scala 41:38:@8550.4]
  assign _T_18785 = select_1 == 5'h1a; // @[Switch.scala 41:52:@8552.4]
  assign output_26_1 = io_outValid_1 & _T_18785; // @[Switch.scala 41:38:@8553.4]
  assign _T_18788 = select_2 == 5'h1a; // @[Switch.scala 41:52:@8555.4]
  assign output_26_2 = io_outValid_2 & _T_18788; // @[Switch.scala 41:38:@8556.4]
  assign _T_18791 = select_3 == 5'h1a; // @[Switch.scala 41:52:@8558.4]
  assign output_26_3 = io_outValid_3 & _T_18791; // @[Switch.scala 41:38:@8559.4]
  assign _T_18794 = select_4 == 5'h1a; // @[Switch.scala 41:52:@8561.4]
  assign output_26_4 = io_outValid_4 & _T_18794; // @[Switch.scala 41:38:@8562.4]
  assign _T_18797 = select_5 == 5'h1a; // @[Switch.scala 41:52:@8564.4]
  assign output_26_5 = io_outValid_5 & _T_18797; // @[Switch.scala 41:38:@8565.4]
  assign _T_18800 = select_6 == 5'h1a; // @[Switch.scala 41:52:@8567.4]
  assign output_26_6 = io_outValid_6 & _T_18800; // @[Switch.scala 41:38:@8568.4]
  assign _T_18803 = select_7 == 5'h1a; // @[Switch.scala 41:52:@8570.4]
  assign output_26_7 = io_outValid_7 & _T_18803; // @[Switch.scala 41:38:@8571.4]
  assign _T_18806 = select_8 == 5'h1a; // @[Switch.scala 41:52:@8573.4]
  assign output_26_8 = io_outValid_8 & _T_18806; // @[Switch.scala 41:38:@8574.4]
  assign _T_18809 = select_9 == 5'h1a; // @[Switch.scala 41:52:@8576.4]
  assign output_26_9 = io_outValid_9 & _T_18809; // @[Switch.scala 41:38:@8577.4]
  assign _T_18812 = select_10 == 5'h1a; // @[Switch.scala 41:52:@8579.4]
  assign output_26_10 = io_outValid_10 & _T_18812; // @[Switch.scala 41:38:@8580.4]
  assign _T_18815 = select_11 == 5'h1a; // @[Switch.scala 41:52:@8582.4]
  assign output_26_11 = io_outValid_11 & _T_18815; // @[Switch.scala 41:38:@8583.4]
  assign _T_18818 = select_12 == 5'h1a; // @[Switch.scala 41:52:@8585.4]
  assign output_26_12 = io_outValid_12 & _T_18818; // @[Switch.scala 41:38:@8586.4]
  assign _T_18821 = select_13 == 5'h1a; // @[Switch.scala 41:52:@8588.4]
  assign output_26_13 = io_outValid_13 & _T_18821; // @[Switch.scala 41:38:@8589.4]
  assign _T_18824 = select_14 == 5'h1a; // @[Switch.scala 41:52:@8591.4]
  assign output_26_14 = io_outValid_14 & _T_18824; // @[Switch.scala 41:38:@8592.4]
  assign _T_18827 = select_15 == 5'h1a; // @[Switch.scala 41:52:@8594.4]
  assign output_26_15 = io_outValid_15 & _T_18827; // @[Switch.scala 41:38:@8595.4]
  assign _T_18830 = select_16 == 5'h1a; // @[Switch.scala 41:52:@8597.4]
  assign output_26_16 = io_outValid_16 & _T_18830; // @[Switch.scala 41:38:@8598.4]
  assign _T_18833 = select_17 == 5'h1a; // @[Switch.scala 41:52:@8600.4]
  assign output_26_17 = io_outValid_17 & _T_18833; // @[Switch.scala 41:38:@8601.4]
  assign _T_18836 = select_18 == 5'h1a; // @[Switch.scala 41:52:@8603.4]
  assign output_26_18 = io_outValid_18 & _T_18836; // @[Switch.scala 41:38:@8604.4]
  assign _T_18839 = select_19 == 5'h1a; // @[Switch.scala 41:52:@8606.4]
  assign output_26_19 = io_outValid_19 & _T_18839; // @[Switch.scala 41:38:@8607.4]
  assign _T_18842 = select_20 == 5'h1a; // @[Switch.scala 41:52:@8609.4]
  assign output_26_20 = io_outValid_20 & _T_18842; // @[Switch.scala 41:38:@8610.4]
  assign _T_18845 = select_21 == 5'h1a; // @[Switch.scala 41:52:@8612.4]
  assign output_26_21 = io_outValid_21 & _T_18845; // @[Switch.scala 41:38:@8613.4]
  assign _T_18848 = select_22 == 5'h1a; // @[Switch.scala 41:52:@8615.4]
  assign output_26_22 = io_outValid_22 & _T_18848; // @[Switch.scala 41:38:@8616.4]
  assign _T_18851 = select_23 == 5'h1a; // @[Switch.scala 41:52:@8618.4]
  assign output_26_23 = io_outValid_23 & _T_18851; // @[Switch.scala 41:38:@8619.4]
  assign _T_18854 = select_24 == 5'h1a; // @[Switch.scala 41:52:@8621.4]
  assign output_26_24 = io_outValid_24 & _T_18854; // @[Switch.scala 41:38:@8622.4]
  assign _T_18857 = select_25 == 5'h1a; // @[Switch.scala 41:52:@8624.4]
  assign output_26_25 = io_outValid_25 & _T_18857; // @[Switch.scala 41:38:@8625.4]
  assign _T_18860 = select_26 == 5'h1a; // @[Switch.scala 41:52:@8627.4]
  assign output_26_26 = io_outValid_26 & _T_18860; // @[Switch.scala 41:38:@8628.4]
  assign _T_18863 = select_27 == 5'h1a; // @[Switch.scala 41:52:@8630.4]
  assign output_26_27 = io_outValid_27 & _T_18863; // @[Switch.scala 41:38:@8631.4]
  assign _T_18866 = select_28 == 5'h1a; // @[Switch.scala 41:52:@8633.4]
  assign output_26_28 = io_outValid_28 & _T_18866; // @[Switch.scala 41:38:@8634.4]
  assign _T_18869 = select_29 == 5'h1a; // @[Switch.scala 41:52:@8636.4]
  assign output_26_29 = io_outValid_29 & _T_18869; // @[Switch.scala 41:38:@8637.4]
  assign _T_18872 = select_30 == 5'h1a; // @[Switch.scala 41:52:@8639.4]
  assign output_26_30 = io_outValid_30 & _T_18872; // @[Switch.scala 41:38:@8640.4]
  assign _T_18875 = select_31 == 5'h1a; // @[Switch.scala 41:52:@8642.4]
  assign output_26_31 = io_outValid_31 & _T_18875; // @[Switch.scala 41:38:@8643.4]
  assign _T_18883 = {output_26_7,output_26_6,output_26_5,output_26_4,output_26_3,output_26_2,output_26_1,output_26_0}; // @[Switch.scala 43:31:@8651.4]
  assign _T_18891 = {output_26_15,output_26_14,output_26_13,output_26_12,output_26_11,output_26_10,output_26_9,output_26_8,_T_18883}; // @[Switch.scala 43:31:@8659.4]
  assign _T_18898 = {output_26_23,output_26_22,output_26_21,output_26_20,output_26_19,output_26_18,output_26_17,output_26_16}; // @[Switch.scala 43:31:@8666.4]
  assign _T_18907 = {output_26_31,output_26_30,output_26_29,output_26_28,output_26_27,output_26_26,output_26_25,output_26_24,_T_18898,_T_18891}; // @[Switch.scala 43:31:@8675.4]
  assign _T_18911 = select_0 == 5'h1b; // @[Switch.scala 41:52:@8678.4]
  assign output_27_0 = io_outValid_0 & _T_18911; // @[Switch.scala 41:38:@8679.4]
  assign _T_18914 = select_1 == 5'h1b; // @[Switch.scala 41:52:@8681.4]
  assign output_27_1 = io_outValid_1 & _T_18914; // @[Switch.scala 41:38:@8682.4]
  assign _T_18917 = select_2 == 5'h1b; // @[Switch.scala 41:52:@8684.4]
  assign output_27_2 = io_outValid_2 & _T_18917; // @[Switch.scala 41:38:@8685.4]
  assign _T_18920 = select_3 == 5'h1b; // @[Switch.scala 41:52:@8687.4]
  assign output_27_3 = io_outValid_3 & _T_18920; // @[Switch.scala 41:38:@8688.4]
  assign _T_18923 = select_4 == 5'h1b; // @[Switch.scala 41:52:@8690.4]
  assign output_27_4 = io_outValid_4 & _T_18923; // @[Switch.scala 41:38:@8691.4]
  assign _T_18926 = select_5 == 5'h1b; // @[Switch.scala 41:52:@8693.4]
  assign output_27_5 = io_outValid_5 & _T_18926; // @[Switch.scala 41:38:@8694.4]
  assign _T_18929 = select_6 == 5'h1b; // @[Switch.scala 41:52:@8696.4]
  assign output_27_6 = io_outValid_6 & _T_18929; // @[Switch.scala 41:38:@8697.4]
  assign _T_18932 = select_7 == 5'h1b; // @[Switch.scala 41:52:@8699.4]
  assign output_27_7 = io_outValid_7 & _T_18932; // @[Switch.scala 41:38:@8700.4]
  assign _T_18935 = select_8 == 5'h1b; // @[Switch.scala 41:52:@8702.4]
  assign output_27_8 = io_outValid_8 & _T_18935; // @[Switch.scala 41:38:@8703.4]
  assign _T_18938 = select_9 == 5'h1b; // @[Switch.scala 41:52:@8705.4]
  assign output_27_9 = io_outValid_9 & _T_18938; // @[Switch.scala 41:38:@8706.4]
  assign _T_18941 = select_10 == 5'h1b; // @[Switch.scala 41:52:@8708.4]
  assign output_27_10 = io_outValid_10 & _T_18941; // @[Switch.scala 41:38:@8709.4]
  assign _T_18944 = select_11 == 5'h1b; // @[Switch.scala 41:52:@8711.4]
  assign output_27_11 = io_outValid_11 & _T_18944; // @[Switch.scala 41:38:@8712.4]
  assign _T_18947 = select_12 == 5'h1b; // @[Switch.scala 41:52:@8714.4]
  assign output_27_12 = io_outValid_12 & _T_18947; // @[Switch.scala 41:38:@8715.4]
  assign _T_18950 = select_13 == 5'h1b; // @[Switch.scala 41:52:@8717.4]
  assign output_27_13 = io_outValid_13 & _T_18950; // @[Switch.scala 41:38:@8718.4]
  assign _T_18953 = select_14 == 5'h1b; // @[Switch.scala 41:52:@8720.4]
  assign output_27_14 = io_outValid_14 & _T_18953; // @[Switch.scala 41:38:@8721.4]
  assign _T_18956 = select_15 == 5'h1b; // @[Switch.scala 41:52:@8723.4]
  assign output_27_15 = io_outValid_15 & _T_18956; // @[Switch.scala 41:38:@8724.4]
  assign _T_18959 = select_16 == 5'h1b; // @[Switch.scala 41:52:@8726.4]
  assign output_27_16 = io_outValid_16 & _T_18959; // @[Switch.scala 41:38:@8727.4]
  assign _T_18962 = select_17 == 5'h1b; // @[Switch.scala 41:52:@8729.4]
  assign output_27_17 = io_outValid_17 & _T_18962; // @[Switch.scala 41:38:@8730.4]
  assign _T_18965 = select_18 == 5'h1b; // @[Switch.scala 41:52:@8732.4]
  assign output_27_18 = io_outValid_18 & _T_18965; // @[Switch.scala 41:38:@8733.4]
  assign _T_18968 = select_19 == 5'h1b; // @[Switch.scala 41:52:@8735.4]
  assign output_27_19 = io_outValid_19 & _T_18968; // @[Switch.scala 41:38:@8736.4]
  assign _T_18971 = select_20 == 5'h1b; // @[Switch.scala 41:52:@8738.4]
  assign output_27_20 = io_outValid_20 & _T_18971; // @[Switch.scala 41:38:@8739.4]
  assign _T_18974 = select_21 == 5'h1b; // @[Switch.scala 41:52:@8741.4]
  assign output_27_21 = io_outValid_21 & _T_18974; // @[Switch.scala 41:38:@8742.4]
  assign _T_18977 = select_22 == 5'h1b; // @[Switch.scala 41:52:@8744.4]
  assign output_27_22 = io_outValid_22 & _T_18977; // @[Switch.scala 41:38:@8745.4]
  assign _T_18980 = select_23 == 5'h1b; // @[Switch.scala 41:52:@8747.4]
  assign output_27_23 = io_outValid_23 & _T_18980; // @[Switch.scala 41:38:@8748.4]
  assign _T_18983 = select_24 == 5'h1b; // @[Switch.scala 41:52:@8750.4]
  assign output_27_24 = io_outValid_24 & _T_18983; // @[Switch.scala 41:38:@8751.4]
  assign _T_18986 = select_25 == 5'h1b; // @[Switch.scala 41:52:@8753.4]
  assign output_27_25 = io_outValid_25 & _T_18986; // @[Switch.scala 41:38:@8754.4]
  assign _T_18989 = select_26 == 5'h1b; // @[Switch.scala 41:52:@8756.4]
  assign output_27_26 = io_outValid_26 & _T_18989; // @[Switch.scala 41:38:@8757.4]
  assign _T_18992 = select_27 == 5'h1b; // @[Switch.scala 41:52:@8759.4]
  assign output_27_27 = io_outValid_27 & _T_18992; // @[Switch.scala 41:38:@8760.4]
  assign _T_18995 = select_28 == 5'h1b; // @[Switch.scala 41:52:@8762.4]
  assign output_27_28 = io_outValid_28 & _T_18995; // @[Switch.scala 41:38:@8763.4]
  assign _T_18998 = select_29 == 5'h1b; // @[Switch.scala 41:52:@8765.4]
  assign output_27_29 = io_outValid_29 & _T_18998; // @[Switch.scala 41:38:@8766.4]
  assign _T_19001 = select_30 == 5'h1b; // @[Switch.scala 41:52:@8768.4]
  assign output_27_30 = io_outValid_30 & _T_19001; // @[Switch.scala 41:38:@8769.4]
  assign _T_19004 = select_31 == 5'h1b; // @[Switch.scala 41:52:@8771.4]
  assign output_27_31 = io_outValid_31 & _T_19004; // @[Switch.scala 41:38:@8772.4]
  assign _T_19012 = {output_27_7,output_27_6,output_27_5,output_27_4,output_27_3,output_27_2,output_27_1,output_27_0}; // @[Switch.scala 43:31:@8780.4]
  assign _T_19020 = {output_27_15,output_27_14,output_27_13,output_27_12,output_27_11,output_27_10,output_27_9,output_27_8,_T_19012}; // @[Switch.scala 43:31:@8788.4]
  assign _T_19027 = {output_27_23,output_27_22,output_27_21,output_27_20,output_27_19,output_27_18,output_27_17,output_27_16}; // @[Switch.scala 43:31:@8795.4]
  assign _T_19036 = {output_27_31,output_27_30,output_27_29,output_27_28,output_27_27,output_27_26,output_27_25,output_27_24,_T_19027,_T_19020}; // @[Switch.scala 43:31:@8804.4]
  assign _T_19040 = select_0 == 5'h1c; // @[Switch.scala 41:52:@8807.4]
  assign output_28_0 = io_outValid_0 & _T_19040; // @[Switch.scala 41:38:@8808.4]
  assign _T_19043 = select_1 == 5'h1c; // @[Switch.scala 41:52:@8810.4]
  assign output_28_1 = io_outValid_1 & _T_19043; // @[Switch.scala 41:38:@8811.4]
  assign _T_19046 = select_2 == 5'h1c; // @[Switch.scala 41:52:@8813.4]
  assign output_28_2 = io_outValid_2 & _T_19046; // @[Switch.scala 41:38:@8814.4]
  assign _T_19049 = select_3 == 5'h1c; // @[Switch.scala 41:52:@8816.4]
  assign output_28_3 = io_outValid_3 & _T_19049; // @[Switch.scala 41:38:@8817.4]
  assign _T_19052 = select_4 == 5'h1c; // @[Switch.scala 41:52:@8819.4]
  assign output_28_4 = io_outValid_4 & _T_19052; // @[Switch.scala 41:38:@8820.4]
  assign _T_19055 = select_5 == 5'h1c; // @[Switch.scala 41:52:@8822.4]
  assign output_28_5 = io_outValid_5 & _T_19055; // @[Switch.scala 41:38:@8823.4]
  assign _T_19058 = select_6 == 5'h1c; // @[Switch.scala 41:52:@8825.4]
  assign output_28_6 = io_outValid_6 & _T_19058; // @[Switch.scala 41:38:@8826.4]
  assign _T_19061 = select_7 == 5'h1c; // @[Switch.scala 41:52:@8828.4]
  assign output_28_7 = io_outValid_7 & _T_19061; // @[Switch.scala 41:38:@8829.4]
  assign _T_19064 = select_8 == 5'h1c; // @[Switch.scala 41:52:@8831.4]
  assign output_28_8 = io_outValid_8 & _T_19064; // @[Switch.scala 41:38:@8832.4]
  assign _T_19067 = select_9 == 5'h1c; // @[Switch.scala 41:52:@8834.4]
  assign output_28_9 = io_outValid_9 & _T_19067; // @[Switch.scala 41:38:@8835.4]
  assign _T_19070 = select_10 == 5'h1c; // @[Switch.scala 41:52:@8837.4]
  assign output_28_10 = io_outValid_10 & _T_19070; // @[Switch.scala 41:38:@8838.4]
  assign _T_19073 = select_11 == 5'h1c; // @[Switch.scala 41:52:@8840.4]
  assign output_28_11 = io_outValid_11 & _T_19073; // @[Switch.scala 41:38:@8841.4]
  assign _T_19076 = select_12 == 5'h1c; // @[Switch.scala 41:52:@8843.4]
  assign output_28_12 = io_outValid_12 & _T_19076; // @[Switch.scala 41:38:@8844.4]
  assign _T_19079 = select_13 == 5'h1c; // @[Switch.scala 41:52:@8846.4]
  assign output_28_13 = io_outValid_13 & _T_19079; // @[Switch.scala 41:38:@8847.4]
  assign _T_19082 = select_14 == 5'h1c; // @[Switch.scala 41:52:@8849.4]
  assign output_28_14 = io_outValid_14 & _T_19082; // @[Switch.scala 41:38:@8850.4]
  assign _T_19085 = select_15 == 5'h1c; // @[Switch.scala 41:52:@8852.4]
  assign output_28_15 = io_outValid_15 & _T_19085; // @[Switch.scala 41:38:@8853.4]
  assign _T_19088 = select_16 == 5'h1c; // @[Switch.scala 41:52:@8855.4]
  assign output_28_16 = io_outValid_16 & _T_19088; // @[Switch.scala 41:38:@8856.4]
  assign _T_19091 = select_17 == 5'h1c; // @[Switch.scala 41:52:@8858.4]
  assign output_28_17 = io_outValid_17 & _T_19091; // @[Switch.scala 41:38:@8859.4]
  assign _T_19094 = select_18 == 5'h1c; // @[Switch.scala 41:52:@8861.4]
  assign output_28_18 = io_outValid_18 & _T_19094; // @[Switch.scala 41:38:@8862.4]
  assign _T_19097 = select_19 == 5'h1c; // @[Switch.scala 41:52:@8864.4]
  assign output_28_19 = io_outValid_19 & _T_19097; // @[Switch.scala 41:38:@8865.4]
  assign _T_19100 = select_20 == 5'h1c; // @[Switch.scala 41:52:@8867.4]
  assign output_28_20 = io_outValid_20 & _T_19100; // @[Switch.scala 41:38:@8868.4]
  assign _T_19103 = select_21 == 5'h1c; // @[Switch.scala 41:52:@8870.4]
  assign output_28_21 = io_outValid_21 & _T_19103; // @[Switch.scala 41:38:@8871.4]
  assign _T_19106 = select_22 == 5'h1c; // @[Switch.scala 41:52:@8873.4]
  assign output_28_22 = io_outValid_22 & _T_19106; // @[Switch.scala 41:38:@8874.4]
  assign _T_19109 = select_23 == 5'h1c; // @[Switch.scala 41:52:@8876.4]
  assign output_28_23 = io_outValid_23 & _T_19109; // @[Switch.scala 41:38:@8877.4]
  assign _T_19112 = select_24 == 5'h1c; // @[Switch.scala 41:52:@8879.4]
  assign output_28_24 = io_outValid_24 & _T_19112; // @[Switch.scala 41:38:@8880.4]
  assign _T_19115 = select_25 == 5'h1c; // @[Switch.scala 41:52:@8882.4]
  assign output_28_25 = io_outValid_25 & _T_19115; // @[Switch.scala 41:38:@8883.4]
  assign _T_19118 = select_26 == 5'h1c; // @[Switch.scala 41:52:@8885.4]
  assign output_28_26 = io_outValid_26 & _T_19118; // @[Switch.scala 41:38:@8886.4]
  assign _T_19121 = select_27 == 5'h1c; // @[Switch.scala 41:52:@8888.4]
  assign output_28_27 = io_outValid_27 & _T_19121; // @[Switch.scala 41:38:@8889.4]
  assign _T_19124 = select_28 == 5'h1c; // @[Switch.scala 41:52:@8891.4]
  assign output_28_28 = io_outValid_28 & _T_19124; // @[Switch.scala 41:38:@8892.4]
  assign _T_19127 = select_29 == 5'h1c; // @[Switch.scala 41:52:@8894.4]
  assign output_28_29 = io_outValid_29 & _T_19127; // @[Switch.scala 41:38:@8895.4]
  assign _T_19130 = select_30 == 5'h1c; // @[Switch.scala 41:52:@8897.4]
  assign output_28_30 = io_outValid_30 & _T_19130; // @[Switch.scala 41:38:@8898.4]
  assign _T_19133 = select_31 == 5'h1c; // @[Switch.scala 41:52:@8900.4]
  assign output_28_31 = io_outValid_31 & _T_19133; // @[Switch.scala 41:38:@8901.4]
  assign _T_19141 = {output_28_7,output_28_6,output_28_5,output_28_4,output_28_3,output_28_2,output_28_1,output_28_0}; // @[Switch.scala 43:31:@8909.4]
  assign _T_19149 = {output_28_15,output_28_14,output_28_13,output_28_12,output_28_11,output_28_10,output_28_9,output_28_8,_T_19141}; // @[Switch.scala 43:31:@8917.4]
  assign _T_19156 = {output_28_23,output_28_22,output_28_21,output_28_20,output_28_19,output_28_18,output_28_17,output_28_16}; // @[Switch.scala 43:31:@8924.4]
  assign _T_19165 = {output_28_31,output_28_30,output_28_29,output_28_28,output_28_27,output_28_26,output_28_25,output_28_24,_T_19156,_T_19149}; // @[Switch.scala 43:31:@8933.4]
  assign _T_19169 = select_0 == 5'h1d; // @[Switch.scala 41:52:@8936.4]
  assign output_29_0 = io_outValid_0 & _T_19169; // @[Switch.scala 41:38:@8937.4]
  assign _T_19172 = select_1 == 5'h1d; // @[Switch.scala 41:52:@8939.4]
  assign output_29_1 = io_outValid_1 & _T_19172; // @[Switch.scala 41:38:@8940.4]
  assign _T_19175 = select_2 == 5'h1d; // @[Switch.scala 41:52:@8942.4]
  assign output_29_2 = io_outValid_2 & _T_19175; // @[Switch.scala 41:38:@8943.4]
  assign _T_19178 = select_3 == 5'h1d; // @[Switch.scala 41:52:@8945.4]
  assign output_29_3 = io_outValid_3 & _T_19178; // @[Switch.scala 41:38:@8946.4]
  assign _T_19181 = select_4 == 5'h1d; // @[Switch.scala 41:52:@8948.4]
  assign output_29_4 = io_outValid_4 & _T_19181; // @[Switch.scala 41:38:@8949.4]
  assign _T_19184 = select_5 == 5'h1d; // @[Switch.scala 41:52:@8951.4]
  assign output_29_5 = io_outValid_5 & _T_19184; // @[Switch.scala 41:38:@8952.4]
  assign _T_19187 = select_6 == 5'h1d; // @[Switch.scala 41:52:@8954.4]
  assign output_29_6 = io_outValid_6 & _T_19187; // @[Switch.scala 41:38:@8955.4]
  assign _T_19190 = select_7 == 5'h1d; // @[Switch.scala 41:52:@8957.4]
  assign output_29_7 = io_outValid_7 & _T_19190; // @[Switch.scala 41:38:@8958.4]
  assign _T_19193 = select_8 == 5'h1d; // @[Switch.scala 41:52:@8960.4]
  assign output_29_8 = io_outValid_8 & _T_19193; // @[Switch.scala 41:38:@8961.4]
  assign _T_19196 = select_9 == 5'h1d; // @[Switch.scala 41:52:@8963.4]
  assign output_29_9 = io_outValid_9 & _T_19196; // @[Switch.scala 41:38:@8964.4]
  assign _T_19199 = select_10 == 5'h1d; // @[Switch.scala 41:52:@8966.4]
  assign output_29_10 = io_outValid_10 & _T_19199; // @[Switch.scala 41:38:@8967.4]
  assign _T_19202 = select_11 == 5'h1d; // @[Switch.scala 41:52:@8969.4]
  assign output_29_11 = io_outValid_11 & _T_19202; // @[Switch.scala 41:38:@8970.4]
  assign _T_19205 = select_12 == 5'h1d; // @[Switch.scala 41:52:@8972.4]
  assign output_29_12 = io_outValid_12 & _T_19205; // @[Switch.scala 41:38:@8973.4]
  assign _T_19208 = select_13 == 5'h1d; // @[Switch.scala 41:52:@8975.4]
  assign output_29_13 = io_outValid_13 & _T_19208; // @[Switch.scala 41:38:@8976.4]
  assign _T_19211 = select_14 == 5'h1d; // @[Switch.scala 41:52:@8978.4]
  assign output_29_14 = io_outValid_14 & _T_19211; // @[Switch.scala 41:38:@8979.4]
  assign _T_19214 = select_15 == 5'h1d; // @[Switch.scala 41:52:@8981.4]
  assign output_29_15 = io_outValid_15 & _T_19214; // @[Switch.scala 41:38:@8982.4]
  assign _T_19217 = select_16 == 5'h1d; // @[Switch.scala 41:52:@8984.4]
  assign output_29_16 = io_outValid_16 & _T_19217; // @[Switch.scala 41:38:@8985.4]
  assign _T_19220 = select_17 == 5'h1d; // @[Switch.scala 41:52:@8987.4]
  assign output_29_17 = io_outValid_17 & _T_19220; // @[Switch.scala 41:38:@8988.4]
  assign _T_19223 = select_18 == 5'h1d; // @[Switch.scala 41:52:@8990.4]
  assign output_29_18 = io_outValid_18 & _T_19223; // @[Switch.scala 41:38:@8991.4]
  assign _T_19226 = select_19 == 5'h1d; // @[Switch.scala 41:52:@8993.4]
  assign output_29_19 = io_outValid_19 & _T_19226; // @[Switch.scala 41:38:@8994.4]
  assign _T_19229 = select_20 == 5'h1d; // @[Switch.scala 41:52:@8996.4]
  assign output_29_20 = io_outValid_20 & _T_19229; // @[Switch.scala 41:38:@8997.4]
  assign _T_19232 = select_21 == 5'h1d; // @[Switch.scala 41:52:@8999.4]
  assign output_29_21 = io_outValid_21 & _T_19232; // @[Switch.scala 41:38:@9000.4]
  assign _T_19235 = select_22 == 5'h1d; // @[Switch.scala 41:52:@9002.4]
  assign output_29_22 = io_outValid_22 & _T_19235; // @[Switch.scala 41:38:@9003.4]
  assign _T_19238 = select_23 == 5'h1d; // @[Switch.scala 41:52:@9005.4]
  assign output_29_23 = io_outValid_23 & _T_19238; // @[Switch.scala 41:38:@9006.4]
  assign _T_19241 = select_24 == 5'h1d; // @[Switch.scala 41:52:@9008.4]
  assign output_29_24 = io_outValid_24 & _T_19241; // @[Switch.scala 41:38:@9009.4]
  assign _T_19244 = select_25 == 5'h1d; // @[Switch.scala 41:52:@9011.4]
  assign output_29_25 = io_outValid_25 & _T_19244; // @[Switch.scala 41:38:@9012.4]
  assign _T_19247 = select_26 == 5'h1d; // @[Switch.scala 41:52:@9014.4]
  assign output_29_26 = io_outValid_26 & _T_19247; // @[Switch.scala 41:38:@9015.4]
  assign _T_19250 = select_27 == 5'h1d; // @[Switch.scala 41:52:@9017.4]
  assign output_29_27 = io_outValid_27 & _T_19250; // @[Switch.scala 41:38:@9018.4]
  assign _T_19253 = select_28 == 5'h1d; // @[Switch.scala 41:52:@9020.4]
  assign output_29_28 = io_outValid_28 & _T_19253; // @[Switch.scala 41:38:@9021.4]
  assign _T_19256 = select_29 == 5'h1d; // @[Switch.scala 41:52:@9023.4]
  assign output_29_29 = io_outValid_29 & _T_19256; // @[Switch.scala 41:38:@9024.4]
  assign _T_19259 = select_30 == 5'h1d; // @[Switch.scala 41:52:@9026.4]
  assign output_29_30 = io_outValid_30 & _T_19259; // @[Switch.scala 41:38:@9027.4]
  assign _T_19262 = select_31 == 5'h1d; // @[Switch.scala 41:52:@9029.4]
  assign output_29_31 = io_outValid_31 & _T_19262; // @[Switch.scala 41:38:@9030.4]
  assign _T_19270 = {output_29_7,output_29_6,output_29_5,output_29_4,output_29_3,output_29_2,output_29_1,output_29_0}; // @[Switch.scala 43:31:@9038.4]
  assign _T_19278 = {output_29_15,output_29_14,output_29_13,output_29_12,output_29_11,output_29_10,output_29_9,output_29_8,_T_19270}; // @[Switch.scala 43:31:@9046.4]
  assign _T_19285 = {output_29_23,output_29_22,output_29_21,output_29_20,output_29_19,output_29_18,output_29_17,output_29_16}; // @[Switch.scala 43:31:@9053.4]
  assign _T_19294 = {output_29_31,output_29_30,output_29_29,output_29_28,output_29_27,output_29_26,output_29_25,output_29_24,_T_19285,_T_19278}; // @[Switch.scala 43:31:@9062.4]
  assign _T_19298 = select_0 == 5'h1e; // @[Switch.scala 41:52:@9065.4]
  assign output_30_0 = io_outValid_0 & _T_19298; // @[Switch.scala 41:38:@9066.4]
  assign _T_19301 = select_1 == 5'h1e; // @[Switch.scala 41:52:@9068.4]
  assign output_30_1 = io_outValid_1 & _T_19301; // @[Switch.scala 41:38:@9069.4]
  assign _T_19304 = select_2 == 5'h1e; // @[Switch.scala 41:52:@9071.4]
  assign output_30_2 = io_outValid_2 & _T_19304; // @[Switch.scala 41:38:@9072.4]
  assign _T_19307 = select_3 == 5'h1e; // @[Switch.scala 41:52:@9074.4]
  assign output_30_3 = io_outValid_3 & _T_19307; // @[Switch.scala 41:38:@9075.4]
  assign _T_19310 = select_4 == 5'h1e; // @[Switch.scala 41:52:@9077.4]
  assign output_30_4 = io_outValid_4 & _T_19310; // @[Switch.scala 41:38:@9078.4]
  assign _T_19313 = select_5 == 5'h1e; // @[Switch.scala 41:52:@9080.4]
  assign output_30_5 = io_outValid_5 & _T_19313; // @[Switch.scala 41:38:@9081.4]
  assign _T_19316 = select_6 == 5'h1e; // @[Switch.scala 41:52:@9083.4]
  assign output_30_6 = io_outValid_6 & _T_19316; // @[Switch.scala 41:38:@9084.4]
  assign _T_19319 = select_7 == 5'h1e; // @[Switch.scala 41:52:@9086.4]
  assign output_30_7 = io_outValid_7 & _T_19319; // @[Switch.scala 41:38:@9087.4]
  assign _T_19322 = select_8 == 5'h1e; // @[Switch.scala 41:52:@9089.4]
  assign output_30_8 = io_outValid_8 & _T_19322; // @[Switch.scala 41:38:@9090.4]
  assign _T_19325 = select_9 == 5'h1e; // @[Switch.scala 41:52:@9092.4]
  assign output_30_9 = io_outValid_9 & _T_19325; // @[Switch.scala 41:38:@9093.4]
  assign _T_19328 = select_10 == 5'h1e; // @[Switch.scala 41:52:@9095.4]
  assign output_30_10 = io_outValid_10 & _T_19328; // @[Switch.scala 41:38:@9096.4]
  assign _T_19331 = select_11 == 5'h1e; // @[Switch.scala 41:52:@9098.4]
  assign output_30_11 = io_outValid_11 & _T_19331; // @[Switch.scala 41:38:@9099.4]
  assign _T_19334 = select_12 == 5'h1e; // @[Switch.scala 41:52:@9101.4]
  assign output_30_12 = io_outValid_12 & _T_19334; // @[Switch.scala 41:38:@9102.4]
  assign _T_19337 = select_13 == 5'h1e; // @[Switch.scala 41:52:@9104.4]
  assign output_30_13 = io_outValid_13 & _T_19337; // @[Switch.scala 41:38:@9105.4]
  assign _T_19340 = select_14 == 5'h1e; // @[Switch.scala 41:52:@9107.4]
  assign output_30_14 = io_outValid_14 & _T_19340; // @[Switch.scala 41:38:@9108.4]
  assign _T_19343 = select_15 == 5'h1e; // @[Switch.scala 41:52:@9110.4]
  assign output_30_15 = io_outValid_15 & _T_19343; // @[Switch.scala 41:38:@9111.4]
  assign _T_19346 = select_16 == 5'h1e; // @[Switch.scala 41:52:@9113.4]
  assign output_30_16 = io_outValid_16 & _T_19346; // @[Switch.scala 41:38:@9114.4]
  assign _T_19349 = select_17 == 5'h1e; // @[Switch.scala 41:52:@9116.4]
  assign output_30_17 = io_outValid_17 & _T_19349; // @[Switch.scala 41:38:@9117.4]
  assign _T_19352 = select_18 == 5'h1e; // @[Switch.scala 41:52:@9119.4]
  assign output_30_18 = io_outValid_18 & _T_19352; // @[Switch.scala 41:38:@9120.4]
  assign _T_19355 = select_19 == 5'h1e; // @[Switch.scala 41:52:@9122.4]
  assign output_30_19 = io_outValid_19 & _T_19355; // @[Switch.scala 41:38:@9123.4]
  assign _T_19358 = select_20 == 5'h1e; // @[Switch.scala 41:52:@9125.4]
  assign output_30_20 = io_outValid_20 & _T_19358; // @[Switch.scala 41:38:@9126.4]
  assign _T_19361 = select_21 == 5'h1e; // @[Switch.scala 41:52:@9128.4]
  assign output_30_21 = io_outValid_21 & _T_19361; // @[Switch.scala 41:38:@9129.4]
  assign _T_19364 = select_22 == 5'h1e; // @[Switch.scala 41:52:@9131.4]
  assign output_30_22 = io_outValid_22 & _T_19364; // @[Switch.scala 41:38:@9132.4]
  assign _T_19367 = select_23 == 5'h1e; // @[Switch.scala 41:52:@9134.4]
  assign output_30_23 = io_outValid_23 & _T_19367; // @[Switch.scala 41:38:@9135.4]
  assign _T_19370 = select_24 == 5'h1e; // @[Switch.scala 41:52:@9137.4]
  assign output_30_24 = io_outValid_24 & _T_19370; // @[Switch.scala 41:38:@9138.4]
  assign _T_19373 = select_25 == 5'h1e; // @[Switch.scala 41:52:@9140.4]
  assign output_30_25 = io_outValid_25 & _T_19373; // @[Switch.scala 41:38:@9141.4]
  assign _T_19376 = select_26 == 5'h1e; // @[Switch.scala 41:52:@9143.4]
  assign output_30_26 = io_outValid_26 & _T_19376; // @[Switch.scala 41:38:@9144.4]
  assign _T_19379 = select_27 == 5'h1e; // @[Switch.scala 41:52:@9146.4]
  assign output_30_27 = io_outValid_27 & _T_19379; // @[Switch.scala 41:38:@9147.4]
  assign _T_19382 = select_28 == 5'h1e; // @[Switch.scala 41:52:@9149.4]
  assign output_30_28 = io_outValid_28 & _T_19382; // @[Switch.scala 41:38:@9150.4]
  assign _T_19385 = select_29 == 5'h1e; // @[Switch.scala 41:52:@9152.4]
  assign output_30_29 = io_outValid_29 & _T_19385; // @[Switch.scala 41:38:@9153.4]
  assign _T_19388 = select_30 == 5'h1e; // @[Switch.scala 41:52:@9155.4]
  assign output_30_30 = io_outValid_30 & _T_19388; // @[Switch.scala 41:38:@9156.4]
  assign _T_19391 = select_31 == 5'h1e; // @[Switch.scala 41:52:@9158.4]
  assign output_30_31 = io_outValid_31 & _T_19391; // @[Switch.scala 41:38:@9159.4]
  assign _T_19399 = {output_30_7,output_30_6,output_30_5,output_30_4,output_30_3,output_30_2,output_30_1,output_30_0}; // @[Switch.scala 43:31:@9167.4]
  assign _T_19407 = {output_30_15,output_30_14,output_30_13,output_30_12,output_30_11,output_30_10,output_30_9,output_30_8,_T_19399}; // @[Switch.scala 43:31:@9175.4]
  assign _T_19414 = {output_30_23,output_30_22,output_30_21,output_30_20,output_30_19,output_30_18,output_30_17,output_30_16}; // @[Switch.scala 43:31:@9182.4]
  assign _T_19423 = {output_30_31,output_30_30,output_30_29,output_30_28,output_30_27,output_30_26,output_30_25,output_30_24,_T_19414,_T_19407}; // @[Switch.scala 43:31:@9191.4]
  assign _T_19427 = select_0 == 5'h1f; // @[Switch.scala 41:52:@9194.4]
  assign output_31_0 = io_outValid_0 & _T_19427; // @[Switch.scala 41:38:@9195.4]
  assign _T_19430 = select_1 == 5'h1f; // @[Switch.scala 41:52:@9197.4]
  assign output_31_1 = io_outValid_1 & _T_19430; // @[Switch.scala 41:38:@9198.4]
  assign _T_19433 = select_2 == 5'h1f; // @[Switch.scala 41:52:@9200.4]
  assign output_31_2 = io_outValid_2 & _T_19433; // @[Switch.scala 41:38:@9201.4]
  assign _T_19436 = select_3 == 5'h1f; // @[Switch.scala 41:52:@9203.4]
  assign output_31_3 = io_outValid_3 & _T_19436; // @[Switch.scala 41:38:@9204.4]
  assign _T_19439 = select_4 == 5'h1f; // @[Switch.scala 41:52:@9206.4]
  assign output_31_4 = io_outValid_4 & _T_19439; // @[Switch.scala 41:38:@9207.4]
  assign _T_19442 = select_5 == 5'h1f; // @[Switch.scala 41:52:@9209.4]
  assign output_31_5 = io_outValid_5 & _T_19442; // @[Switch.scala 41:38:@9210.4]
  assign _T_19445 = select_6 == 5'h1f; // @[Switch.scala 41:52:@9212.4]
  assign output_31_6 = io_outValid_6 & _T_19445; // @[Switch.scala 41:38:@9213.4]
  assign _T_19448 = select_7 == 5'h1f; // @[Switch.scala 41:52:@9215.4]
  assign output_31_7 = io_outValid_7 & _T_19448; // @[Switch.scala 41:38:@9216.4]
  assign _T_19451 = select_8 == 5'h1f; // @[Switch.scala 41:52:@9218.4]
  assign output_31_8 = io_outValid_8 & _T_19451; // @[Switch.scala 41:38:@9219.4]
  assign _T_19454 = select_9 == 5'h1f; // @[Switch.scala 41:52:@9221.4]
  assign output_31_9 = io_outValid_9 & _T_19454; // @[Switch.scala 41:38:@9222.4]
  assign _T_19457 = select_10 == 5'h1f; // @[Switch.scala 41:52:@9224.4]
  assign output_31_10 = io_outValid_10 & _T_19457; // @[Switch.scala 41:38:@9225.4]
  assign _T_19460 = select_11 == 5'h1f; // @[Switch.scala 41:52:@9227.4]
  assign output_31_11 = io_outValid_11 & _T_19460; // @[Switch.scala 41:38:@9228.4]
  assign _T_19463 = select_12 == 5'h1f; // @[Switch.scala 41:52:@9230.4]
  assign output_31_12 = io_outValid_12 & _T_19463; // @[Switch.scala 41:38:@9231.4]
  assign _T_19466 = select_13 == 5'h1f; // @[Switch.scala 41:52:@9233.4]
  assign output_31_13 = io_outValid_13 & _T_19466; // @[Switch.scala 41:38:@9234.4]
  assign _T_19469 = select_14 == 5'h1f; // @[Switch.scala 41:52:@9236.4]
  assign output_31_14 = io_outValid_14 & _T_19469; // @[Switch.scala 41:38:@9237.4]
  assign _T_19472 = select_15 == 5'h1f; // @[Switch.scala 41:52:@9239.4]
  assign output_31_15 = io_outValid_15 & _T_19472; // @[Switch.scala 41:38:@9240.4]
  assign _T_19475 = select_16 == 5'h1f; // @[Switch.scala 41:52:@9242.4]
  assign output_31_16 = io_outValid_16 & _T_19475; // @[Switch.scala 41:38:@9243.4]
  assign _T_19478 = select_17 == 5'h1f; // @[Switch.scala 41:52:@9245.4]
  assign output_31_17 = io_outValid_17 & _T_19478; // @[Switch.scala 41:38:@9246.4]
  assign _T_19481 = select_18 == 5'h1f; // @[Switch.scala 41:52:@9248.4]
  assign output_31_18 = io_outValid_18 & _T_19481; // @[Switch.scala 41:38:@9249.4]
  assign _T_19484 = select_19 == 5'h1f; // @[Switch.scala 41:52:@9251.4]
  assign output_31_19 = io_outValid_19 & _T_19484; // @[Switch.scala 41:38:@9252.4]
  assign _T_19487 = select_20 == 5'h1f; // @[Switch.scala 41:52:@9254.4]
  assign output_31_20 = io_outValid_20 & _T_19487; // @[Switch.scala 41:38:@9255.4]
  assign _T_19490 = select_21 == 5'h1f; // @[Switch.scala 41:52:@9257.4]
  assign output_31_21 = io_outValid_21 & _T_19490; // @[Switch.scala 41:38:@9258.4]
  assign _T_19493 = select_22 == 5'h1f; // @[Switch.scala 41:52:@9260.4]
  assign output_31_22 = io_outValid_22 & _T_19493; // @[Switch.scala 41:38:@9261.4]
  assign _T_19496 = select_23 == 5'h1f; // @[Switch.scala 41:52:@9263.4]
  assign output_31_23 = io_outValid_23 & _T_19496; // @[Switch.scala 41:38:@9264.4]
  assign _T_19499 = select_24 == 5'h1f; // @[Switch.scala 41:52:@9266.4]
  assign output_31_24 = io_outValid_24 & _T_19499; // @[Switch.scala 41:38:@9267.4]
  assign _T_19502 = select_25 == 5'h1f; // @[Switch.scala 41:52:@9269.4]
  assign output_31_25 = io_outValid_25 & _T_19502; // @[Switch.scala 41:38:@9270.4]
  assign _T_19505 = select_26 == 5'h1f; // @[Switch.scala 41:52:@9272.4]
  assign output_31_26 = io_outValid_26 & _T_19505; // @[Switch.scala 41:38:@9273.4]
  assign _T_19508 = select_27 == 5'h1f; // @[Switch.scala 41:52:@9275.4]
  assign output_31_27 = io_outValid_27 & _T_19508; // @[Switch.scala 41:38:@9276.4]
  assign _T_19511 = select_28 == 5'h1f; // @[Switch.scala 41:52:@9278.4]
  assign output_31_28 = io_outValid_28 & _T_19511; // @[Switch.scala 41:38:@9279.4]
  assign _T_19514 = select_29 == 5'h1f; // @[Switch.scala 41:52:@9281.4]
  assign output_31_29 = io_outValid_29 & _T_19514; // @[Switch.scala 41:38:@9282.4]
  assign _T_19517 = select_30 == 5'h1f; // @[Switch.scala 41:52:@9284.4]
  assign output_31_30 = io_outValid_30 & _T_19517; // @[Switch.scala 41:38:@9285.4]
  assign _T_19520 = select_31 == 5'h1f; // @[Switch.scala 41:52:@9287.4]
  assign output_31_31 = io_outValid_31 & _T_19520; // @[Switch.scala 41:38:@9288.4]
  assign _T_19528 = {output_31_7,output_31_6,output_31_5,output_31_4,output_31_3,output_31_2,output_31_1,output_31_0}; // @[Switch.scala 43:31:@9296.4]
  assign _T_19536 = {output_31_15,output_31_14,output_31_13,output_31_12,output_31_11,output_31_10,output_31_9,output_31_8,_T_19528}; // @[Switch.scala 43:31:@9304.4]
  assign _T_19543 = {output_31_23,output_31_22,output_31_21,output_31_20,output_31_19,output_31_18,output_31_17,output_31_16}; // @[Switch.scala 43:31:@9311.4]
  assign _T_19552 = {output_31_31,output_31_30,output_31_29,output_31_28,output_31_27,output_31_26,output_31_25,output_31_24,_T_19543,_T_19536}; // @[Switch.scala 43:31:@9320.4]
  assign io_outAck_0 = _T_15553 != 32'h0; // @[Switch.scala 43:18:@5323.4]
  assign io_outAck_1 = _T_15682 != 32'h0; // @[Switch.scala 43:18:@5452.4]
  assign io_outAck_2 = _T_15811 != 32'h0; // @[Switch.scala 43:18:@5581.4]
  assign io_outAck_3 = _T_15940 != 32'h0; // @[Switch.scala 43:18:@5710.4]
  assign io_outAck_4 = _T_16069 != 32'h0; // @[Switch.scala 43:18:@5839.4]
  assign io_outAck_5 = _T_16198 != 32'h0; // @[Switch.scala 43:18:@5968.4]
  assign io_outAck_6 = _T_16327 != 32'h0; // @[Switch.scala 43:18:@6097.4]
  assign io_outAck_7 = _T_16456 != 32'h0; // @[Switch.scala 43:18:@6226.4]
  assign io_outAck_8 = _T_16585 != 32'h0; // @[Switch.scala 43:18:@6355.4]
  assign io_outAck_9 = _T_16714 != 32'h0; // @[Switch.scala 43:18:@6484.4]
  assign io_outAck_10 = _T_16843 != 32'h0; // @[Switch.scala 43:18:@6613.4]
  assign io_outAck_11 = _T_16972 != 32'h0; // @[Switch.scala 43:18:@6742.4]
  assign io_outAck_12 = _T_17101 != 32'h0; // @[Switch.scala 43:18:@6871.4]
  assign io_outAck_13 = _T_17230 != 32'h0; // @[Switch.scala 43:18:@7000.4]
  assign io_outAck_14 = _T_17359 != 32'h0; // @[Switch.scala 43:18:@7129.4]
  assign io_outAck_15 = _T_17488 != 32'h0; // @[Switch.scala 43:18:@7258.4]
  assign io_outAck_16 = _T_17617 != 32'h0; // @[Switch.scala 43:18:@7387.4]
  assign io_outAck_17 = _T_17746 != 32'h0; // @[Switch.scala 43:18:@7516.4]
  assign io_outAck_18 = _T_17875 != 32'h0; // @[Switch.scala 43:18:@7645.4]
  assign io_outAck_19 = _T_18004 != 32'h0; // @[Switch.scala 43:18:@7774.4]
  assign io_outAck_20 = _T_18133 != 32'h0; // @[Switch.scala 43:18:@7903.4]
  assign io_outAck_21 = _T_18262 != 32'h0; // @[Switch.scala 43:18:@8032.4]
  assign io_outAck_22 = _T_18391 != 32'h0; // @[Switch.scala 43:18:@8161.4]
  assign io_outAck_23 = _T_18520 != 32'h0; // @[Switch.scala 43:18:@8290.4]
  assign io_outAck_24 = _T_18649 != 32'h0; // @[Switch.scala 43:18:@8419.4]
  assign io_outAck_25 = _T_18778 != 32'h0; // @[Switch.scala 43:18:@8548.4]
  assign io_outAck_26 = _T_18907 != 32'h0; // @[Switch.scala 43:18:@8677.4]
  assign io_outAck_27 = _T_19036 != 32'h0; // @[Switch.scala 43:18:@8806.4]
  assign io_outAck_28 = _T_19165 != 32'h0; // @[Switch.scala 43:18:@8935.4]
  assign io_outAck_29 = _T_19294 != 32'h0; // @[Switch.scala 43:18:@9064.4]
  assign io_outAck_30 = _T_19423 != 32'h0; // @[Switch.scala 43:18:@9193.4]
  assign io_outAck_31 = _T_19552 != 32'h0; // @[Switch.scala 43:18:@9322.4]
  assign io_outData_0 = 5'h1f == select_0 ? io_inData_31 : _GEN_30; // @[Switch.scala 33:19:@138.4]
  assign io_outData_1 = 5'h1f == select_1 ? io_inData_31 : _GEN_62; // @[Switch.scala 33:19:@300.4]
  assign io_outData_2 = 5'h1f == select_2 ? io_inData_31 : _GEN_94; // @[Switch.scala 33:19:@462.4]
  assign io_outData_3 = 5'h1f == select_3 ? io_inData_31 : _GEN_126; // @[Switch.scala 33:19:@624.4]
  assign io_outData_4 = 5'h1f == select_4 ? io_inData_31 : _GEN_158; // @[Switch.scala 33:19:@786.4]
  assign io_outData_5 = 5'h1f == select_5 ? io_inData_31 : _GEN_190; // @[Switch.scala 33:19:@948.4]
  assign io_outData_6 = 5'h1f == select_6 ? io_inData_31 : _GEN_222; // @[Switch.scala 33:19:@1110.4]
  assign io_outData_7 = 5'h1f == select_7 ? io_inData_31 : _GEN_254; // @[Switch.scala 33:19:@1272.4]
  assign io_outData_8 = 5'h1f == select_8 ? io_inData_31 : _GEN_286; // @[Switch.scala 33:19:@1434.4]
  assign io_outData_9 = 5'h1f == select_9 ? io_inData_31 : _GEN_318; // @[Switch.scala 33:19:@1596.4]
  assign io_outData_10 = 5'h1f == select_10 ? io_inData_31 : _GEN_350; // @[Switch.scala 33:19:@1758.4]
  assign io_outData_11 = 5'h1f == select_11 ? io_inData_31 : _GEN_382; // @[Switch.scala 33:19:@1920.4]
  assign io_outData_12 = 5'h1f == select_12 ? io_inData_31 : _GEN_414; // @[Switch.scala 33:19:@2082.4]
  assign io_outData_13 = 5'h1f == select_13 ? io_inData_31 : _GEN_446; // @[Switch.scala 33:19:@2244.4]
  assign io_outData_14 = 5'h1f == select_14 ? io_inData_31 : _GEN_478; // @[Switch.scala 33:19:@2406.4]
  assign io_outData_15 = 5'h1f == select_15 ? io_inData_31 : _GEN_510; // @[Switch.scala 33:19:@2568.4]
  assign io_outData_16 = 5'h1f == select_16 ? io_inData_31 : _GEN_542; // @[Switch.scala 33:19:@2730.4]
  assign io_outData_17 = 5'h1f == select_17 ? io_inData_31 : _GEN_574; // @[Switch.scala 33:19:@2892.4]
  assign io_outData_18 = 5'h1f == select_18 ? io_inData_31 : _GEN_606; // @[Switch.scala 33:19:@3054.4]
  assign io_outData_19 = 5'h1f == select_19 ? io_inData_31 : _GEN_638; // @[Switch.scala 33:19:@3216.4]
  assign io_outData_20 = 5'h1f == select_20 ? io_inData_31 : _GEN_670; // @[Switch.scala 33:19:@3378.4]
  assign io_outData_21 = 5'h1f == select_21 ? io_inData_31 : _GEN_702; // @[Switch.scala 33:19:@3540.4]
  assign io_outData_22 = 5'h1f == select_22 ? io_inData_31 : _GEN_734; // @[Switch.scala 33:19:@3702.4]
  assign io_outData_23 = 5'h1f == select_23 ? io_inData_31 : _GEN_766; // @[Switch.scala 33:19:@3864.4]
  assign io_outData_24 = 5'h1f == select_24 ? io_inData_31 : _GEN_798; // @[Switch.scala 33:19:@4026.4]
  assign io_outData_25 = 5'h1f == select_25 ? io_inData_31 : _GEN_830; // @[Switch.scala 33:19:@4188.4]
  assign io_outData_26 = 5'h1f == select_26 ? io_inData_31 : _GEN_862; // @[Switch.scala 33:19:@4350.4]
  assign io_outData_27 = 5'h1f == select_27 ? io_inData_31 : _GEN_894; // @[Switch.scala 33:19:@4512.4]
  assign io_outData_28 = 5'h1f == select_28 ? io_inData_31 : _GEN_926; // @[Switch.scala 33:19:@4674.4]
  assign io_outData_29 = 5'h1f == select_29 ? io_inData_31 : _GEN_958; // @[Switch.scala 33:19:@4836.4]
  assign io_outData_30 = 5'h1f == select_30 ? io_inData_31 : _GEN_990; // @[Switch.scala 33:19:@4998.4]
  assign io_outData_31 = 5'h1f == select_31 ? io_inData_31 : _GEN_1022; // @[Switch.scala 33:19:@5160.4]
  assign io_outValid_0 = _T_4947 != 32'h0; // @[Switch.scala 34:20:@171.4]
  assign io_outValid_1 = _T_5140 != 32'h0; // @[Switch.scala 34:20:@333.4]
  assign io_outValid_2 = _T_5333 != 32'h0; // @[Switch.scala 34:20:@495.4]
  assign io_outValid_3 = _T_5526 != 32'h0; // @[Switch.scala 34:20:@657.4]
  assign io_outValid_4 = _T_5719 != 32'h0; // @[Switch.scala 34:20:@819.4]
  assign io_outValid_5 = _T_5912 != 32'h0; // @[Switch.scala 34:20:@981.4]
  assign io_outValid_6 = _T_6105 != 32'h0; // @[Switch.scala 34:20:@1143.4]
  assign io_outValid_7 = _T_6298 != 32'h0; // @[Switch.scala 34:20:@1305.4]
  assign io_outValid_8 = _T_6491 != 32'h0; // @[Switch.scala 34:20:@1467.4]
  assign io_outValid_9 = _T_6684 != 32'h0; // @[Switch.scala 34:20:@1629.4]
  assign io_outValid_10 = _T_6877 != 32'h0; // @[Switch.scala 34:20:@1791.4]
  assign io_outValid_11 = _T_7070 != 32'h0; // @[Switch.scala 34:20:@1953.4]
  assign io_outValid_12 = _T_7263 != 32'h0; // @[Switch.scala 34:20:@2115.4]
  assign io_outValid_13 = _T_7456 != 32'h0; // @[Switch.scala 34:20:@2277.4]
  assign io_outValid_14 = _T_7649 != 32'h0; // @[Switch.scala 34:20:@2439.4]
  assign io_outValid_15 = _T_7842 != 32'h0; // @[Switch.scala 34:20:@2601.4]
  assign io_outValid_16 = _T_8035 != 32'h0; // @[Switch.scala 34:20:@2763.4]
  assign io_outValid_17 = _T_8228 != 32'h0; // @[Switch.scala 34:20:@2925.4]
  assign io_outValid_18 = _T_8421 != 32'h0; // @[Switch.scala 34:20:@3087.4]
  assign io_outValid_19 = _T_8614 != 32'h0; // @[Switch.scala 34:20:@3249.4]
  assign io_outValid_20 = _T_8807 != 32'h0; // @[Switch.scala 34:20:@3411.4]
  assign io_outValid_21 = _T_9000 != 32'h0; // @[Switch.scala 34:20:@3573.4]
  assign io_outValid_22 = _T_9193 != 32'h0; // @[Switch.scala 34:20:@3735.4]
  assign io_outValid_23 = _T_9386 != 32'h0; // @[Switch.scala 34:20:@3897.4]
  assign io_outValid_24 = _T_9579 != 32'h0; // @[Switch.scala 34:20:@4059.4]
  assign io_outValid_25 = _T_9772 != 32'h0; // @[Switch.scala 34:20:@4221.4]
  assign io_outValid_26 = _T_9965 != 32'h0; // @[Switch.scala 34:20:@4383.4]
  assign io_outValid_27 = _T_10158 != 32'h0; // @[Switch.scala 34:20:@4545.4]
  assign io_outValid_28 = _T_10351 != 32'h0; // @[Switch.scala 34:20:@4707.4]
  assign io_outValid_29 = _T_10544 != 32'h0; // @[Switch.scala 34:20:@4869.4]
  assign io_outValid_30 = _T_10737 != 32'h0; // @[Switch.scala 34:20:@5031.4]
  assign io_outValid_31 = _T_10930 != 32'h0; // @[Switch.scala 34:20:@5193.4]
endmodule
module SwitchWrapper( // @[:@9324.2]
  input         clock, // @[:@9325.4]
  input         reset, // @[:@9326.4]
  input  [4:0]  io_inAddr_0, // @[:@9327.4]
  input  [4:0]  io_inAddr_1, // @[:@9327.4]
  input  [4:0]  io_inAddr_2, // @[:@9327.4]
  input  [4:0]  io_inAddr_3, // @[:@9327.4]
  input  [4:0]  io_inAddr_4, // @[:@9327.4]
  input  [4:0]  io_inAddr_5, // @[:@9327.4]
  input  [4:0]  io_inAddr_6, // @[:@9327.4]
  input  [4:0]  io_inAddr_7, // @[:@9327.4]
  input  [4:0]  io_inAddr_8, // @[:@9327.4]
  input  [4:0]  io_inAddr_9, // @[:@9327.4]
  input  [4:0]  io_inAddr_10, // @[:@9327.4]
  input  [4:0]  io_inAddr_11, // @[:@9327.4]
  input  [4:0]  io_inAddr_12, // @[:@9327.4]
  input  [4:0]  io_inAddr_13, // @[:@9327.4]
  input  [4:0]  io_inAddr_14, // @[:@9327.4]
  input  [4:0]  io_inAddr_15, // @[:@9327.4]
  input  [4:0]  io_inAddr_16, // @[:@9327.4]
  input  [4:0]  io_inAddr_17, // @[:@9327.4]
  input  [4:0]  io_inAddr_18, // @[:@9327.4]
  input  [4:0]  io_inAddr_19, // @[:@9327.4]
  input  [4:0]  io_inAddr_20, // @[:@9327.4]
  input  [4:0]  io_inAddr_21, // @[:@9327.4]
  input  [4:0]  io_inAddr_22, // @[:@9327.4]
  input  [4:0]  io_inAddr_23, // @[:@9327.4]
  input  [4:0]  io_inAddr_24, // @[:@9327.4]
  input  [4:0]  io_inAddr_25, // @[:@9327.4]
  input  [4:0]  io_inAddr_26, // @[:@9327.4]
  input  [4:0]  io_inAddr_27, // @[:@9327.4]
  input  [4:0]  io_inAddr_28, // @[:@9327.4]
  input  [4:0]  io_inAddr_29, // @[:@9327.4]
  input  [4:0]  io_inAddr_30, // @[:@9327.4]
  input  [4:0]  io_inAddr_31, // @[:@9327.4]
  input  [47:0] io_inData_0, // @[:@9327.4]
  input  [47:0] io_inData_1, // @[:@9327.4]
  input  [47:0] io_inData_2, // @[:@9327.4]
  input  [47:0] io_inData_3, // @[:@9327.4]
  input  [47:0] io_inData_4, // @[:@9327.4]
  input  [47:0] io_inData_5, // @[:@9327.4]
  input  [47:0] io_inData_6, // @[:@9327.4]
  input  [47:0] io_inData_7, // @[:@9327.4]
  input  [47:0] io_inData_8, // @[:@9327.4]
  input  [47:0] io_inData_9, // @[:@9327.4]
  input  [47:0] io_inData_10, // @[:@9327.4]
  input  [47:0] io_inData_11, // @[:@9327.4]
  input  [47:0] io_inData_12, // @[:@9327.4]
  input  [47:0] io_inData_13, // @[:@9327.4]
  input  [47:0] io_inData_14, // @[:@9327.4]
  input  [47:0] io_inData_15, // @[:@9327.4]
  input  [47:0] io_inData_16, // @[:@9327.4]
  input  [47:0] io_inData_17, // @[:@9327.4]
  input  [47:0] io_inData_18, // @[:@9327.4]
  input  [47:0] io_inData_19, // @[:@9327.4]
  input  [47:0] io_inData_20, // @[:@9327.4]
  input  [47:0] io_inData_21, // @[:@9327.4]
  input  [47:0] io_inData_22, // @[:@9327.4]
  input  [47:0] io_inData_23, // @[:@9327.4]
  input  [47:0] io_inData_24, // @[:@9327.4]
  input  [47:0] io_inData_25, // @[:@9327.4]
  input  [47:0] io_inData_26, // @[:@9327.4]
  input  [47:0] io_inData_27, // @[:@9327.4]
  input  [47:0] io_inData_28, // @[:@9327.4]
  input  [47:0] io_inData_29, // @[:@9327.4]
  input  [47:0] io_inData_30, // @[:@9327.4]
  input  [47:0] io_inData_31, // @[:@9327.4]
  input         io_inValid_0, // @[:@9327.4]
  input         io_inValid_1, // @[:@9327.4]
  input         io_inValid_2, // @[:@9327.4]
  input         io_inValid_3, // @[:@9327.4]
  input         io_inValid_4, // @[:@9327.4]
  input         io_inValid_5, // @[:@9327.4]
  input         io_inValid_6, // @[:@9327.4]
  input         io_inValid_7, // @[:@9327.4]
  input         io_inValid_8, // @[:@9327.4]
  input         io_inValid_9, // @[:@9327.4]
  input         io_inValid_10, // @[:@9327.4]
  input         io_inValid_11, // @[:@9327.4]
  input         io_inValid_12, // @[:@9327.4]
  input         io_inValid_13, // @[:@9327.4]
  input         io_inValid_14, // @[:@9327.4]
  input         io_inValid_15, // @[:@9327.4]
  input         io_inValid_16, // @[:@9327.4]
  input         io_inValid_17, // @[:@9327.4]
  input         io_inValid_18, // @[:@9327.4]
  input         io_inValid_19, // @[:@9327.4]
  input         io_inValid_20, // @[:@9327.4]
  input         io_inValid_21, // @[:@9327.4]
  input         io_inValid_22, // @[:@9327.4]
  input         io_inValid_23, // @[:@9327.4]
  input         io_inValid_24, // @[:@9327.4]
  input         io_inValid_25, // @[:@9327.4]
  input         io_inValid_26, // @[:@9327.4]
  input         io_inValid_27, // @[:@9327.4]
  input         io_inValid_28, // @[:@9327.4]
  input         io_inValid_29, // @[:@9327.4]
  input         io_inValid_30, // @[:@9327.4]
  input         io_inValid_31, // @[:@9327.4]
  output        io_outAck_0, // @[:@9327.4]
  output        io_outAck_1, // @[:@9327.4]
  output        io_outAck_2, // @[:@9327.4]
  output        io_outAck_3, // @[:@9327.4]
  output        io_outAck_4, // @[:@9327.4]
  output        io_outAck_5, // @[:@9327.4]
  output        io_outAck_6, // @[:@9327.4]
  output        io_outAck_7, // @[:@9327.4]
  output        io_outAck_8, // @[:@9327.4]
  output        io_outAck_9, // @[:@9327.4]
  output        io_outAck_10, // @[:@9327.4]
  output        io_outAck_11, // @[:@9327.4]
  output        io_outAck_12, // @[:@9327.4]
  output        io_outAck_13, // @[:@9327.4]
  output        io_outAck_14, // @[:@9327.4]
  output        io_outAck_15, // @[:@9327.4]
  output        io_outAck_16, // @[:@9327.4]
  output        io_outAck_17, // @[:@9327.4]
  output        io_outAck_18, // @[:@9327.4]
  output        io_outAck_19, // @[:@9327.4]
  output        io_outAck_20, // @[:@9327.4]
  output        io_outAck_21, // @[:@9327.4]
  output        io_outAck_22, // @[:@9327.4]
  output        io_outAck_23, // @[:@9327.4]
  output        io_outAck_24, // @[:@9327.4]
  output        io_outAck_25, // @[:@9327.4]
  output        io_outAck_26, // @[:@9327.4]
  output        io_outAck_27, // @[:@9327.4]
  output        io_outAck_28, // @[:@9327.4]
  output        io_outAck_29, // @[:@9327.4]
  output        io_outAck_30, // @[:@9327.4]
  output        io_outAck_31, // @[:@9327.4]
  output [47:0] io_outData_0, // @[:@9327.4]
  output [47:0] io_outData_1, // @[:@9327.4]
  output [47:0] io_outData_2, // @[:@9327.4]
  output [47:0] io_outData_3, // @[:@9327.4]
  output [47:0] io_outData_4, // @[:@9327.4]
  output [47:0] io_outData_5, // @[:@9327.4]
  output [47:0] io_outData_6, // @[:@9327.4]
  output [47:0] io_outData_7, // @[:@9327.4]
  output [47:0] io_outData_8, // @[:@9327.4]
  output [47:0] io_outData_9, // @[:@9327.4]
  output [47:0] io_outData_10, // @[:@9327.4]
  output [47:0] io_outData_11, // @[:@9327.4]
  output [47:0] io_outData_12, // @[:@9327.4]
  output [47:0] io_outData_13, // @[:@9327.4]
  output [47:0] io_outData_14, // @[:@9327.4]
  output [47:0] io_outData_15, // @[:@9327.4]
  output [47:0] io_outData_16, // @[:@9327.4]
  output [47:0] io_outData_17, // @[:@9327.4]
  output [47:0] io_outData_18, // @[:@9327.4]
  output [47:0] io_outData_19, // @[:@9327.4]
  output [47:0] io_outData_20, // @[:@9327.4]
  output [47:0] io_outData_21, // @[:@9327.4]
  output [47:0] io_outData_22, // @[:@9327.4]
  output [47:0] io_outData_23, // @[:@9327.4]
  output [47:0] io_outData_24, // @[:@9327.4]
  output [47:0] io_outData_25, // @[:@9327.4]
  output [47:0] io_outData_26, // @[:@9327.4]
  output [47:0] io_outData_27, // @[:@9327.4]
  output [47:0] io_outData_28, // @[:@9327.4]
  output [47:0] io_outData_29, // @[:@9327.4]
  output [47:0] io_outData_30, // @[:@9327.4]
  output [47:0] io_outData_31, // @[:@9327.4]
  output        io_outValid_0, // @[:@9327.4]
  output        io_outValid_1, // @[:@9327.4]
  output        io_outValid_2, // @[:@9327.4]
  output        io_outValid_3, // @[:@9327.4]
  output        io_outValid_4, // @[:@9327.4]
  output        io_outValid_5, // @[:@9327.4]
  output        io_outValid_6, // @[:@9327.4]
  output        io_outValid_7, // @[:@9327.4]
  output        io_outValid_8, // @[:@9327.4]
  output        io_outValid_9, // @[:@9327.4]
  output        io_outValid_10, // @[:@9327.4]
  output        io_outValid_11, // @[:@9327.4]
  output        io_outValid_12, // @[:@9327.4]
  output        io_outValid_13, // @[:@9327.4]
  output        io_outValid_14, // @[:@9327.4]
  output        io_outValid_15, // @[:@9327.4]
  output        io_outValid_16, // @[:@9327.4]
  output        io_outValid_17, // @[:@9327.4]
  output        io_outValid_18, // @[:@9327.4]
  output        io_outValid_19, // @[:@9327.4]
  output        io_outValid_20, // @[:@9327.4]
  output        io_outValid_21, // @[:@9327.4]
  output        io_outValid_22, // @[:@9327.4]
  output        io_outValid_23, // @[:@9327.4]
  output        io_outValid_24, // @[:@9327.4]
  output        io_outValid_25, // @[:@9327.4]
  output        io_outValid_26, // @[:@9327.4]
  output        io_outValid_27, // @[:@9327.4]
  output        io_outValid_28, // @[:@9327.4]
  output        io_outValid_29, // @[:@9327.4]
  output        io_outValid_30, // @[:@9327.4]
  output        io_outValid_31 // @[:@9327.4]
);
  wire [4:0] switch_io_inAddr_0; // @[Switch.scala 50:22:@9329.4]
  wire [4:0] switch_io_inAddr_1; // @[Switch.scala 50:22:@9329.4]
  wire [4:0] switch_io_inAddr_2; // @[Switch.scala 50:22:@9329.4]
  wire [4:0] switch_io_inAddr_3; // @[Switch.scala 50:22:@9329.4]
  wire [4:0] switch_io_inAddr_4; // @[Switch.scala 50:22:@9329.4]
  wire [4:0] switch_io_inAddr_5; // @[Switch.scala 50:22:@9329.4]
  wire [4:0] switch_io_inAddr_6; // @[Switch.scala 50:22:@9329.4]
  wire [4:0] switch_io_inAddr_7; // @[Switch.scala 50:22:@9329.4]
  wire [4:0] switch_io_inAddr_8; // @[Switch.scala 50:22:@9329.4]
  wire [4:0] switch_io_inAddr_9; // @[Switch.scala 50:22:@9329.4]
  wire [4:0] switch_io_inAddr_10; // @[Switch.scala 50:22:@9329.4]
  wire [4:0] switch_io_inAddr_11; // @[Switch.scala 50:22:@9329.4]
  wire [4:0] switch_io_inAddr_12; // @[Switch.scala 50:22:@9329.4]
  wire [4:0] switch_io_inAddr_13; // @[Switch.scala 50:22:@9329.4]
  wire [4:0] switch_io_inAddr_14; // @[Switch.scala 50:22:@9329.4]
  wire [4:0] switch_io_inAddr_15; // @[Switch.scala 50:22:@9329.4]
  wire [4:0] switch_io_inAddr_16; // @[Switch.scala 50:22:@9329.4]
  wire [4:0] switch_io_inAddr_17; // @[Switch.scala 50:22:@9329.4]
  wire [4:0] switch_io_inAddr_18; // @[Switch.scala 50:22:@9329.4]
  wire [4:0] switch_io_inAddr_19; // @[Switch.scala 50:22:@9329.4]
  wire [4:0] switch_io_inAddr_20; // @[Switch.scala 50:22:@9329.4]
  wire [4:0] switch_io_inAddr_21; // @[Switch.scala 50:22:@9329.4]
  wire [4:0] switch_io_inAddr_22; // @[Switch.scala 50:22:@9329.4]
  wire [4:0] switch_io_inAddr_23; // @[Switch.scala 50:22:@9329.4]
  wire [4:0] switch_io_inAddr_24; // @[Switch.scala 50:22:@9329.4]
  wire [4:0] switch_io_inAddr_25; // @[Switch.scala 50:22:@9329.4]
  wire [4:0] switch_io_inAddr_26; // @[Switch.scala 50:22:@9329.4]
  wire [4:0] switch_io_inAddr_27; // @[Switch.scala 50:22:@9329.4]
  wire [4:0] switch_io_inAddr_28; // @[Switch.scala 50:22:@9329.4]
  wire [4:0] switch_io_inAddr_29; // @[Switch.scala 50:22:@9329.4]
  wire [4:0] switch_io_inAddr_30; // @[Switch.scala 50:22:@9329.4]
  wire [4:0] switch_io_inAddr_31; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_inData_0; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_inData_1; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_inData_2; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_inData_3; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_inData_4; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_inData_5; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_inData_6; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_inData_7; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_inData_8; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_inData_9; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_inData_10; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_inData_11; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_inData_12; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_inData_13; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_inData_14; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_inData_15; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_inData_16; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_inData_17; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_inData_18; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_inData_19; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_inData_20; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_inData_21; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_inData_22; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_inData_23; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_inData_24; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_inData_25; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_inData_26; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_inData_27; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_inData_28; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_inData_29; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_inData_30; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_inData_31; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_inValid_0; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_inValid_1; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_inValid_2; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_inValid_3; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_inValid_4; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_inValid_5; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_inValid_6; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_inValid_7; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_inValid_8; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_inValid_9; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_inValid_10; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_inValid_11; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_inValid_12; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_inValid_13; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_inValid_14; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_inValid_15; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_inValid_16; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_inValid_17; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_inValid_18; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_inValid_19; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_inValid_20; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_inValid_21; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_inValid_22; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_inValid_23; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_inValid_24; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_inValid_25; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_inValid_26; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_inValid_27; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_inValid_28; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_inValid_29; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_inValid_30; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_inValid_31; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outAck_0; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outAck_1; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outAck_2; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outAck_3; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outAck_4; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outAck_5; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outAck_6; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outAck_7; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outAck_8; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outAck_9; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outAck_10; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outAck_11; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outAck_12; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outAck_13; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outAck_14; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outAck_15; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outAck_16; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outAck_17; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outAck_18; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outAck_19; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outAck_20; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outAck_21; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outAck_22; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outAck_23; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outAck_24; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outAck_25; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outAck_26; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outAck_27; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outAck_28; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outAck_29; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outAck_30; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outAck_31; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_outData_0; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_outData_1; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_outData_2; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_outData_3; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_outData_4; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_outData_5; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_outData_6; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_outData_7; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_outData_8; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_outData_9; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_outData_10; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_outData_11; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_outData_12; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_outData_13; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_outData_14; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_outData_15; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_outData_16; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_outData_17; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_outData_18; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_outData_19; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_outData_20; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_outData_21; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_outData_22; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_outData_23; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_outData_24; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_outData_25; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_outData_26; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_outData_27; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_outData_28; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_outData_29; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_outData_30; // @[Switch.scala 50:22:@9329.4]
  wire [47:0] switch_io_outData_31; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outValid_0; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outValid_1; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outValid_2; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outValid_3; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outValid_4; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outValid_5; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outValid_6; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outValid_7; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outValid_8; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outValid_9; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outValid_10; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outValid_11; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outValid_12; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outValid_13; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outValid_14; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outValid_15; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outValid_16; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outValid_17; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outValid_18; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outValid_19; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outValid_20; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outValid_21; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outValid_22; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outValid_23; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outValid_24; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outValid_25; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outValid_26; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outValid_27; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outValid_28; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outValid_29; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outValid_30; // @[Switch.scala 50:22:@9329.4]
  wire  switch_io_outValid_31; // @[Switch.scala 50:22:@9329.4]
  reg [4:0] _T_294_0; // @[Switch.scala 51:30:@9332.4]
  reg [31:0] _RAND_0;
  reg [4:0] _T_294_1; // @[Switch.scala 51:30:@9332.4]
  reg [31:0] _RAND_1;
  reg [4:0] _T_294_2; // @[Switch.scala 51:30:@9332.4]
  reg [31:0] _RAND_2;
  reg [4:0] _T_294_3; // @[Switch.scala 51:30:@9332.4]
  reg [31:0] _RAND_3;
  reg [4:0] _T_294_4; // @[Switch.scala 51:30:@9332.4]
  reg [31:0] _RAND_4;
  reg [4:0] _T_294_5; // @[Switch.scala 51:30:@9332.4]
  reg [31:0] _RAND_5;
  reg [4:0] _T_294_6; // @[Switch.scala 51:30:@9332.4]
  reg [31:0] _RAND_6;
  reg [4:0] _T_294_7; // @[Switch.scala 51:30:@9332.4]
  reg [31:0] _RAND_7;
  reg [4:0] _T_294_8; // @[Switch.scala 51:30:@9332.4]
  reg [31:0] _RAND_8;
  reg [4:0] _T_294_9; // @[Switch.scala 51:30:@9332.4]
  reg [31:0] _RAND_9;
  reg [4:0] _T_294_10; // @[Switch.scala 51:30:@9332.4]
  reg [31:0] _RAND_10;
  reg [4:0] _T_294_11; // @[Switch.scala 51:30:@9332.4]
  reg [31:0] _RAND_11;
  reg [4:0] _T_294_12; // @[Switch.scala 51:30:@9332.4]
  reg [31:0] _RAND_12;
  reg [4:0] _T_294_13; // @[Switch.scala 51:30:@9332.4]
  reg [31:0] _RAND_13;
  reg [4:0] _T_294_14; // @[Switch.scala 51:30:@9332.4]
  reg [31:0] _RAND_14;
  reg [4:0] _T_294_15; // @[Switch.scala 51:30:@9332.4]
  reg [31:0] _RAND_15;
  reg [4:0] _T_294_16; // @[Switch.scala 51:30:@9332.4]
  reg [31:0] _RAND_16;
  reg [4:0] _T_294_17; // @[Switch.scala 51:30:@9332.4]
  reg [31:0] _RAND_17;
  reg [4:0] _T_294_18; // @[Switch.scala 51:30:@9332.4]
  reg [31:0] _RAND_18;
  reg [4:0] _T_294_19; // @[Switch.scala 51:30:@9332.4]
  reg [31:0] _RAND_19;
  reg [4:0] _T_294_20; // @[Switch.scala 51:30:@9332.4]
  reg [31:0] _RAND_20;
  reg [4:0] _T_294_21; // @[Switch.scala 51:30:@9332.4]
  reg [31:0] _RAND_21;
  reg [4:0] _T_294_22; // @[Switch.scala 51:30:@9332.4]
  reg [31:0] _RAND_22;
  reg [4:0] _T_294_23; // @[Switch.scala 51:30:@9332.4]
  reg [31:0] _RAND_23;
  reg [4:0] _T_294_24; // @[Switch.scala 51:30:@9332.4]
  reg [31:0] _RAND_24;
  reg [4:0] _T_294_25; // @[Switch.scala 51:30:@9332.4]
  reg [31:0] _RAND_25;
  reg [4:0] _T_294_26; // @[Switch.scala 51:30:@9332.4]
  reg [31:0] _RAND_26;
  reg [4:0] _T_294_27; // @[Switch.scala 51:30:@9332.4]
  reg [31:0] _RAND_27;
  reg [4:0] _T_294_28; // @[Switch.scala 51:30:@9332.4]
  reg [31:0] _RAND_28;
  reg [4:0] _T_294_29; // @[Switch.scala 51:30:@9332.4]
  reg [31:0] _RAND_29;
  reg [4:0] _T_294_30; // @[Switch.scala 51:30:@9332.4]
  reg [31:0] _RAND_30;
  reg [4:0] _T_294_31; // @[Switch.scala 51:30:@9332.4]
  reg [31:0] _RAND_31;
  reg [47:0] _T_463_0; // @[Switch.scala 52:30:@9397.4]
  reg [63:0] _RAND_32;
  reg [47:0] _T_463_1; // @[Switch.scala 52:30:@9397.4]
  reg [63:0] _RAND_33;
  reg [47:0] _T_463_2; // @[Switch.scala 52:30:@9397.4]
  reg [63:0] _RAND_34;
  reg [47:0] _T_463_3; // @[Switch.scala 52:30:@9397.4]
  reg [63:0] _RAND_35;
  reg [47:0] _T_463_4; // @[Switch.scala 52:30:@9397.4]
  reg [63:0] _RAND_36;
  reg [47:0] _T_463_5; // @[Switch.scala 52:30:@9397.4]
  reg [63:0] _RAND_37;
  reg [47:0] _T_463_6; // @[Switch.scala 52:30:@9397.4]
  reg [63:0] _RAND_38;
  reg [47:0] _T_463_7; // @[Switch.scala 52:30:@9397.4]
  reg [63:0] _RAND_39;
  reg [47:0] _T_463_8; // @[Switch.scala 52:30:@9397.4]
  reg [63:0] _RAND_40;
  reg [47:0] _T_463_9; // @[Switch.scala 52:30:@9397.4]
  reg [63:0] _RAND_41;
  reg [47:0] _T_463_10; // @[Switch.scala 52:30:@9397.4]
  reg [63:0] _RAND_42;
  reg [47:0] _T_463_11; // @[Switch.scala 52:30:@9397.4]
  reg [63:0] _RAND_43;
  reg [47:0] _T_463_12; // @[Switch.scala 52:30:@9397.4]
  reg [63:0] _RAND_44;
  reg [47:0] _T_463_13; // @[Switch.scala 52:30:@9397.4]
  reg [63:0] _RAND_45;
  reg [47:0] _T_463_14; // @[Switch.scala 52:30:@9397.4]
  reg [63:0] _RAND_46;
  reg [47:0] _T_463_15; // @[Switch.scala 52:30:@9397.4]
  reg [63:0] _RAND_47;
  reg [47:0] _T_463_16; // @[Switch.scala 52:30:@9397.4]
  reg [63:0] _RAND_48;
  reg [47:0] _T_463_17; // @[Switch.scala 52:30:@9397.4]
  reg [63:0] _RAND_49;
  reg [47:0] _T_463_18; // @[Switch.scala 52:30:@9397.4]
  reg [63:0] _RAND_50;
  reg [47:0] _T_463_19; // @[Switch.scala 52:30:@9397.4]
  reg [63:0] _RAND_51;
  reg [47:0] _T_463_20; // @[Switch.scala 52:30:@9397.4]
  reg [63:0] _RAND_52;
  reg [47:0] _T_463_21; // @[Switch.scala 52:30:@9397.4]
  reg [63:0] _RAND_53;
  reg [47:0] _T_463_22; // @[Switch.scala 52:30:@9397.4]
  reg [63:0] _RAND_54;
  reg [47:0] _T_463_23; // @[Switch.scala 52:30:@9397.4]
  reg [63:0] _RAND_55;
  reg [47:0] _T_463_24; // @[Switch.scala 52:30:@9397.4]
  reg [63:0] _RAND_56;
  reg [47:0] _T_463_25; // @[Switch.scala 52:30:@9397.4]
  reg [63:0] _RAND_57;
  reg [47:0] _T_463_26; // @[Switch.scala 52:30:@9397.4]
  reg [63:0] _RAND_58;
  reg [47:0] _T_463_27; // @[Switch.scala 52:30:@9397.4]
  reg [63:0] _RAND_59;
  reg [47:0] _T_463_28; // @[Switch.scala 52:30:@9397.4]
  reg [63:0] _RAND_60;
  reg [47:0] _T_463_29; // @[Switch.scala 52:30:@9397.4]
  reg [63:0] _RAND_61;
  reg [47:0] _T_463_30; // @[Switch.scala 52:30:@9397.4]
  reg [63:0] _RAND_62;
  reg [47:0] _T_463_31; // @[Switch.scala 52:30:@9397.4]
  reg [63:0] _RAND_63;
  reg  _T_632_0; // @[Switch.scala 53:31:@9462.4]
  reg [31:0] _RAND_64;
  reg  _T_632_1; // @[Switch.scala 53:31:@9462.4]
  reg [31:0] _RAND_65;
  reg  _T_632_2; // @[Switch.scala 53:31:@9462.4]
  reg [31:0] _RAND_66;
  reg  _T_632_3; // @[Switch.scala 53:31:@9462.4]
  reg [31:0] _RAND_67;
  reg  _T_632_4; // @[Switch.scala 53:31:@9462.4]
  reg [31:0] _RAND_68;
  reg  _T_632_5; // @[Switch.scala 53:31:@9462.4]
  reg [31:0] _RAND_69;
  reg  _T_632_6; // @[Switch.scala 53:31:@9462.4]
  reg [31:0] _RAND_70;
  reg  _T_632_7; // @[Switch.scala 53:31:@9462.4]
  reg [31:0] _RAND_71;
  reg  _T_632_8; // @[Switch.scala 53:31:@9462.4]
  reg [31:0] _RAND_72;
  reg  _T_632_9; // @[Switch.scala 53:31:@9462.4]
  reg [31:0] _RAND_73;
  reg  _T_632_10; // @[Switch.scala 53:31:@9462.4]
  reg [31:0] _RAND_74;
  reg  _T_632_11; // @[Switch.scala 53:31:@9462.4]
  reg [31:0] _RAND_75;
  reg  _T_632_12; // @[Switch.scala 53:31:@9462.4]
  reg [31:0] _RAND_76;
  reg  _T_632_13; // @[Switch.scala 53:31:@9462.4]
  reg [31:0] _RAND_77;
  reg  _T_632_14; // @[Switch.scala 53:31:@9462.4]
  reg [31:0] _RAND_78;
  reg  _T_632_15; // @[Switch.scala 53:31:@9462.4]
  reg [31:0] _RAND_79;
  reg  _T_632_16; // @[Switch.scala 53:31:@9462.4]
  reg [31:0] _RAND_80;
  reg  _T_632_17; // @[Switch.scala 53:31:@9462.4]
  reg [31:0] _RAND_81;
  reg  _T_632_18; // @[Switch.scala 53:31:@9462.4]
  reg [31:0] _RAND_82;
  reg  _T_632_19; // @[Switch.scala 53:31:@9462.4]
  reg [31:0] _RAND_83;
  reg  _T_632_20; // @[Switch.scala 53:31:@9462.4]
  reg [31:0] _RAND_84;
  reg  _T_632_21; // @[Switch.scala 53:31:@9462.4]
  reg [31:0] _RAND_85;
  reg  _T_632_22; // @[Switch.scala 53:31:@9462.4]
  reg [31:0] _RAND_86;
  reg  _T_632_23; // @[Switch.scala 53:31:@9462.4]
  reg [31:0] _RAND_87;
  reg  _T_632_24; // @[Switch.scala 53:31:@9462.4]
  reg [31:0] _RAND_88;
  reg  _T_632_25; // @[Switch.scala 53:31:@9462.4]
  reg [31:0] _RAND_89;
  reg  _T_632_26; // @[Switch.scala 53:31:@9462.4]
  reg [31:0] _RAND_90;
  reg  _T_632_27; // @[Switch.scala 53:31:@9462.4]
  reg [31:0] _RAND_91;
  reg  _T_632_28; // @[Switch.scala 53:31:@9462.4]
  reg [31:0] _RAND_92;
  reg  _T_632_29; // @[Switch.scala 53:31:@9462.4]
  reg [31:0] _RAND_93;
  reg  _T_632_30; // @[Switch.scala 53:31:@9462.4]
  reg [31:0] _RAND_94;
  reg  _T_632_31; // @[Switch.scala 53:31:@9462.4]
  reg [31:0] _RAND_95;
  reg  _T_801_0; // @[Switch.scala 54:23:@9527.4]
  reg [31:0] _RAND_96;
  reg  _T_801_1; // @[Switch.scala 54:23:@9527.4]
  reg [31:0] _RAND_97;
  reg  _T_801_2; // @[Switch.scala 54:23:@9527.4]
  reg [31:0] _RAND_98;
  reg  _T_801_3; // @[Switch.scala 54:23:@9527.4]
  reg [31:0] _RAND_99;
  reg  _T_801_4; // @[Switch.scala 54:23:@9527.4]
  reg [31:0] _RAND_100;
  reg  _T_801_5; // @[Switch.scala 54:23:@9527.4]
  reg [31:0] _RAND_101;
  reg  _T_801_6; // @[Switch.scala 54:23:@9527.4]
  reg [31:0] _RAND_102;
  reg  _T_801_7; // @[Switch.scala 54:23:@9527.4]
  reg [31:0] _RAND_103;
  reg  _T_801_8; // @[Switch.scala 54:23:@9527.4]
  reg [31:0] _RAND_104;
  reg  _T_801_9; // @[Switch.scala 54:23:@9527.4]
  reg [31:0] _RAND_105;
  reg  _T_801_10; // @[Switch.scala 54:23:@9527.4]
  reg [31:0] _RAND_106;
  reg  _T_801_11; // @[Switch.scala 54:23:@9527.4]
  reg [31:0] _RAND_107;
  reg  _T_801_12; // @[Switch.scala 54:23:@9527.4]
  reg [31:0] _RAND_108;
  reg  _T_801_13; // @[Switch.scala 54:23:@9527.4]
  reg [31:0] _RAND_109;
  reg  _T_801_14; // @[Switch.scala 54:23:@9527.4]
  reg [31:0] _RAND_110;
  reg  _T_801_15; // @[Switch.scala 54:23:@9527.4]
  reg [31:0] _RAND_111;
  reg  _T_801_16; // @[Switch.scala 54:23:@9527.4]
  reg [31:0] _RAND_112;
  reg  _T_801_17; // @[Switch.scala 54:23:@9527.4]
  reg [31:0] _RAND_113;
  reg  _T_801_18; // @[Switch.scala 54:23:@9527.4]
  reg [31:0] _RAND_114;
  reg  _T_801_19; // @[Switch.scala 54:23:@9527.4]
  reg [31:0] _RAND_115;
  reg  _T_801_20; // @[Switch.scala 54:23:@9527.4]
  reg [31:0] _RAND_116;
  reg  _T_801_21; // @[Switch.scala 54:23:@9527.4]
  reg [31:0] _RAND_117;
  reg  _T_801_22; // @[Switch.scala 54:23:@9527.4]
  reg [31:0] _RAND_118;
  reg  _T_801_23; // @[Switch.scala 54:23:@9527.4]
  reg [31:0] _RAND_119;
  reg  _T_801_24; // @[Switch.scala 54:23:@9527.4]
  reg [31:0] _RAND_120;
  reg  _T_801_25; // @[Switch.scala 54:23:@9527.4]
  reg [31:0] _RAND_121;
  reg  _T_801_26; // @[Switch.scala 54:23:@9527.4]
  reg [31:0] _RAND_122;
  reg  _T_801_27; // @[Switch.scala 54:23:@9527.4]
  reg [31:0] _RAND_123;
  reg  _T_801_28; // @[Switch.scala 54:23:@9527.4]
  reg [31:0] _RAND_124;
  reg  _T_801_29; // @[Switch.scala 54:23:@9527.4]
  reg [31:0] _RAND_125;
  reg  _T_801_30; // @[Switch.scala 54:23:@9527.4]
  reg [31:0] _RAND_126;
  reg  _T_801_31; // @[Switch.scala 54:23:@9527.4]
  reg [31:0] _RAND_127;
  reg [47:0] _T_970_0; // @[Switch.scala 55:24:@9592.4]
  reg [63:0] _RAND_128;
  reg [47:0] _T_970_1; // @[Switch.scala 55:24:@9592.4]
  reg [63:0] _RAND_129;
  reg [47:0] _T_970_2; // @[Switch.scala 55:24:@9592.4]
  reg [63:0] _RAND_130;
  reg [47:0] _T_970_3; // @[Switch.scala 55:24:@9592.4]
  reg [63:0] _RAND_131;
  reg [47:0] _T_970_4; // @[Switch.scala 55:24:@9592.4]
  reg [63:0] _RAND_132;
  reg [47:0] _T_970_5; // @[Switch.scala 55:24:@9592.4]
  reg [63:0] _RAND_133;
  reg [47:0] _T_970_6; // @[Switch.scala 55:24:@9592.4]
  reg [63:0] _RAND_134;
  reg [47:0] _T_970_7; // @[Switch.scala 55:24:@9592.4]
  reg [63:0] _RAND_135;
  reg [47:0] _T_970_8; // @[Switch.scala 55:24:@9592.4]
  reg [63:0] _RAND_136;
  reg [47:0] _T_970_9; // @[Switch.scala 55:24:@9592.4]
  reg [63:0] _RAND_137;
  reg [47:0] _T_970_10; // @[Switch.scala 55:24:@9592.4]
  reg [63:0] _RAND_138;
  reg [47:0] _T_970_11; // @[Switch.scala 55:24:@9592.4]
  reg [63:0] _RAND_139;
  reg [47:0] _T_970_12; // @[Switch.scala 55:24:@9592.4]
  reg [63:0] _RAND_140;
  reg [47:0] _T_970_13; // @[Switch.scala 55:24:@9592.4]
  reg [63:0] _RAND_141;
  reg [47:0] _T_970_14; // @[Switch.scala 55:24:@9592.4]
  reg [63:0] _RAND_142;
  reg [47:0] _T_970_15; // @[Switch.scala 55:24:@9592.4]
  reg [63:0] _RAND_143;
  reg [47:0] _T_970_16; // @[Switch.scala 55:24:@9592.4]
  reg [63:0] _RAND_144;
  reg [47:0] _T_970_17; // @[Switch.scala 55:24:@9592.4]
  reg [63:0] _RAND_145;
  reg [47:0] _T_970_18; // @[Switch.scala 55:24:@9592.4]
  reg [63:0] _RAND_146;
  reg [47:0] _T_970_19; // @[Switch.scala 55:24:@9592.4]
  reg [63:0] _RAND_147;
  reg [47:0] _T_970_20; // @[Switch.scala 55:24:@9592.4]
  reg [63:0] _RAND_148;
  reg [47:0] _T_970_21; // @[Switch.scala 55:24:@9592.4]
  reg [63:0] _RAND_149;
  reg [47:0] _T_970_22; // @[Switch.scala 55:24:@9592.4]
  reg [63:0] _RAND_150;
  reg [47:0] _T_970_23; // @[Switch.scala 55:24:@9592.4]
  reg [63:0] _RAND_151;
  reg [47:0] _T_970_24; // @[Switch.scala 55:24:@9592.4]
  reg [63:0] _RAND_152;
  reg [47:0] _T_970_25; // @[Switch.scala 55:24:@9592.4]
  reg [63:0] _RAND_153;
  reg [47:0] _T_970_26; // @[Switch.scala 55:24:@9592.4]
  reg [63:0] _RAND_154;
  reg [47:0] _T_970_27; // @[Switch.scala 55:24:@9592.4]
  reg [63:0] _RAND_155;
  reg [47:0] _T_970_28; // @[Switch.scala 55:24:@9592.4]
  reg [63:0] _RAND_156;
  reg [47:0] _T_970_29; // @[Switch.scala 55:24:@9592.4]
  reg [63:0] _RAND_157;
  reg [47:0] _T_970_30; // @[Switch.scala 55:24:@9592.4]
  reg [63:0] _RAND_158;
  reg [47:0] _T_970_31; // @[Switch.scala 55:24:@9592.4]
  reg [63:0] _RAND_159;
  reg  _T_1139_0; // @[Switch.scala 56:25:@9657.4]
  reg [31:0] _RAND_160;
  reg  _T_1139_1; // @[Switch.scala 56:25:@9657.4]
  reg [31:0] _RAND_161;
  reg  _T_1139_2; // @[Switch.scala 56:25:@9657.4]
  reg [31:0] _RAND_162;
  reg  _T_1139_3; // @[Switch.scala 56:25:@9657.4]
  reg [31:0] _RAND_163;
  reg  _T_1139_4; // @[Switch.scala 56:25:@9657.4]
  reg [31:0] _RAND_164;
  reg  _T_1139_5; // @[Switch.scala 56:25:@9657.4]
  reg [31:0] _RAND_165;
  reg  _T_1139_6; // @[Switch.scala 56:25:@9657.4]
  reg [31:0] _RAND_166;
  reg  _T_1139_7; // @[Switch.scala 56:25:@9657.4]
  reg [31:0] _RAND_167;
  reg  _T_1139_8; // @[Switch.scala 56:25:@9657.4]
  reg [31:0] _RAND_168;
  reg  _T_1139_9; // @[Switch.scala 56:25:@9657.4]
  reg [31:0] _RAND_169;
  reg  _T_1139_10; // @[Switch.scala 56:25:@9657.4]
  reg [31:0] _RAND_170;
  reg  _T_1139_11; // @[Switch.scala 56:25:@9657.4]
  reg [31:0] _RAND_171;
  reg  _T_1139_12; // @[Switch.scala 56:25:@9657.4]
  reg [31:0] _RAND_172;
  reg  _T_1139_13; // @[Switch.scala 56:25:@9657.4]
  reg [31:0] _RAND_173;
  reg  _T_1139_14; // @[Switch.scala 56:25:@9657.4]
  reg [31:0] _RAND_174;
  reg  _T_1139_15; // @[Switch.scala 56:25:@9657.4]
  reg [31:0] _RAND_175;
  reg  _T_1139_16; // @[Switch.scala 56:25:@9657.4]
  reg [31:0] _RAND_176;
  reg  _T_1139_17; // @[Switch.scala 56:25:@9657.4]
  reg [31:0] _RAND_177;
  reg  _T_1139_18; // @[Switch.scala 56:25:@9657.4]
  reg [31:0] _RAND_178;
  reg  _T_1139_19; // @[Switch.scala 56:25:@9657.4]
  reg [31:0] _RAND_179;
  reg  _T_1139_20; // @[Switch.scala 56:25:@9657.4]
  reg [31:0] _RAND_180;
  reg  _T_1139_21; // @[Switch.scala 56:25:@9657.4]
  reg [31:0] _RAND_181;
  reg  _T_1139_22; // @[Switch.scala 56:25:@9657.4]
  reg [31:0] _RAND_182;
  reg  _T_1139_23; // @[Switch.scala 56:25:@9657.4]
  reg [31:0] _RAND_183;
  reg  _T_1139_24; // @[Switch.scala 56:25:@9657.4]
  reg [31:0] _RAND_184;
  reg  _T_1139_25; // @[Switch.scala 56:25:@9657.4]
  reg [31:0] _RAND_185;
  reg  _T_1139_26; // @[Switch.scala 56:25:@9657.4]
  reg [31:0] _RAND_186;
  reg  _T_1139_27; // @[Switch.scala 56:25:@9657.4]
  reg [31:0] _RAND_187;
  reg  _T_1139_28; // @[Switch.scala 56:25:@9657.4]
  reg [31:0] _RAND_188;
  reg  _T_1139_29; // @[Switch.scala 56:25:@9657.4]
  reg [31:0] _RAND_189;
  reg  _T_1139_30; // @[Switch.scala 56:25:@9657.4]
  reg [31:0] _RAND_190;
  reg  _T_1139_31; // @[Switch.scala 56:25:@9657.4]
  reg [31:0] _RAND_191;
  Switch switch ( // @[Switch.scala 50:22:@9329.4]
    .io_inAddr_0(switch_io_inAddr_0),
    .io_inAddr_1(switch_io_inAddr_1),
    .io_inAddr_2(switch_io_inAddr_2),
    .io_inAddr_3(switch_io_inAddr_3),
    .io_inAddr_4(switch_io_inAddr_4),
    .io_inAddr_5(switch_io_inAddr_5),
    .io_inAddr_6(switch_io_inAddr_6),
    .io_inAddr_7(switch_io_inAddr_7),
    .io_inAddr_8(switch_io_inAddr_8),
    .io_inAddr_9(switch_io_inAddr_9),
    .io_inAddr_10(switch_io_inAddr_10),
    .io_inAddr_11(switch_io_inAddr_11),
    .io_inAddr_12(switch_io_inAddr_12),
    .io_inAddr_13(switch_io_inAddr_13),
    .io_inAddr_14(switch_io_inAddr_14),
    .io_inAddr_15(switch_io_inAddr_15),
    .io_inAddr_16(switch_io_inAddr_16),
    .io_inAddr_17(switch_io_inAddr_17),
    .io_inAddr_18(switch_io_inAddr_18),
    .io_inAddr_19(switch_io_inAddr_19),
    .io_inAddr_20(switch_io_inAddr_20),
    .io_inAddr_21(switch_io_inAddr_21),
    .io_inAddr_22(switch_io_inAddr_22),
    .io_inAddr_23(switch_io_inAddr_23),
    .io_inAddr_24(switch_io_inAddr_24),
    .io_inAddr_25(switch_io_inAddr_25),
    .io_inAddr_26(switch_io_inAddr_26),
    .io_inAddr_27(switch_io_inAddr_27),
    .io_inAddr_28(switch_io_inAddr_28),
    .io_inAddr_29(switch_io_inAddr_29),
    .io_inAddr_30(switch_io_inAddr_30),
    .io_inAddr_31(switch_io_inAddr_31),
    .io_inData_0(switch_io_inData_0),
    .io_inData_1(switch_io_inData_1),
    .io_inData_2(switch_io_inData_2),
    .io_inData_3(switch_io_inData_3),
    .io_inData_4(switch_io_inData_4),
    .io_inData_5(switch_io_inData_5),
    .io_inData_6(switch_io_inData_6),
    .io_inData_7(switch_io_inData_7),
    .io_inData_8(switch_io_inData_8),
    .io_inData_9(switch_io_inData_9),
    .io_inData_10(switch_io_inData_10),
    .io_inData_11(switch_io_inData_11),
    .io_inData_12(switch_io_inData_12),
    .io_inData_13(switch_io_inData_13),
    .io_inData_14(switch_io_inData_14),
    .io_inData_15(switch_io_inData_15),
    .io_inData_16(switch_io_inData_16),
    .io_inData_17(switch_io_inData_17),
    .io_inData_18(switch_io_inData_18),
    .io_inData_19(switch_io_inData_19),
    .io_inData_20(switch_io_inData_20),
    .io_inData_21(switch_io_inData_21),
    .io_inData_22(switch_io_inData_22),
    .io_inData_23(switch_io_inData_23),
    .io_inData_24(switch_io_inData_24),
    .io_inData_25(switch_io_inData_25),
    .io_inData_26(switch_io_inData_26),
    .io_inData_27(switch_io_inData_27),
    .io_inData_28(switch_io_inData_28),
    .io_inData_29(switch_io_inData_29),
    .io_inData_30(switch_io_inData_30),
    .io_inData_31(switch_io_inData_31),
    .io_inValid_0(switch_io_inValid_0),
    .io_inValid_1(switch_io_inValid_1),
    .io_inValid_2(switch_io_inValid_2),
    .io_inValid_3(switch_io_inValid_3),
    .io_inValid_4(switch_io_inValid_4),
    .io_inValid_5(switch_io_inValid_5),
    .io_inValid_6(switch_io_inValid_6),
    .io_inValid_7(switch_io_inValid_7),
    .io_inValid_8(switch_io_inValid_8),
    .io_inValid_9(switch_io_inValid_9),
    .io_inValid_10(switch_io_inValid_10),
    .io_inValid_11(switch_io_inValid_11),
    .io_inValid_12(switch_io_inValid_12),
    .io_inValid_13(switch_io_inValid_13),
    .io_inValid_14(switch_io_inValid_14),
    .io_inValid_15(switch_io_inValid_15),
    .io_inValid_16(switch_io_inValid_16),
    .io_inValid_17(switch_io_inValid_17),
    .io_inValid_18(switch_io_inValid_18),
    .io_inValid_19(switch_io_inValid_19),
    .io_inValid_20(switch_io_inValid_20),
    .io_inValid_21(switch_io_inValid_21),
    .io_inValid_22(switch_io_inValid_22),
    .io_inValid_23(switch_io_inValid_23),
    .io_inValid_24(switch_io_inValid_24),
    .io_inValid_25(switch_io_inValid_25),
    .io_inValid_26(switch_io_inValid_26),
    .io_inValid_27(switch_io_inValid_27),
    .io_inValid_28(switch_io_inValid_28),
    .io_inValid_29(switch_io_inValid_29),
    .io_inValid_30(switch_io_inValid_30),
    .io_inValid_31(switch_io_inValid_31),
    .io_outAck_0(switch_io_outAck_0),
    .io_outAck_1(switch_io_outAck_1),
    .io_outAck_2(switch_io_outAck_2),
    .io_outAck_3(switch_io_outAck_3),
    .io_outAck_4(switch_io_outAck_4),
    .io_outAck_5(switch_io_outAck_5),
    .io_outAck_6(switch_io_outAck_6),
    .io_outAck_7(switch_io_outAck_7),
    .io_outAck_8(switch_io_outAck_8),
    .io_outAck_9(switch_io_outAck_9),
    .io_outAck_10(switch_io_outAck_10),
    .io_outAck_11(switch_io_outAck_11),
    .io_outAck_12(switch_io_outAck_12),
    .io_outAck_13(switch_io_outAck_13),
    .io_outAck_14(switch_io_outAck_14),
    .io_outAck_15(switch_io_outAck_15),
    .io_outAck_16(switch_io_outAck_16),
    .io_outAck_17(switch_io_outAck_17),
    .io_outAck_18(switch_io_outAck_18),
    .io_outAck_19(switch_io_outAck_19),
    .io_outAck_20(switch_io_outAck_20),
    .io_outAck_21(switch_io_outAck_21),
    .io_outAck_22(switch_io_outAck_22),
    .io_outAck_23(switch_io_outAck_23),
    .io_outAck_24(switch_io_outAck_24),
    .io_outAck_25(switch_io_outAck_25),
    .io_outAck_26(switch_io_outAck_26),
    .io_outAck_27(switch_io_outAck_27),
    .io_outAck_28(switch_io_outAck_28),
    .io_outAck_29(switch_io_outAck_29),
    .io_outAck_30(switch_io_outAck_30),
    .io_outAck_31(switch_io_outAck_31),
    .io_outData_0(switch_io_outData_0),
    .io_outData_1(switch_io_outData_1),
    .io_outData_2(switch_io_outData_2),
    .io_outData_3(switch_io_outData_3),
    .io_outData_4(switch_io_outData_4),
    .io_outData_5(switch_io_outData_5),
    .io_outData_6(switch_io_outData_6),
    .io_outData_7(switch_io_outData_7),
    .io_outData_8(switch_io_outData_8),
    .io_outData_9(switch_io_outData_9),
    .io_outData_10(switch_io_outData_10),
    .io_outData_11(switch_io_outData_11),
    .io_outData_12(switch_io_outData_12),
    .io_outData_13(switch_io_outData_13),
    .io_outData_14(switch_io_outData_14),
    .io_outData_15(switch_io_outData_15),
    .io_outData_16(switch_io_outData_16),
    .io_outData_17(switch_io_outData_17),
    .io_outData_18(switch_io_outData_18),
    .io_outData_19(switch_io_outData_19),
    .io_outData_20(switch_io_outData_20),
    .io_outData_21(switch_io_outData_21),
    .io_outData_22(switch_io_outData_22),
    .io_outData_23(switch_io_outData_23),
    .io_outData_24(switch_io_outData_24),
    .io_outData_25(switch_io_outData_25),
    .io_outData_26(switch_io_outData_26),
    .io_outData_27(switch_io_outData_27),
    .io_outData_28(switch_io_outData_28),
    .io_outData_29(switch_io_outData_29),
    .io_outData_30(switch_io_outData_30),
    .io_outData_31(switch_io_outData_31),
    .io_outValid_0(switch_io_outValid_0),
    .io_outValid_1(switch_io_outValid_1),
    .io_outValid_2(switch_io_outValid_2),
    .io_outValid_3(switch_io_outValid_3),
    .io_outValid_4(switch_io_outValid_4),
    .io_outValid_5(switch_io_outValid_5),
    .io_outValid_6(switch_io_outValid_6),
    .io_outValid_7(switch_io_outValid_7),
    .io_outValid_8(switch_io_outValid_8),
    .io_outValid_9(switch_io_outValid_9),
    .io_outValid_10(switch_io_outValid_10),
    .io_outValid_11(switch_io_outValid_11),
    .io_outValid_12(switch_io_outValid_12),
    .io_outValid_13(switch_io_outValid_13),
    .io_outValid_14(switch_io_outValid_14),
    .io_outValid_15(switch_io_outValid_15),
    .io_outValid_16(switch_io_outValid_16),
    .io_outValid_17(switch_io_outValid_17),
    .io_outValid_18(switch_io_outValid_18),
    .io_outValid_19(switch_io_outValid_19),
    .io_outValid_20(switch_io_outValid_20),
    .io_outValid_21(switch_io_outValid_21),
    .io_outValid_22(switch_io_outValid_22),
    .io_outValid_23(switch_io_outValid_23),
    .io_outValid_24(switch_io_outValid_24),
    .io_outValid_25(switch_io_outValid_25),
    .io_outValid_26(switch_io_outValid_26),
    .io_outValid_27(switch_io_outValid_27),
    .io_outValid_28(switch_io_outValid_28),
    .io_outValid_29(switch_io_outValid_29),
    .io_outValid_30(switch_io_outValid_30),
    .io_outValid_31(switch_io_outValid_31)
  );
  assign io_outAck_0 = _T_801_0; // @[Switch.scala 54:13:@9560.4]
  assign io_outAck_1 = _T_801_1; // @[Switch.scala 54:13:@9561.4]
  assign io_outAck_2 = _T_801_2; // @[Switch.scala 54:13:@9562.4]
  assign io_outAck_3 = _T_801_3; // @[Switch.scala 54:13:@9563.4]
  assign io_outAck_4 = _T_801_4; // @[Switch.scala 54:13:@9564.4]
  assign io_outAck_5 = _T_801_5; // @[Switch.scala 54:13:@9565.4]
  assign io_outAck_6 = _T_801_6; // @[Switch.scala 54:13:@9566.4]
  assign io_outAck_7 = _T_801_7; // @[Switch.scala 54:13:@9567.4]
  assign io_outAck_8 = _T_801_8; // @[Switch.scala 54:13:@9568.4]
  assign io_outAck_9 = _T_801_9; // @[Switch.scala 54:13:@9569.4]
  assign io_outAck_10 = _T_801_10; // @[Switch.scala 54:13:@9570.4]
  assign io_outAck_11 = _T_801_11; // @[Switch.scala 54:13:@9571.4]
  assign io_outAck_12 = _T_801_12; // @[Switch.scala 54:13:@9572.4]
  assign io_outAck_13 = _T_801_13; // @[Switch.scala 54:13:@9573.4]
  assign io_outAck_14 = _T_801_14; // @[Switch.scala 54:13:@9574.4]
  assign io_outAck_15 = _T_801_15; // @[Switch.scala 54:13:@9575.4]
  assign io_outAck_16 = _T_801_16; // @[Switch.scala 54:13:@9576.4]
  assign io_outAck_17 = _T_801_17; // @[Switch.scala 54:13:@9577.4]
  assign io_outAck_18 = _T_801_18; // @[Switch.scala 54:13:@9578.4]
  assign io_outAck_19 = _T_801_19; // @[Switch.scala 54:13:@9579.4]
  assign io_outAck_20 = _T_801_20; // @[Switch.scala 54:13:@9580.4]
  assign io_outAck_21 = _T_801_21; // @[Switch.scala 54:13:@9581.4]
  assign io_outAck_22 = _T_801_22; // @[Switch.scala 54:13:@9582.4]
  assign io_outAck_23 = _T_801_23; // @[Switch.scala 54:13:@9583.4]
  assign io_outAck_24 = _T_801_24; // @[Switch.scala 54:13:@9584.4]
  assign io_outAck_25 = _T_801_25; // @[Switch.scala 54:13:@9585.4]
  assign io_outAck_26 = _T_801_26; // @[Switch.scala 54:13:@9586.4]
  assign io_outAck_27 = _T_801_27; // @[Switch.scala 54:13:@9587.4]
  assign io_outAck_28 = _T_801_28; // @[Switch.scala 54:13:@9588.4]
  assign io_outAck_29 = _T_801_29; // @[Switch.scala 54:13:@9589.4]
  assign io_outAck_30 = _T_801_30; // @[Switch.scala 54:13:@9590.4]
  assign io_outAck_31 = _T_801_31; // @[Switch.scala 54:13:@9591.4]
  assign io_outData_0 = _T_970_0; // @[Switch.scala 55:14:@9625.4]
  assign io_outData_1 = _T_970_1; // @[Switch.scala 55:14:@9626.4]
  assign io_outData_2 = _T_970_2; // @[Switch.scala 55:14:@9627.4]
  assign io_outData_3 = _T_970_3; // @[Switch.scala 55:14:@9628.4]
  assign io_outData_4 = _T_970_4; // @[Switch.scala 55:14:@9629.4]
  assign io_outData_5 = _T_970_5; // @[Switch.scala 55:14:@9630.4]
  assign io_outData_6 = _T_970_6; // @[Switch.scala 55:14:@9631.4]
  assign io_outData_7 = _T_970_7; // @[Switch.scala 55:14:@9632.4]
  assign io_outData_8 = _T_970_8; // @[Switch.scala 55:14:@9633.4]
  assign io_outData_9 = _T_970_9; // @[Switch.scala 55:14:@9634.4]
  assign io_outData_10 = _T_970_10; // @[Switch.scala 55:14:@9635.4]
  assign io_outData_11 = _T_970_11; // @[Switch.scala 55:14:@9636.4]
  assign io_outData_12 = _T_970_12; // @[Switch.scala 55:14:@9637.4]
  assign io_outData_13 = _T_970_13; // @[Switch.scala 55:14:@9638.4]
  assign io_outData_14 = _T_970_14; // @[Switch.scala 55:14:@9639.4]
  assign io_outData_15 = _T_970_15; // @[Switch.scala 55:14:@9640.4]
  assign io_outData_16 = _T_970_16; // @[Switch.scala 55:14:@9641.4]
  assign io_outData_17 = _T_970_17; // @[Switch.scala 55:14:@9642.4]
  assign io_outData_18 = _T_970_18; // @[Switch.scala 55:14:@9643.4]
  assign io_outData_19 = _T_970_19; // @[Switch.scala 55:14:@9644.4]
  assign io_outData_20 = _T_970_20; // @[Switch.scala 55:14:@9645.4]
  assign io_outData_21 = _T_970_21; // @[Switch.scala 55:14:@9646.4]
  assign io_outData_22 = _T_970_22; // @[Switch.scala 55:14:@9647.4]
  assign io_outData_23 = _T_970_23; // @[Switch.scala 55:14:@9648.4]
  assign io_outData_24 = _T_970_24; // @[Switch.scala 55:14:@9649.4]
  assign io_outData_25 = _T_970_25; // @[Switch.scala 55:14:@9650.4]
  assign io_outData_26 = _T_970_26; // @[Switch.scala 55:14:@9651.4]
  assign io_outData_27 = _T_970_27; // @[Switch.scala 55:14:@9652.4]
  assign io_outData_28 = _T_970_28; // @[Switch.scala 55:14:@9653.4]
  assign io_outData_29 = _T_970_29; // @[Switch.scala 55:14:@9654.4]
  assign io_outData_30 = _T_970_30; // @[Switch.scala 55:14:@9655.4]
  assign io_outData_31 = _T_970_31; // @[Switch.scala 55:14:@9656.4]
  assign io_outValid_0 = _T_1139_0; // @[Switch.scala 56:15:@9690.4]
  assign io_outValid_1 = _T_1139_1; // @[Switch.scala 56:15:@9691.4]
  assign io_outValid_2 = _T_1139_2; // @[Switch.scala 56:15:@9692.4]
  assign io_outValid_3 = _T_1139_3; // @[Switch.scala 56:15:@9693.4]
  assign io_outValid_4 = _T_1139_4; // @[Switch.scala 56:15:@9694.4]
  assign io_outValid_5 = _T_1139_5; // @[Switch.scala 56:15:@9695.4]
  assign io_outValid_6 = _T_1139_6; // @[Switch.scala 56:15:@9696.4]
  assign io_outValid_7 = _T_1139_7; // @[Switch.scala 56:15:@9697.4]
  assign io_outValid_8 = _T_1139_8; // @[Switch.scala 56:15:@9698.4]
  assign io_outValid_9 = _T_1139_9; // @[Switch.scala 56:15:@9699.4]
  assign io_outValid_10 = _T_1139_10; // @[Switch.scala 56:15:@9700.4]
  assign io_outValid_11 = _T_1139_11; // @[Switch.scala 56:15:@9701.4]
  assign io_outValid_12 = _T_1139_12; // @[Switch.scala 56:15:@9702.4]
  assign io_outValid_13 = _T_1139_13; // @[Switch.scala 56:15:@9703.4]
  assign io_outValid_14 = _T_1139_14; // @[Switch.scala 56:15:@9704.4]
  assign io_outValid_15 = _T_1139_15; // @[Switch.scala 56:15:@9705.4]
  assign io_outValid_16 = _T_1139_16; // @[Switch.scala 56:15:@9706.4]
  assign io_outValid_17 = _T_1139_17; // @[Switch.scala 56:15:@9707.4]
  assign io_outValid_18 = _T_1139_18; // @[Switch.scala 56:15:@9708.4]
  assign io_outValid_19 = _T_1139_19; // @[Switch.scala 56:15:@9709.4]
  assign io_outValid_20 = _T_1139_20; // @[Switch.scala 56:15:@9710.4]
  assign io_outValid_21 = _T_1139_21; // @[Switch.scala 56:15:@9711.4]
  assign io_outValid_22 = _T_1139_22; // @[Switch.scala 56:15:@9712.4]
  assign io_outValid_23 = _T_1139_23; // @[Switch.scala 56:15:@9713.4]
  assign io_outValid_24 = _T_1139_24; // @[Switch.scala 56:15:@9714.4]
  assign io_outValid_25 = _T_1139_25; // @[Switch.scala 56:15:@9715.4]
  assign io_outValid_26 = _T_1139_26; // @[Switch.scala 56:15:@9716.4]
  assign io_outValid_27 = _T_1139_27; // @[Switch.scala 56:15:@9717.4]
  assign io_outValid_28 = _T_1139_28; // @[Switch.scala 56:15:@9718.4]
  assign io_outValid_29 = _T_1139_29; // @[Switch.scala 56:15:@9719.4]
  assign io_outValid_30 = _T_1139_30; // @[Switch.scala 56:15:@9720.4]
  assign io_outValid_31 = _T_1139_31; // @[Switch.scala 56:15:@9721.4]
  assign switch_io_inAddr_0 = _T_294_0; // @[Switch.scala 51:20:@9365.4]
  assign switch_io_inAddr_1 = _T_294_1; // @[Switch.scala 51:20:@9366.4]
  assign switch_io_inAddr_2 = _T_294_2; // @[Switch.scala 51:20:@9367.4]
  assign switch_io_inAddr_3 = _T_294_3; // @[Switch.scala 51:20:@9368.4]
  assign switch_io_inAddr_4 = _T_294_4; // @[Switch.scala 51:20:@9369.4]
  assign switch_io_inAddr_5 = _T_294_5; // @[Switch.scala 51:20:@9370.4]
  assign switch_io_inAddr_6 = _T_294_6; // @[Switch.scala 51:20:@9371.4]
  assign switch_io_inAddr_7 = _T_294_7; // @[Switch.scala 51:20:@9372.4]
  assign switch_io_inAddr_8 = _T_294_8; // @[Switch.scala 51:20:@9373.4]
  assign switch_io_inAddr_9 = _T_294_9; // @[Switch.scala 51:20:@9374.4]
  assign switch_io_inAddr_10 = _T_294_10; // @[Switch.scala 51:20:@9375.4]
  assign switch_io_inAddr_11 = _T_294_11; // @[Switch.scala 51:20:@9376.4]
  assign switch_io_inAddr_12 = _T_294_12; // @[Switch.scala 51:20:@9377.4]
  assign switch_io_inAddr_13 = _T_294_13; // @[Switch.scala 51:20:@9378.4]
  assign switch_io_inAddr_14 = _T_294_14; // @[Switch.scala 51:20:@9379.4]
  assign switch_io_inAddr_15 = _T_294_15; // @[Switch.scala 51:20:@9380.4]
  assign switch_io_inAddr_16 = _T_294_16; // @[Switch.scala 51:20:@9381.4]
  assign switch_io_inAddr_17 = _T_294_17; // @[Switch.scala 51:20:@9382.4]
  assign switch_io_inAddr_18 = _T_294_18; // @[Switch.scala 51:20:@9383.4]
  assign switch_io_inAddr_19 = _T_294_19; // @[Switch.scala 51:20:@9384.4]
  assign switch_io_inAddr_20 = _T_294_20; // @[Switch.scala 51:20:@9385.4]
  assign switch_io_inAddr_21 = _T_294_21; // @[Switch.scala 51:20:@9386.4]
  assign switch_io_inAddr_22 = _T_294_22; // @[Switch.scala 51:20:@9387.4]
  assign switch_io_inAddr_23 = _T_294_23; // @[Switch.scala 51:20:@9388.4]
  assign switch_io_inAddr_24 = _T_294_24; // @[Switch.scala 51:20:@9389.4]
  assign switch_io_inAddr_25 = _T_294_25; // @[Switch.scala 51:20:@9390.4]
  assign switch_io_inAddr_26 = _T_294_26; // @[Switch.scala 51:20:@9391.4]
  assign switch_io_inAddr_27 = _T_294_27; // @[Switch.scala 51:20:@9392.4]
  assign switch_io_inAddr_28 = _T_294_28; // @[Switch.scala 51:20:@9393.4]
  assign switch_io_inAddr_29 = _T_294_29; // @[Switch.scala 51:20:@9394.4]
  assign switch_io_inAddr_30 = _T_294_30; // @[Switch.scala 51:20:@9395.4]
  assign switch_io_inAddr_31 = _T_294_31; // @[Switch.scala 51:20:@9396.4]
  assign switch_io_inData_0 = _T_463_0; // @[Switch.scala 52:20:@9430.4]
  assign switch_io_inData_1 = _T_463_1; // @[Switch.scala 52:20:@9431.4]
  assign switch_io_inData_2 = _T_463_2; // @[Switch.scala 52:20:@9432.4]
  assign switch_io_inData_3 = _T_463_3; // @[Switch.scala 52:20:@9433.4]
  assign switch_io_inData_4 = _T_463_4; // @[Switch.scala 52:20:@9434.4]
  assign switch_io_inData_5 = _T_463_5; // @[Switch.scala 52:20:@9435.4]
  assign switch_io_inData_6 = _T_463_6; // @[Switch.scala 52:20:@9436.4]
  assign switch_io_inData_7 = _T_463_7; // @[Switch.scala 52:20:@9437.4]
  assign switch_io_inData_8 = _T_463_8; // @[Switch.scala 52:20:@9438.4]
  assign switch_io_inData_9 = _T_463_9; // @[Switch.scala 52:20:@9439.4]
  assign switch_io_inData_10 = _T_463_10; // @[Switch.scala 52:20:@9440.4]
  assign switch_io_inData_11 = _T_463_11; // @[Switch.scala 52:20:@9441.4]
  assign switch_io_inData_12 = _T_463_12; // @[Switch.scala 52:20:@9442.4]
  assign switch_io_inData_13 = _T_463_13; // @[Switch.scala 52:20:@9443.4]
  assign switch_io_inData_14 = _T_463_14; // @[Switch.scala 52:20:@9444.4]
  assign switch_io_inData_15 = _T_463_15; // @[Switch.scala 52:20:@9445.4]
  assign switch_io_inData_16 = _T_463_16; // @[Switch.scala 52:20:@9446.4]
  assign switch_io_inData_17 = _T_463_17; // @[Switch.scala 52:20:@9447.4]
  assign switch_io_inData_18 = _T_463_18; // @[Switch.scala 52:20:@9448.4]
  assign switch_io_inData_19 = _T_463_19; // @[Switch.scala 52:20:@9449.4]
  assign switch_io_inData_20 = _T_463_20; // @[Switch.scala 52:20:@9450.4]
  assign switch_io_inData_21 = _T_463_21; // @[Switch.scala 52:20:@9451.4]
  assign switch_io_inData_22 = _T_463_22; // @[Switch.scala 52:20:@9452.4]
  assign switch_io_inData_23 = _T_463_23; // @[Switch.scala 52:20:@9453.4]
  assign switch_io_inData_24 = _T_463_24; // @[Switch.scala 52:20:@9454.4]
  assign switch_io_inData_25 = _T_463_25; // @[Switch.scala 52:20:@9455.4]
  assign switch_io_inData_26 = _T_463_26; // @[Switch.scala 52:20:@9456.4]
  assign switch_io_inData_27 = _T_463_27; // @[Switch.scala 52:20:@9457.4]
  assign switch_io_inData_28 = _T_463_28; // @[Switch.scala 52:20:@9458.4]
  assign switch_io_inData_29 = _T_463_29; // @[Switch.scala 52:20:@9459.4]
  assign switch_io_inData_30 = _T_463_30; // @[Switch.scala 52:20:@9460.4]
  assign switch_io_inData_31 = _T_463_31; // @[Switch.scala 52:20:@9461.4]
  assign switch_io_inValid_0 = _T_632_0; // @[Switch.scala 53:21:@9495.4]
  assign switch_io_inValid_1 = _T_632_1; // @[Switch.scala 53:21:@9496.4]
  assign switch_io_inValid_2 = _T_632_2; // @[Switch.scala 53:21:@9497.4]
  assign switch_io_inValid_3 = _T_632_3; // @[Switch.scala 53:21:@9498.4]
  assign switch_io_inValid_4 = _T_632_4; // @[Switch.scala 53:21:@9499.4]
  assign switch_io_inValid_5 = _T_632_5; // @[Switch.scala 53:21:@9500.4]
  assign switch_io_inValid_6 = _T_632_6; // @[Switch.scala 53:21:@9501.4]
  assign switch_io_inValid_7 = _T_632_7; // @[Switch.scala 53:21:@9502.4]
  assign switch_io_inValid_8 = _T_632_8; // @[Switch.scala 53:21:@9503.4]
  assign switch_io_inValid_9 = _T_632_9; // @[Switch.scala 53:21:@9504.4]
  assign switch_io_inValid_10 = _T_632_10; // @[Switch.scala 53:21:@9505.4]
  assign switch_io_inValid_11 = _T_632_11; // @[Switch.scala 53:21:@9506.4]
  assign switch_io_inValid_12 = _T_632_12; // @[Switch.scala 53:21:@9507.4]
  assign switch_io_inValid_13 = _T_632_13; // @[Switch.scala 53:21:@9508.4]
  assign switch_io_inValid_14 = _T_632_14; // @[Switch.scala 53:21:@9509.4]
  assign switch_io_inValid_15 = _T_632_15; // @[Switch.scala 53:21:@9510.4]
  assign switch_io_inValid_16 = _T_632_16; // @[Switch.scala 53:21:@9511.4]
  assign switch_io_inValid_17 = _T_632_17; // @[Switch.scala 53:21:@9512.4]
  assign switch_io_inValid_18 = _T_632_18; // @[Switch.scala 53:21:@9513.4]
  assign switch_io_inValid_19 = _T_632_19; // @[Switch.scala 53:21:@9514.4]
  assign switch_io_inValid_20 = _T_632_20; // @[Switch.scala 53:21:@9515.4]
  assign switch_io_inValid_21 = _T_632_21; // @[Switch.scala 53:21:@9516.4]
  assign switch_io_inValid_22 = _T_632_22; // @[Switch.scala 53:21:@9517.4]
  assign switch_io_inValid_23 = _T_632_23; // @[Switch.scala 53:21:@9518.4]
  assign switch_io_inValid_24 = _T_632_24; // @[Switch.scala 53:21:@9519.4]
  assign switch_io_inValid_25 = _T_632_25; // @[Switch.scala 53:21:@9520.4]
  assign switch_io_inValid_26 = _T_632_26; // @[Switch.scala 53:21:@9521.4]
  assign switch_io_inValid_27 = _T_632_27; // @[Switch.scala 53:21:@9522.4]
  assign switch_io_inValid_28 = _T_632_28; // @[Switch.scala 53:21:@9523.4]
  assign switch_io_inValid_29 = _T_632_29; // @[Switch.scala 53:21:@9524.4]
  assign switch_io_inValid_30 = _T_632_30; // @[Switch.scala 53:21:@9525.4]
  assign switch_io_inValid_31 = _T_632_31; // @[Switch.scala 53:21:@9526.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_294_0 = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_294_1 = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_294_2 = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_294_3 = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_294_4 = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_294_5 = _RAND_5[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_294_6 = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_294_7 = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_294_8 = _RAND_8[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_294_9 = _RAND_9[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_294_10 = _RAND_10[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_294_11 = _RAND_11[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_294_12 = _RAND_12[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_294_13 = _RAND_13[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_294_14 = _RAND_14[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_294_15 = _RAND_15[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_294_16 = _RAND_16[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_294_17 = _RAND_17[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_294_18 = _RAND_18[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_294_19 = _RAND_19[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_294_20 = _RAND_20[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_294_21 = _RAND_21[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_294_22 = _RAND_22[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_294_23 = _RAND_23[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_294_24 = _RAND_24[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_294_25 = _RAND_25[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_294_26 = _RAND_26[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_294_27 = _RAND_27[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_294_28 = _RAND_28[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_294_29 = _RAND_29[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_294_30 = _RAND_30[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_294_31 = _RAND_31[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {2{`RANDOM}};
  _T_463_0 = _RAND_32[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {2{`RANDOM}};
  _T_463_1 = _RAND_33[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {2{`RANDOM}};
  _T_463_2 = _RAND_34[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {2{`RANDOM}};
  _T_463_3 = _RAND_35[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {2{`RANDOM}};
  _T_463_4 = _RAND_36[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {2{`RANDOM}};
  _T_463_5 = _RAND_37[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {2{`RANDOM}};
  _T_463_6 = _RAND_38[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {2{`RANDOM}};
  _T_463_7 = _RAND_39[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {2{`RANDOM}};
  _T_463_8 = _RAND_40[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {2{`RANDOM}};
  _T_463_9 = _RAND_41[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {2{`RANDOM}};
  _T_463_10 = _RAND_42[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {2{`RANDOM}};
  _T_463_11 = _RAND_43[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {2{`RANDOM}};
  _T_463_12 = _RAND_44[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {2{`RANDOM}};
  _T_463_13 = _RAND_45[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {2{`RANDOM}};
  _T_463_14 = _RAND_46[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {2{`RANDOM}};
  _T_463_15 = _RAND_47[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {2{`RANDOM}};
  _T_463_16 = _RAND_48[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {2{`RANDOM}};
  _T_463_17 = _RAND_49[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {2{`RANDOM}};
  _T_463_18 = _RAND_50[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {2{`RANDOM}};
  _T_463_19 = _RAND_51[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {2{`RANDOM}};
  _T_463_20 = _RAND_52[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {2{`RANDOM}};
  _T_463_21 = _RAND_53[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {2{`RANDOM}};
  _T_463_22 = _RAND_54[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {2{`RANDOM}};
  _T_463_23 = _RAND_55[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {2{`RANDOM}};
  _T_463_24 = _RAND_56[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {2{`RANDOM}};
  _T_463_25 = _RAND_57[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {2{`RANDOM}};
  _T_463_26 = _RAND_58[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {2{`RANDOM}};
  _T_463_27 = _RAND_59[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {2{`RANDOM}};
  _T_463_28 = _RAND_60[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {2{`RANDOM}};
  _T_463_29 = _RAND_61[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {2{`RANDOM}};
  _T_463_30 = _RAND_62[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {2{`RANDOM}};
  _T_463_31 = _RAND_63[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_632_0 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_632_1 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_632_2 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_632_3 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_632_4 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_632_5 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_632_6 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_632_7 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_632_8 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_632_9 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_632_10 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_632_11 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_632_12 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_632_13 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_632_14 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_632_15 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_632_16 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_632_17 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_632_18 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_632_19 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_632_20 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_632_21 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_632_22 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_632_23 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_632_24 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_632_25 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_632_26 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_632_27 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_632_28 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_632_29 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_632_30 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_632_31 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_801_0 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_801_1 = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_801_2 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_801_3 = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_801_4 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_801_5 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_801_6 = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_801_7 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_801_8 = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_801_9 = _RAND_105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_801_10 = _RAND_106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_801_11 = _RAND_107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_801_12 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_801_13 = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_801_14 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_801_15 = _RAND_111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_801_16 = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_801_17 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_801_18 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_801_19 = _RAND_115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_801_20 = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_801_21 = _RAND_117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_801_22 = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_801_23 = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_801_24 = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_801_25 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_801_26 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_801_27 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_801_28 = _RAND_124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T_801_29 = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_801_30 = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_801_31 = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {2{`RANDOM}};
  _T_970_0 = _RAND_128[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {2{`RANDOM}};
  _T_970_1 = _RAND_129[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {2{`RANDOM}};
  _T_970_2 = _RAND_130[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {2{`RANDOM}};
  _T_970_3 = _RAND_131[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {2{`RANDOM}};
  _T_970_4 = _RAND_132[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {2{`RANDOM}};
  _T_970_5 = _RAND_133[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {2{`RANDOM}};
  _T_970_6 = _RAND_134[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {2{`RANDOM}};
  _T_970_7 = _RAND_135[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {2{`RANDOM}};
  _T_970_8 = _RAND_136[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {2{`RANDOM}};
  _T_970_9 = _RAND_137[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {2{`RANDOM}};
  _T_970_10 = _RAND_138[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {2{`RANDOM}};
  _T_970_11 = _RAND_139[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {2{`RANDOM}};
  _T_970_12 = _RAND_140[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {2{`RANDOM}};
  _T_970_13 = _RAND_141[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {2{`RANDOM}};
  _T_970_14 = _RAND_142[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {2{`RANDOM}};
  _T_970_15 = _RAND_143[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {2{`RANDOM}};
  _T_970_16 = _RAND_144[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {2{`RANDOM}};
  _T_970_17 = _RAND_145[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {2{`RANDOM}};
  _T_970_18 = _RAND_146[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {2{`RANDOM}};
  _T_970_19 = _RAND_147[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {2{`RANDOM}};
  _T_970_20 = _RAND_148[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {2{`RANDOM}};
  _T_970_21 = _RAND_149[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {2{`RANDOM}};
  _T_970_22 = _RAND_150[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {2{`RANDOM}};
  _T_970_23 = _RAND_151[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {2{`RANDOM}};
  _T_970_24 = _RAND_152[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {2{`RANDOM}};
  _T_970_25 = _RAND_153[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {2{`RANDOM}};
  _T_970_26 = _RAND_154[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {2{`RANDOM}};
  _T_970_27 = _RAND_155[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {2{`RANDOM}};
  _T_970_28 = _RAND_156[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {2{`RANDOM}};
  _T_970_29 = _RAND_157[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {2{`RANDOM}};
  _T_970_30 = _RAND_158[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {2{`RANDOM}};
  _T_970_31 = _RAND_159[47:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _T_1139_0 = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _T_1139_1 = _RAND_161[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _T_1139_2 = _RAND_162[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _T_1139_3 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _T_1139_4 = _RAND_164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _T_1139_5 = _RAND_165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _T_1139_6 = _RAND_166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _T_1139_7 = _RAND_167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _T_1139_8 = _RAND_168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _T_1139_9 = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _T_1139_10 = _RAND_170[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _T_1139_11 = _RAND_171[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _T_1139_12 = _RAND_172[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _T_1139_13 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _T_1139_14 = _RAND_174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _T_1139_15 = _RAND_175[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _T_1139_16 = _RAND_176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _T_1139_17 = _RAND_177[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _T_1139_18 = _RAND_178[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _T_1139_19 = _RAND_179[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  _T_1139_20 = _RAND_180[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _T_1139_21 = _RAND_181[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _T_1139_22 = _RAND_182[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _T_1139_23 = _RAND_183[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _T_1139_24 = _RAND_184[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _T_1139_25 = _RAND_185[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _T_1139_26 = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _T_1139_27 = _RAND_187[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _T_1139_28 = _RAND_188[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _T_1139_29 = _RAND_189[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _T_1139_30 = _RAND_190[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  _T_1139_31 = _RAND_191[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    _T_294_0 <= io_inAddr_0;
    _T_294_1 <= io_inAddr_1;
    _T_294_2 <= io_inAddr_2;
    _T_294_3 <= io_inAddr_3;
    _T_294_4 <= io_inAddr_4;
    _T_294_5 <= io_inAddr_5;
    _T_294_6 <= io_inAddr_6;
    _T_294_7 <= io_inAddr_7;
    _T_294_8 <= io_inAddr_8;
    _T_294_9 <= io_inAddr_9;
    _T_294_10 <= io_inAddr_10;
    _T_294_11 <= io_inAddr_11;
    _T_294_12 <= io_inAddr_12;
    _T_294_13 <= io_inAddr_13;
    _T_294_14 <= io_inAddr_14;
    _T_294_15 <= io_inAddr_15;
    _T_294_16 <= io_inAddr_16;
    _T_294_17 <= io_inAddr_17;
    _T_294_18 <= io_inAddr_18;
    _T_294_19 <= io_inAddr_19;
    _T_294_20 <= io_inAddr_20;
    _T_294_21 <= io_inAddr_21;
    _T_294_22 <= io_inAddr_22;
    _T_294_23 <= io_inAddr_23;
    _T_294_24 <= io_inAddr_24;
    _T_294_25 <= io_inAddr_25;
    _T_294_26 <= io_inAddr_26;
    _T_294_27 <= io_inAddr_27;
    _T_294_28 <= io_inAddr_28;
    _T_294_29 <= io_inAddr_29;
    _T_294_30 <= io_inAddr_30;
    _T_294_31 <= io_inAddr_31;
    _T_463_0 <= io_inData_0;
    _T_463_1 <= io_inData_1;
    _T_463_2 <= io_inData_2;
    _T_463_3 <= io_inData_3;
    _T_463_4 <= io_inData_4;
    _T_463_5 <= io_inData_5;
    _T_463_6 <= io_inData_6;
    _T_463_7 <= io_inData_7;
    _T_463_8 <= io_inData_8;
    _T_463_9 <= io_inData_9;
    _T_463_10 <= io_inData_10;
    _T_463_11 <= io_inData_11;
    _T_463_12 <= io_inData_12;
    _T_463_13 <= io_inData_13;
    _T_463_14 <= io_inData_14;
    _T_463_15 <= io_inData_15;
    _T_463_16 <= io_inData_16;
    _T_463_17 <= io_inData_17;
    _T_463_18 <= io_inData_18;
    _T_463_19 <= io_inData_19;
    _T_463_20 <= io_inData_20;
    _T_463_21 <= io_inData_21;
    _T_463_22 <= io_inData_22;
    _T_463_23 <= io_inData_23;
    _T_463_24 <= io_inData_24;
    _T_463_25 <= io_inData_25;
    _T_463_26 <= io_inData_26;
    _T_463_27 <= io_inData_27;
    _T_463_28 <= io_inData_28;
    _T_463_29 <= io_inData_29;
    _T_463_30 <= io_inData_30;
    _T_463_31 <= io_inData_31;
    _T_632_0 <= io_inValid_0;
    _T_632_1 <= io_inValid_1;
    _T_632_2 <= io_inValid_2;
    _T_632_3 <= io_inValid_3;
    _T_632_4 <= io_inValid_4;
    _T_632_5 <= io_inValid_5;
    _T_632_6 <= io_inValid_6;
    _T_632_7 <= io_inValid_7;
    _T_632_8 <= io_inValid_8;
    _T_632_9 <= io_inValid_9;
    _T_632_10 <= io_inValid_10;
    _T_632_11 <= io_inValid_11;
    _T_632_12 <= io_inValid_12;
    _T_632_13 <= io_inValid_13;
    _T_632_14 <= io_inValid_14;
    _T_632_15 <= io_inValid_15;
    _T_632_16 <= io_inValid_16;
    _T_632_17 <= io_inValid_17;
    _T_632_18 <= io_inValid_18;
    _T_632_19 <= io_inValid_19;
    _T_632_20 <= io_inValid_20;
    _T_632_21 <= io_inValid_21;
    _T_632_22 <= io_inValid_22;
    _T_632_23 <= io_inValid_23;
    _T_632_24 <= io_inValid_24;
    _T_632_25 <= io_inValid_25;
    _T_632_26 <= io_inValid_26;
    _T_632_27 <= io_inValid_27;
    _T_632_28 <= io_inValid_28;
    _T_632_29 <= io_inValid_29;
    _T_632_30 <= io_inValid_30;
    _T_632_31 <= io_inValid_31;
    _T_801_0 <= switch_io_outAck_0;
    _T_801_1 <= switch_io_outAck_1;
    _T_801_2 <= switch_io_outAck_2;
    _T_801_3 <= switch_io_outAck_3;
    _T_801_4 <= switch_io_outAck_4;
    _T_801_5 <= switch_io_outAck_5;
    _T_801_6 <= switch_io_outAck_6;
    _T_801_7 <= switch_io_outAck_7;
    _T_801_8 <= switch_io_outAck_8;
    _T_801_9 <= switch_io_outAck_9;
    _T_801_10 <= switch_io_outAck_10;
    _T_801_11 <= switch_io_outAck_11;
    _T_801_12 <= switch_io_outAck_12;
    _T_801_13 <= switch_io_outAck_13;
    _T_801_14 <= switch_io_outAck_14;
    _T_801_15 <= switch_io_outAck_15;
    _T_801_16 <= switch_io_outAck_16;
    _T_801_17 <= switch_io_outAck_17;
    _T_801_18 <= switch_io_outAck_18;
    _T_801_19 <= switch_io_outAck_19;
    _T_801_20 <= switch_io_outAck_20;
    _T_801_21 <= switch_io_outAck_21;
    _T_801_22 <= switch_io_outAck_22;
    _T_801_23 <= switch_io_outAck_23;
    _T_801_24 <= switch_io_outAck_24;
    _T_801_25 <= switch_io_outAck_25;
    _T_801_26 <= switch_io_outAck_26;
    _T_801_27 <= switch_io_outAck_27;
    _T_801_28 <= switch_io_outAck_28;
    _T_801_29 <= switch_io_outAck_29;
    _T_801_30 <= switch_io_outAck_30;
    _T_801_31 <= switch_io_outAck_31;
    _T_970_0 <= switch_io_outData_0;
    _T_970_1 <= switch_io_outData_1;
    _T_970_2 <= switch_io_outData_2;
    _T_970_3 <= switch_io_outData_3;
    _T_970_4 <= switch_io_outData_4;
    _T_970_5 <= switch_io_outData_5;
    _T_970_6 <= switch_io_outData_6;
    _T_970_7 <= switch_io_outData_7;
    _T_970_8 <= switch_io_outData_8;
    _T_970_9 <= switch_io_outData_9;
    _T_970_10 <= switch_io_outData_10;
    _T_970_11 <= switch_io_outData_11;
    _T_970_12 <= switch_io_outData_12;
    _T_970_13 <= switch_io_outData_13;
    _T_970_14 <= switch_io_outData_14;
    _T_970_15 <= switch_io_outData_15;
    _T_970_16 <= switch_io_outData_16;
    _T_970_17 <= switch_io_outData_17;
    _T_970_18 <= switch_io_outData_18;
    _T_970_19 <= switch_io_outData_19;
    _T_970_20 <= switch_io_outData_20;
    _T_970_21 <= switch_io_outData_21;
    _T_970_22 <= switch_io_outData_22;
    _T_970_23 <= switch_io_outData_23;
    _T_970_24 <= switch_io_outData_24;
    _T_970_25 <= switch_io_outData_25;
    _T_970_26 <= switch_io_outData_26;
    _T_970_27 <= switch_io_outData_27;
    _T_970_28 <= switch_io_outData_28;
    _T_970_29 <= switch_io_outData_29;
    _T_970_30 <= switch_io_outData_30;
    _T_970_31 <= switch_io_outData_31;
    _T_1139_0 <= switch_io_outValid_0;
    _T_1139_1 <= switch_io_outValid_1;
    _T_1139_2 <= switch_io_outValid_2;
    _T_1139_3 <= switch_io_outValid_3;
    _T_1139_4 <= switch_io_outValid_4;
    _T_1139_5 <= switch_io_outValid_5;
    _T_1139_6 <= switch_io_outValid_6;
    _T_1139_7 <= switch_io_outValid_7;
    _T_1139_8 <= switch_io_outValid_8;
    _T_1139_9 <= switch_io_outValid_9;
    _T_1139_10 <= switch_io_outValid_10;
    _T_1139_11 <= switch_io_outValid_11;
    _T_1139_12 <= switch_io_outValid_12;
    _T_1139_13 <= switch_io_outValid_13;
    _T_1139_14 <= switch_io_outValid_14;
    _T_1139_15 <= switch_io_outValid_15;
    _T_1139_16 <= switch_io_outValid_16;
    _T_1139_17 <= switch_io_outValid_17;
    _T_1139_18 <= switch_io_outValid_18;
    _T_1139_19 <= switch_io_outValid_19;
    _T_1139_20 <= switch_io_outValid_20;
    _T_1139_21 <= switch_io_outValid_21;
    _T_1139_22 <= switch_io_outValid_22;
    _T_1139_23 <= switch_io_outValid_23;
    _T_1139_24 <= switch_io_outValid_24;
    _T_1139_25 <= switch_io_outValid_25;
    _T_1139_26 <= switch_io_outValid_26;
    _T_1139_27 <= switch_io_outValid_27;
    _T_1139_28 <= switch_io_outValid_28;
    _T_1139_29 <= switch_io_outValid_29;
    _T_1139_30 <= switch_io_outValid_30;
    _T_1139_31 <= switch_io_outValid_31;
  end
endmodule
